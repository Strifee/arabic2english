RÅDETS FÖRSTA DIREKTIV av den 23 juli 1962 om fastställande av vissa gemensamma regler för internationella transporter (yrkesmässiga godstransporter på väg)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 75.1 i detta,
med beaktande av Europaparlamentets yttrande, och
med beaktande av följande: Antagandet av en gemensam transportpolitik innebär bland annat att man fastställer gemensamma regler för internationella godstransporter på väg till eller från en medlemsstat eller genom en eller flera medlemsstater.
Den gemensamma marknadens successiva uppbyggnad får inte försvåras av hinder inom transportsektorn. Det är nödvändigt att säkerställa en gradvis utbyggnad av de internationella godstransporterna på väg med tanke på utvecklingen av handeln och varuflödena inom gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Senast vid utgången av år 1962 skall varje medlemsstat, på det sätt som fastställts i punkterna 2 och 3 av denna artikel, liberalisera de typer av internationella yrkesmässiga vägtransporter som berör andra medlemsstater och som är förtecknade i bilagorna 1 och 2 till detta direktiv, om sådan transport utförs till eller från medlemsstaten eller passerar dess territorium i transit.
2. De typer av transporter som är förtecknade i bilaga 1 skall vara undantagna från kvoterings- eller tillståndssystem.
3. De typer av transporter som är förtecknade i bilaga 2 skall inte längre regleras av något kvoteringssystem. Dock får tillståndskrav behållas som villkor för denna transportverksamhet, förutsatt att ingen restriktion av kvantitativ natur förekommer; i sådant fall skall medlemsstaterna ombesörja att beslut i tillståndsärenden fattas senast fem dagar efter mottagandet av tillståndsansökan.
4. De båda bilagorna till detta direktiv skall utgöra en del av själva direktivet.
Artikel 2
Medlemsstaterna skall senast tre månader efter detta direktivs ikraftträdande och i vart fall före utgången av år 1962 underrätta kommissionen om de åtgärder som vidtagits för att genomföra det.
Artikel 3
Detta direktiv skall inte påverka de villkor som en medlemsstat uppställer för sina egna medborgare för att bedriva sådan verksamhet som avses i detta direktiv.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EEG) nr 1397/68 av den 6 september 1968 om ändring av förordning nr 474/67/EEG om förutfastställelse av exportbidraget för ris och brutet ris
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning nr 359/67/EEG av den 25 juli 1967 om den gemensamma organisationen av marknaden för ris(1), särskilt artikel 17.6 i denna, och
med beaktande av följande: Enligt artikel 17.4 i förordning nr 359/67/EEG får det exportbidrag som gäller den dag då ansökan om exportlicens inlämnas, tillämpas vid export som sker inom licensens giltighetstid och att ett korrektionsbelopp i så fall skall användas för exportbidraget. Enligt artikel 1 i kommissionens förordning nr 474/67/EEG om förutfastställelse av exportbidraget för ris och brutet ris(2), är korrektionsbeloppet lika med skillnaden mellan cif-priset och cif-priset vid terminsköp.
Exportlicenser för ris och brutet ris gäller till och med den femte månaden efter utfärdandemånaden men det finns för sådana produkter sällan en verkligt representativ terminsmarknad, annat än för den eller de närmaste terminerna. Det bör därför vara möjligt att fastställa ett korrektionsbelopp som är lägre än den ovannämnda skillnaden.
Det är därför nödvändigt att ändra förordning nr 474/67/EEG.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 1 i förordning nr 474/67/EEG skall första och andra stycket ersättas med följande:
"När det exportbidrag för ris och brutet ris som anges i artikel 17.4 första stycket i förordning nr 359/67/EEG förutfastställs, skall exportbidraget vara det som gäller för export den dag då ansökan om exportlicens inlämnas - med avdrag för ett belopp som inte överstiger skillnaden mellan cif-priset för terminsköp och cif-priset, när det förstnämnda överstiger det sistnämnda med mer än 0,025 räkneenheter per 100 kg,
- med tillägg av ett belopp som inte överstiger skillnaden mellan cif-priset och cif-priset för terminsköp, när det förstnämnda överstiger det sistnämnda med mer än 0,025 räkneenheter per 100 kg.
Under tiden mellan de veckovisa fastställelserna skall det bidragsbelopp som gäller vid förutfastställelse endast justeras om tillämpningen av ovannämnda bestämmelse medför att beloppet ändras med mer än 0,025 räkneenheter per 100 kg."
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS DIREKTIV av den 20 mars 1970 om tillnärmning av medlemsstaternas lagstiftning om åtgärder mot luftförorening genom avgaser från motorfordon (70/220/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: Förordningen av den 14 oktober 1968 med ändring i Straßenverkehrs-Zulassungs-Ordnung publicerades i Tyskland i Bundesgesetzblatt Del 1 den 18 oktober 1968. Denna förordning innehåller bestämmelser om åtgärder mot luftföroreningar från förbränningsmotorer i motorfordon. Bestämmelserna kommer att träda i kraft den 1 oktober 1970.
Förordningen av den 31 mars 1969 om "Sammansättningen hos avgaser som släpps ut från bensinmotorer i motorfordon" publicerades i Frankrike den 17 maj 1969 i Journal officiel. Förordningen gäller - från och med den 1 september 1971 för typgodkända fordon med en ny motortyp, dvs. en motortyp som inte tidigare monterats i ett typgodkänt fordon,
- från och med den 1 september 1972 för fordon som tas i bruk för första gången.
Varje medlemsstat som skall utfärda ett nationellt typgodkännande för en fordonstyp måste genom det nämnda meddelandet kunna förvissa sig om att fordonstypen genomgått de prov som krävs enligt detta direktiv. Därför bör varje medlemsstat underrätta övriga medlemsstater om sina resultat genom att sända dem en kopia av det meddelande som upprättats för varje motorfordonstyp som provats.
Vidare måste de tekniska kraven snabbt anpassas med hänsyn till tekniska framsteg. Därför bör det förfarande kunna tillämpas som fastslås i artikel 13 i rådets direktiv av den 6 februari 1970 om typgodkännande av motorfordon och släpvagnar till dessa fordon.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I detta direktiv avses med fordon varje fordon med förbränningsmotor med styrd tändning, avsett att användas på väg, med eller utan karosseri, som har minst fyra hjul, med en tillåten totalvikt på minst 400 kg och som är konstruerat för en högsta hastighet som uppgår till minst 50 km/tim. Jordbrukstraktorer, lantbruksmaskiner och arbetsfordon är undantagna.
Artikel 2
Ingen medlemsstat får vägra att bevilja EEG-typgodkännande eller nationellt typgodkännande för ett fordon av skäl som hänför sig till luftförorening genom gaser från förbränningsmotorer med styrd tändning i fordonet - från och med den 1 oktober 1970, om fordonet uppfyller både kraven i bilaga 1, med undantag för kraven i punkt 3.2.1.1 och 3.2.2.1, och kraven i bilagorna 2, 4, 5 och 6,
- från och med den 1 oktober 1971, om fordonet även uppfyller kraven i punkt 3.2.1.1 och 3.2.2.1 i bilaga 1 och kraven i bilaga 3.
Artikel 3
1. När en ansökan kommer in från en tillverkare eller dennes representant skall de behöriga myndigheterna i den berörda medlemsstaten fylla i uppgifterna i meddelandet enligt bilaga 7. En kopia av meddelandet skall sändas till övriga medlemsstater och till sökanden. Andra medlemsstater som får en ansökan om nationellt typgodkännande för samma fordonstyp skall godta det nämnda dokumentet som bevis för att de föreskrivna proven har utförts.
2. Bestämmelserna i 1 skall upphävas så snart rådets direktiv av den 6 februari 1970 om typgodkännande av motorfordon och släpvagnar till dessa fordon träder i kraft.
Artikel 4
Den medlemsstat som har beviljat ett typgodkännande skall vidta de åtgärder som krävs för att säkerställa att den underrättas om varje ändring i fråga om delar eller egenskaper som avses i punkt 1.1 i bilaga 1. De behöriga myndigheterna i medlemsstaten skall avgöra om nya prov måste utföras på den ändrade prototypen och om en ny rapport måste upprättas. Om dessa prov visar att kraven i detta direktiv inte uppfylls skall ändringen inte godkännas.
Artikel 5
De ändringar som är nödvändiga för att anpassa kraven i bilaga 1 7 till tekniska framsteg skall beslutas enligt det förfarande som fastslås i artikel 13 i rådets direktiv av den 6 februari 1970 om typgodkännande av motorfordon och släpvagnar till dessa fordon.
Artikel 6
1. Medlemsstaterna skall anta bestämmelser som innehåller de krav som är nödvändiga för att följa detta direktiv före den 30 juni 1970 och skall genast underrätta kommissionen om detta.
2. Medlemsstaterna skall se till att till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 7
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 24 juli 1973 om åtgärder för att dämpa verkningarna av svårigheter vid försörjningen med råolja eller petroleumprodukter (73/238/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 103 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande,
med beaktande av Ekonomiska och sociala kommitténs yttrande, och
med beaktande av följande: Fastställandet av en gemensam energipolitik tillhör de mål som gemenskaperna har ställt upp.
Råolja och petroleumprodukter är av allt större betydelse för gemenskapens försörjning med energi. Varje svårighet, även om den är tillfällig, som väsentligt begränsar leveranserna av dessa produkter, skulle kunna vålla allvarliga störningar i gemenskapens ekonomiska verksamhet. Gemenskapen bör därför kunna upphäva eller i vart fall minska de skadliga verkningar som skulle kunna uppstå i ett sådant fall.
Förfaranden och instrument, lämpade att säkerställa ett snabbt genomförande av de åtgärder som är avsedda att dämpa försörjningssvårigheterna i fråga om råolja eller petroleumprodukter, bör fastställas i förväg.
Medlemsstaterna bör därför ges de nödvändiga befogenheterna för att, om så erfordras, omedelbart kunna vidta lämpliga åtgärder i enlighet med bestämmelserna i fördraget, särskilt artikel 103 i detta.
En viss överensstämmelse mellan dessa befogenheter är nödvändig för att underlätta en samordning av de enskilda staternas åtgärder inom ramen för samråd på gemenskapsnivå.
I övrigt är det lämpligt att omedelbart bilda ett samrådsorgan som kan underlätta samordningen av konkreta åtgärder som medlemsstaterna kan ha vidtagit eller planerat på detta område.
Det är nödvändigt att varje medlemsstat upprättar en plan som kan följas vid svårigheter i försörjningen med råolja eller petroleumprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 3
1. Om svårigheter i försörjningen med råolja eller petroleumprodukter uppkommer i gemenskapen eller i en av medlemsstaterna skall kommissionen på begäran av en medlemsstat eller på eget initiativ snarast sammankalla en grupp av företrädare för medlemsstaterna, i vilken kommissionens företrädare skall vara ordförande.
Artikel 5
Medlemsstaterna skall senast den 30 juni 1974 sätta i kraft de rättsliga och administrativa bestämmelser som är nödvändiga för att följa detta direktiv.
Artikel 6
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EKSG, EEG, Euratom) nr 559/73 av den 26 februari 1973 om ändring av rådets förordning (EEG, Euratom, EKSG) nr 260/68 om villkoren för och förfarandet vid skatt till Europeiska gemenskaperna
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättande av ett gemensamt råd och en gemensam kommission,
med beaktande av protokollet om immunitet och privilegier för Europeiska gemenskaperna, särskilt artikel 13 i detta,
med beaktande av kommissionens förslag, och
med beaktande av följande: Med hänsyn till en dom som nyligen avkunnats av domstolen samt till vissa tvingande sociala krav verkar det önskvärt att ändra en bestämmelse i rådets förordning (EEG, Euratom, EKSG) nr 260/681 av den 29 februari 1968 om villkoren för och förfarandet vid skatt till Europeiska gemenskaperna, senast ändrad genom förordning (Euratom, EKSG, EEG) nr 2531/722.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Rådets förordning (EEG, Euratom, EKSG) nr 260/68 av den 29 februari 1968 ändras på följande sätt:
I artikel 3.3 a första strecksatsen skall "familjeförsörjartillägg" ersättas med "hushållstillägg".
Artikel 2
RÅDETS DIREKTIV av den 17 december 1973 om tillnärmning av medlemsstaternas lagstiftning om inredningsdetaljer i motorfordon (passagerarutrymmets inre delar frånsett inre backspeglar, manöverorganens utformning, taket eller det öppningsbara taket, ryggstödet och sätenas baksida) (74/60/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: De tekniska krav som motorfordon måste uppfylla enligt nationell lagstiftning gäller bl.a. inredning avsedd att skydda föraren och passagerarna.
Dessa krav skiljer sig åt i de olika medlemsstaterna. Det är därför nödvändigt att alla medlemsstater antar samma krav, antingen som tillägg till eller i stället för sina nuvarande bestämmelser, särskilt för att det förfarande med EEG-typgodkännande, som behandlats i rådets direktiv av den 6 februari 1970(3) om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon, skall kunna tillämpas på alla fordonstyper.
Gemensamma krav för inre backspeglar har lagts fram genom rådets direktiv av den 1 mars 1971(4) och krav bör också utarbetas för passagerarutrymmets inredningsdetaljer, manöverorganens utformning, taket och ryggstöden och sätenas baksida. Ytterligare krav avseende inredning kommer att antas senare, särskilt i fråga om förankringspunkter för bilbälten och säten, huvudstöd, skydd för föraren mot styranordningen och identifikation av manöverorganen.
Harmoniserade krav bör minska risken för eller graden av skador i samband med olyckor som motorfordonsförare kan bli offer för och trygga trafiksäkerheten inom hela gemenskapen.
När det gäller tekniska krav är det lämpligt att huvudsakligen tillämpa de som antagits av FNs ekonomiska kommission för Europa i reglemente nr 21 ("Enhetliga krav om godkännande av fordon med avseende på inredningar i dessa"), vilka återges i en bilaga till överenskommelsen av den 20 mars 1958 om antagande av enhetliga villkor för godkännande och ömsesidigt erkännande av utrustning och delar för motorfordon.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I detta direktiv avses med fordon varje motorfordon i kategori M1 (definieras i bilaga 1 till direktivet av den 6 februari 1970) som är avsett att användas på väg, har minst fyra hjul och är konstruerat för en högsta hastighet som överstiger 25 km/tim.
Artikel 2
Ingen medlemsstat får vägra att bevilja EEG-typgodkännande eller nationellt typgodkännande för ett fordon av skäl som hänför sig till sådana inredningsdetaljer som
- passagerarutrymmets inre delar frånsett inre backspeglar, - manöverorganens utformning,
- taket eller det öppningsbara taket,
- ryggstödet eller sätenas baksida,
om dessa uppfyller kraven i bilagorna.
Artikel 3
Ingen medlemsstat får vägra eller förbjuda att ett fordon saluförs, registreras, tas i bruk eller används, av skäl som hänför sig till - passagerarutrymmets inre delar frånsett inre backspeglar,
- manöverorganens utformning,
- taket eller det öppningsbara taket,
- ryggstödet eller sätenas baksida,
om dessa inredningsdetaljer uppfyller kraven i bilagorna.
Artikel 4
Den medlemsstat som har beviljat EEG-typgodkännande måste vidta de åtgärder som krävs för att hålla sig informerad om varje ändring av en sådan del eller egenskap som avses i bilaga 1 punkt 2.2. De behöriga myndigheterna i staten skall avgöra om nya provningar behöver utföras på den ändrade fordonstypen och en ny rapport utformas. Om dessa provningar visar att kraven i detta direktiv inte uppfylls skall ändringen inte godkännas.
Artikel 5
De ändringar som är nödvändiga för att anpassa kraven i bilagorna till den tekniska utvecklingen skall beslutas enligt det förfarande som föreskrivs i artikel 13 i rådets direktiv av den 6 februari 1970 om en anpassning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon.
Artikel 6
1. Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv inom 18 månader från dagen för anmälan och skall genast underrätta kommissionen om detta.
2. Medlemsstaterna ska se till att till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 7
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EEG) nr 668/74 av den 28 mars 1974 om ändring av förordning (EEG) nr 922/72 om allmänna tillämpningsföreskrifter för stöd till silkesodling
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 845/72(1) av den 24 april 1972 om särskilda åtgärder för att främja silkesodling, särskilt artikel 2.4 i denna,
med beaktande av kommissionens förslag, och
med beaktande av följande: I förordning (EEG) nr 922/72(2), ändrad genom förordning (EEG) nr 884/73(3), fastställer rådet allmänna tillämpningsföreskrifter för stöd till silkesmaskar för odlingsåren 1972/1973 och 1973/1974. Erfarenheten har visat att det är lämpligt att fortsätta att tillämpa förordningen under kommande odlingsår.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 1 i förordning (EEG) nr 922/72 skall orden "för odlingsåren 1972/1973 och 1973/1974" utgå.
Artikel 2
Denna förordning skall tillämpas från och med den 1 april 1974.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS DIREKTIV av den 17 december 1974 om utvidgande av tillämpningsområdet för direktiv nr 64/221/EEG om samordningen av särskilda åtgärder som gäller utländska medborgares rörlighet och bosättning och som är berättigade med hänsyn till allmän ordning, säkerhet eller hälsa till att även omfatta medborgare i en medlemsstat som begagnar sig av rätten att stanna kvar inom en annan medlemsstats territorium efter att ha verkat där som egna företagare (75/35/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
med beaktande av följande: Direktiv nr 64/221/EEG (3) samordnade särskilda åtgärder som gäller utländska medborgares rörlighet och bosättning och som är berättigade med hänsyn till allmän ordning, säkerhet eller hälsa, och direktiv nr 75/34/EEG (4) fastställde enligt vilka villkor medborgare i en medlemsstat skall ha rätt att stanna kvar inom en annan medlemsstats territorium efter att ha varit verksamma där som egna företagare.
Direktiv nr 64/221/EEG bör därför gälla för personer som omfattas av direktiv 75/34/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv nr 64/221/EEG skall gälla för medborgare i medlemsstaterna och deras familjemedlemmar som har rätt att stanna kvar inom en medlemsstats territorium i enlighet med direktiv nr 75/34/EEG
Artikel 2
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 20 maj 1975 om tillnärmning av medlemsstaternas lagar och andra författningar beträffande aerosolbehållare (75/324/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: I vissa medlemsstater är det ett obligatoriskt krav att aerosolbehållare motsvarar vissa tekniska specifikationer. Sådana specifikationer varierar från medlemsstat till medlemsstat, vilket hindrar handeln inom gemenskapen.
Dessa hinder för upprättandet av en väl fungerande gemensam marknad kan avlägsnas, om alla medlemsstater antar samma specifikationer, antingen utöver eller i stället för dem som fastlagts i deras nuvarande lagstiftning, och dessa specifikationer speciellt avser tillverkning och fyllning av aerosolbehållare och den volym de får anges ha.
Med hänsyn till det tekniska kunnande som för närvarande har uppnåtts skall tillämpningsområdet för detta direktiv begränsas till aerosolbehållare av metall, glas och plast.
De tekniska specifikationer som anges i bilagan till detta direktiv kommer inom kort att behöva anpassas till tekniska framsteg. För att underlätta att nödvändiga åtgärder genomförs på ett effektivt sätt skall former fastställas för ett nära samarbete mellan medlemsstaterna och kommissionen inom ramen för en kommitté för anpassning av direktivet om aerosolbehållare till teknisk utveckling.
Det är möjligt att vissa aerosolbehållare som finns på marknaden kan innebära en säkerhetsrisk, trots att de uppfyller kraven i detta direktiv och dess bilaga. Ett förfarande måste därför fastläggas för att motverka denna risk.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Detta direktiv skall gälla aerosolbehållare enligt definitionen i artikel 2 med undantag av sådana som har mindre volym än maximalt 50 ml och sådana som har större volym än vad som anges i punkt 3.1, 4.1.1, 4.2.1, 5.1 och 5.2 i bilagan till detta direktiv.
Artikel 2
I detta direktiv avses med aerosolbehållare varje behållare som inte kan återanvändas, är tillverkad av metall, glas eller plast, innehåller gas som komprimerats, kondenserats eller lösts under tryck, med eller utan vätska, pasta eller pulver, och som är försedd med en utlösningsanordning för att spruta ut innehållet som en suspension av fasta eller flytande partiklar i gas, som lödder, pasta eller pulver eller i flytande tillstånd.
Artikel 3
Den som svarar för att aerosolbehållare släpps ut på marknaden skall förse dessa med symbolen "3" (omvänt epsilon) som bevis för att de uppfyller kraven i detta direktiv och dess bilaga.
Artikel 4
Medlemsstaterna får inte, av skäl som sammanhänger med kraven i detta direktiv och dess bilaga, begränsa, hindra eller förbjuda att sådana aerosolbehållare släpps ut på marknaden som uppfyller kraven i detta direktiv och dess bilaga.
Artikel 6
1. En kommitté för anpassning av direktivet om aerosolbehållare till teknisk utveckling, nedan kallad "kommittén", inrättas härmed. Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
2. Kommittén skall själv fastställa sin arbetsordning.
Artikel 7
1. När det förfarande som anges i denna artikel skall tillämpas, skall ordföranden hänskjuta ärendet till kommittén, antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom två månader. Yttranden skall antas med 41 rösters majoritet, varvid medlemsstaternas röster skall vägas enligt förslagets artikel 148.2. Ordföranden får inte rösta.
3. a) Kommissionen skall själv anta förslaget, om det har tillstyrkts av kommittén.
b) Om förslaget inte har tillstyrkts av kommittén eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet åtgärder. Rådet skall fatta sitt beslut med kvalificerad majoritet.
c) Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen anta förslaget till åtgärder.
Artikel 8
1. Varje aerosolbehållare skall vara försedd med följande uppgifter i väl synlig, läslig och varaktig skrift som, om förpackningen är av liten volym (högst 150 ml), kan anbringas på en vidfäst etikett; denna bestämmelse gäller utöver krav i andra av gemenskapens direktiv, särskilt direktiven om farliga ämnen och beredningar: a) Namn och adress eller varumärke för den person som svarar för utsläppandet på marknaden av aerosolbehållaren.
b) Symbolen "3" (omvänt epsilon) som bevis för att produkten motsvarar kraven i detta direktiv.
c) Kodbeteckningar som gör det möjligt att identifiera varuparti.
d) De uppgifter som anges i punkt 2.2 i bilagan.
e) Innehållets nettovikt och -volym.
2. Medlemsstaterna kan ställa som villkor för försäljning inom sitt territorium att nationalspråket eller -språken används för förpackningstexten.
Artikel 9
Medlemsstaterna skall vidta nödvändiga åtgärder för att förhindra att märken eller påskrift som kan förväxlas med symbolen "3" (omvänt epsilon) används på aerosolbehållare.
Artikel 10
1. Om någon medlemsstat uppmärksammar att en eller flera aerosolbehållare på goda grunder kan antas medföra fara för hälsa och säkerhet, trots att den eller de motsvarar kraven i detta direktiv, har denna stat rätt att provisoriskt förbjuda försäljning av dessa behållare inom sina nationsgränser eller förena försäljningen med särskilda villkor. Medlemsstaten skall omedelbart underrätta de andra medlemsstaterna och kommissionen om detta och ange skälen till sitt beslut.
2. Kommissionen skall inom sex veckor rådfråga berörda medlemsstater och därefter utan dröjsmål avge sitt yttrande och vidta lämpliga åtgärder.
3. Om kommissionen anser att direktivet behöver bearbetas i tekniskt avseende, skall sådana bearbetningar godkännas av antingen kommissionen eller rådet i enlighet med det förfarande som anges i artikel 7. Om så är fallet kan den medlemsstat som infört säkerhetsåtgärder behålla dessa, tills de nya bestämmelserna trätt i kraft.
Artikel 11
1. Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv inom 18 månader efter dagen för anmälan och skall genast underrätta kommissionen om detta.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 12
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 26 juni 1975 om ändring av direktiven 66/400/EEG, 66/401/EEG, 66/402/EEG, 66/403/EEG och 69/208/EEG om saluföring av betutsäde, utsäde av foderväxter, utsäde av stråsäd, utsädespotatis och utsäde av olje- och spånadsväxter (75/444/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 43 och 100 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: Vissa direktiv om saluföring av utsäde bör ändras av nedan angivna skäl.
Under den tid då direktiven tillämpats har det framkommit att små förpackningar av betutsäde och utsäde av foderväxter utgör en handelsvara inom gemenskapen.
Det är följaktligen lämpligt att harmonisera denna sektor som hittills har omfattats av nationell lagstiftning.
Det är i detta sammanhang lämpligt att, å ena sidan, underlätta saluföring och plombering av sådana små förpackningar och, å andra sidan, göra tillräcklig äkthetskontroll av utsädet obligatorisk.
Vissa av ovannämnda direktiv innehåller bestämmelser om att likvärdighet hos utsäde som skördats i andra länder, särskilt i tredje land, fr.o.m. den 1 juli 1975 inte längre får beslutas nationellt av medlemsstaterna. Eftersom det inte har varit möjligt att utföra gemensam undersökning av utsäde av foder-, olje- och spånadsväxter i samtliga fall bör dock ovannämnda period förlängas för dessa utsäden för att undvika att nuvarande handelsförbindelser störs.
Det är lämpligt att tillåta att medlemsstaterna antar bestämmelser som underlättar plombering av små förpackningar med utsäde av stråsäd, utsädespotatis och utsäde av olje- och spånadsväxter.
Det är också nödvändigt att göra vissa ändringar av det sätt på vilket utsädeskvantiteterna anges.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Rådets direktiv 66/400/EEG(3) av den 14 juni 1966 om saluföring av betutsäde, senast ändrat genom direktiv 73/438/EEG(4) skall ändras på följande sätt: 1. Följande stycke skall läggas till artikel 2.1:
"G. EEG-småförpackningar: förpackningar med följande certifikatutsäden: - Monogermt frö eller tekniskt monogermfrö (precisionsfrö): högst 100 000 frögyttringar eller frön eller med en nettovikt om 2,5 kg, exklusive, i förekommande fall, pesticider i pulverform, pelleteringsmedel eller andra fasta tillsatser.
- Annat frö än monogermt frö eller tekniskt monogermfrö (precisionsfrö): högsta nettovikt 10 kg, exklusive, i förekommande fall, pesticider i pulverform, pelleteringsmedel eller andra fasta tillsatser."
1. Medlemsstaterna skall kräva att förpackningar med basutsäde och certifikatutsäde, förutom då utsäde av den sistnämnda kategorin förpackas i EEG-småförpackningar, skall plomberas officiellt på sådant sätt att plomberingen skadas och inte kan anbringas på nytt när förpackningen öppnats.
2. Medlemsstaterna skall kräva, förutom för EEG-småförpackningar, att förpackningar inte omplomberas, varken en eller flera gånger, annat än genom officiell plombering. Om förpackningar omplomberas, skall detta samt ansvarig myndighet och datum för omplombering anges på den etikett som krävs enligt artikel 11.1.
3. Medlemsstaterna skall kräva att EEG-småförpackningar plomberas på sådant sätt att plomberingen skadas och inte kan anbringas på nytt när förpackningen öppnats. Förpackningar får inte omplomberas, varken en eller flera gånger, annat än under officiell övervakning.
4. Medlemsstaterna får anta bestämmelser om undantag från punkt 1 och 2 för småförpackningar med basutsäde."
4. Det inledande avsnittet i artikel 11.1 skall ersättas med följande:
"1. Medlemsstaterna skall kräva att förpackningar med basutsäde och certifikatutsäde, förutom då utsäde av den sistnämnda kategorin förpackas i EEG-småförpackningar..."
5. Texten i artikel 11.2 b skall ersättas med följande:
"b) anta bestämmelser om undantag från punkt 1 för småförpackningar med basutsäde om dessa är märkta med: "Endast godkänt för saluföring i . . . . . . (den berörda medlemsstaten)"."
6. Följande artiklar skall läggas till efter artikel 11:
Obligatoriska uppgifter 1. "EEG-småförpackning".
RÅDETS FÖRORDNING (EEG) nr 2777/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för fjäderfäkött
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 42 och 43 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1), och
med beaktande av följande. De grundläggande bestämmelserna om organisationen av marknaden för fjäderfäkött har ändrats ett flertal gånger sedan de antogs. Eftersom bestämmelserna är många och komplicerade och dessutom återfinns i ett antal olika nummer av Europeiska gemenskapernas officiella tidning, är de svåra att tillämpa och saknar följaktligen den klarhet som bör vara ett väsentligt drag i all lagstiftning. De bör därför sammanföras i en enda text.
För att den gemensamma marknaden för jordbruksprodukter skall kunna fungera och utvecklas måste den kompletteras av en gemensam jordbrukspolitik som framför allt innefattar gemensam organisation av marknaderna för olika jordbruksprodukter. En sådan organisation kan utformas på olika sätt beroende på vilket produkt det är fråga om.
Syftet med den gemensamma jordbrukspolitiken är att uppnå de mål som fastställs i artikel 39 i fördraget. För att stabilisera marknaderna och tillförsäkra den berörda jordbruksbefolkningen en skälig levnadsstandard bör det inom fjäderfäköttsektorn införas bestämmelser om åtgärder för att underlätta anpassningen av utbudet till marknadens behov.
Förverkligandet av en enhetlig marknad för fjäderfäkött inbegriper införandet av ett enhetligt system för handeln över gemenskapens yttre gränser, innefattande importavgifter och exportbidrag.
För att uppnå detta syfte bör det i regel vara tillräckligt att i samband med import från tredje land införa importavgifter som bestäms med hänsyn till effekten på foderkostnaderna av den skillnad som råder mellan priserna på foderspannmål inom gemenskapen och på världsmarknaden, och till behovet att skydda gemenskapens förädlingsindustri.
Det är nödvändigt att undvika störningar på gemenskapsmarknaden till följd av utbud på världsmarknaden till extremt låga priser. Därför bör slusspriser fastställas och om anbudspriserna fritt gränsen är lägre än slusspriserna bör importavgifterna höjas med en tilläggsavgift.
Gemenskapens deltagande i den internationella handeln med fjäderfäkött skulle säkras av möjligheten att vid export till tredje land bevilja ett exportbidrag som motsvarar skillnaden mellan priserna inom gemenskapen och priserna på världsmarknaden. För att garantera gemenskapens exportörer ett visst mått av trygghet med avseende på exportbidragens stabilitet, bör det göras möjligt att fastställa exportbidraget för fjäderfäkött på förhand.
Utöver det ovan beskrivna systemet bör möjligheter skapas att, när marknadssituationen så kräver, helt eller delvis förbjuda tillämpningen av aktiv förädling.
Beviljandet av vissa former av stöd kan äventyra förverkligandet av en enhetlig marknad. Följaktligen bör de bestämmelser i fördraget som gör det möjligt att värdera stödåtgärder som beviljats av medlemsstaterna och att förbjuda stödåtgärder som är oförenliga med den gemensamma marknaden göras tillämpliga på marknaden för fjäderfä.
Den gemensamma organisationen av marknaden för fjäderfäkött skall på lämpligt sätt och samtidigt ta hänsyn till de mål som fastställs i artikel 39 och artikel 110 i fördraget.
De utgifter som medlemsstaterna ådrar sig till följd av förpliktelser som uppstår vid tillämpningen av denna förordning skall finansieras av gemenskapen i enlighet med bestämmelserna i artikel 2 och 3 i rådets förordning (EEG) nr 729/70(2) av den 21 april 1970 om finansieringen av den gemensamma jordbrukspolitiken, ändrad genom förordning (EEG) nr 1566/72(3).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. I denna förordning avses med: a) levande fjäderfä: levande höns, ankor, gäss, kalkoner och pärlhöns med en vikt på över 185 gram.
b) kycklingar: levande höns, ankor, gäss, kalkoner och pärlhöns med en högsta vikt på 185 gram.
c) slaktade fjäderfä: döda höns, ankor, gäss, kalkoner och pärlhöns, hela och med eller utan slaktbiprodukter.
d) härledda produkter: 1. produkter enligt punkt 1 a utom kycklingar.
2. produkter enligt punkt 1 b utom slaktade fjäderfä och ätbara slaktbiprodukter så kallade styckningsdelar av fjäderfä,
3. ätbara slaktbiprodukter enligt punkt 1 b,
4. produkter enligt punkt 1 c,
5. produkter enligt punkt 1 d och e,
6. produkter enligt punkt 1 f.
e) kvartal: tremånadersperiod som börjar den 1 februari, den 1 maj, den 1 augusti eller den 1 november.
Artikel 2
- Åtgärder för att förbättra kvaliteten.
- Åtgärder för att möjliggöra kort- och långsiktiga prognoser på grundval av de produktionsmedel som används.
- Åtgärder för att underlätta registreringen av prisutvecklingen på marknaden.
Allmänna bestämmelser om dessa åtgärder skall antas i enlighet med det förfarande som föreskrivs i artikel 43.2 i fördraget.
2. Handelsnormer - skall antas för en eller flera av de produkter som anges i artikel 1.1 b,
- får antas för de produkter som anges i artikel 1.1 a, c, d, e och f.
Dessa normer får särskilt avse klassificering efter kvalitet och vikt, förpackning, lagring, transport, presentation och märkning.
På förslag av kommissionen skall rådet med kvalificerad majoritet fastställa normerna och deras användningsområde samt allmänna tillämpningsföreskrifter för dem.
Artikel 3
De produkter som anges i artikel 1.1 skall vid import till gemenskapen beläggas med en importavgift som fastställs på förhand för varje kvartal i enlighet med det förfarande som föreskrivs i artikel 17.
Artikel 4
1. Importavgiften på slaktat fjäderfä skall bestå av följande delar: a) En del som motsvarar skillnaden mellan gemenskapens och världsmarknadens priser på den kvantitet fodersäd, differentierad med hänsyn till art av fjäderfä, som åtgår till att inom gemenskapen producera 1 kg slaktat fjäderfä.
Priserna på foderspannmål inom gemenskapen skall fastställas en gång om året för en tolvmånadersperiod som börjar den 1 augusti. Dessa priser skall baseras på tröskelpriserna på sådan spannmål och den månatliga höjningen av dessa priser.
Världsmarknadspriserna på foderspannmål skall fastställas kvartalsvis på basis av priserna på sådan spannmål under de sex månader som föregår det kvartal under vilket nämnda del beräknas.
Vid fastställande av de importavgifter som skall tillämpas från och med den 1 november, den 1 februari och den 1 maj, skall emellertid hänsyn tas till utvecklingen av världsmarknadspriserna på foderspannmål endast om ett nytt slusspris fastställs samtidigt.
2. Importavgiften för kycklingar skall beräknas på samma sätt som importavgiften för slaktat fjäderfä. Dock skall den kvantitet foderspannmål som skall användas vid beräkningen vara den kvantitet som åtgår till att inom gemenskapen producera en kyckling. Slusspriset skall vara det som gäller för kycklingar.
3. På förslag av kommissionen skall rådet med kvalificerad majoritet - fastställa den kvantitet foderspannmål, differentierad med hänsyn till art av fjäderfä, som åtgår till att producera 1 kg slaktat fjäderfä och den kvantitet foderspannmål som åtgår till att producera en kyckling, samt procentsatserna av de olika slag av foderspannmål som ingår i dessa kvantiteter,
- anta tillämpningsföreskrifter för denna artikel.
Artikel 5
1. För de produkter som anges i artikel 1.2 d skall importavgiften härledas från importavgiften för slaktat fjäderfä, på basis av viktförhållandet mellan dessa olika produkter och slaktat fjäderfä och, vid behov, det genomsnittliga förhållandet mellan deras marknadsvärden.
2. Trots bestämmelserna i punkt 1 skall importavgiften för de produkter som anges under Gemensamma tulltaxans nummer 02.03, 15.01 B och 16.02 B I och för vilka tullsatsen har bundits inom GATT, begränsas till det belopp som följer av denna bundenhet.
3. Koefficienterna som uttrycker de förhållanden som avses i punkt 1 skall fastställas i enlighet med det förfarande som föreskrivs i artikel 17. De uppgifter som används vid fastställande av koefficienterna skall omprövas minst en gång om året.
Artikel 6
Om en betydande prisökning noteras på gemenskapsmarknaden och denna situation sannolikt kommer att bestå och därigenom stör eller hotar att störa marknaden, får nödvändiga åtgärder vidtas.
Rådet skall på förslag av kommissionen och med kvalificerad majoritet anta allmänna tillämpningsföreskrifter för denna artikel.
Artikel 7
1. Slusspriserna skall fastställas på förhand för varje kvartal i enlighet med artikel 17.
2. Slusspriserna på slaktat fjäderfä skall utgöras av följande delar: a) Ett belopp som motsvarar världsmarknadspriset på den kvantitet foderspannmål, differentierad med hänsyn till art av fjäderfä, som åtgår till att i tredje land producera 1 kg slaktat fjäderfä.
b) Ett standardbelopp som representerar övriga foderkostnader och omkostnader för produktion och försäljning, differentierad med hänsyn till art av fjäderfä.
Världsmarknadspriset på kvantiteten av foderspannmål skall fastställas kvartalsvis på basis av priserna på sådan spannmål under de sex månader som föregår det kvartal under vilket slusspriset fastställs.
Vid fastställande av det slusspris som skall gälla från den 1 november, den 1 februari och den 1 maj skall emellertid hänsyn tas till prisutvecklingen på världsmarknaden för foderspannmål endast om priset på kvantiteten foderspannmål uppvisar en minimiavvikelse från det pris som användes vid beräkning av slusspriset för föregående kvartal. De uppgifter som används för att fastställa det standardbelopp som avses i b skall omprövas minst en gång om året.
3. Slusspriset på kycklingar skall beräknas på samma sätt som slusspriset på slaktat fjäderfä. Dock skall världsmarknadspriset på kvantiteten foderspannmål vara priset på den kvantitet som åtgår till att i tredje land producera en kyckling och standardbeloppet skall vara det belopp som representerar övriga foderkostnader och omkostnader för produktion och försäljning för en kyckling. Mängden foderspannmål och standardbeloppet skall inte variera beroende på art.
4. För de produkter som anges i artikel 1.2 d skall slusspriserna härledas från slusspriset på slaktat fjäderfä på basis av de koefficienter som fastställts för sådana produkter i enlighet med artikel 5.3.
5. Rådet skall på förslag av kommissionen och med kvalificerad majoritet anta tillämpningsföreskrifter för denna artikel.
Artikel 8
1. Om anbudspriset fritt gränsen för en produkt ligger under slusspriset, skall importavgiften för denna vara höjas med en tilläggsavgift som motsvarar skillnaden mellan slusspriset och anbudspriset fritt gränsen.
2. Importavgiften skall emellertid inte höjas med denna tilläggsavgift när det gäller tredje land som vill och är i stånd att garantera att importpriset till gemenskapen på produkter som har sitt ursprung i och kommer från deras territorium inte kommer att bli lägre än slusspriset för produkten i fråga och att varje snedvridning av handeln kommer att undvikas.
3. Anbudspriset fritt gränsen skall fastställas för all import från tredje land.
Om exporten från ett eller flera tredje länder sker till onormalt låga priser, lägre än de priser som gäller i andra tredje länder, skall ett andra anbudspris fritt gränsen fastställas för export från dessa länder.
4. Närmare tillämpningsföreskrifter för denna artikel skall antas i enlighet med förfarandet i artikel 17.
Då tilläggsavgifter krävs, skall dessa fastställas i enlighet med samma förfarande.
Artikel 9
1. I den mån det är nödvändigt för att göra det möjligt att exportera de produkter som avses i artikel 1.1 på grundval av världsmarknadspriserna på dessa produkter, får skillnaden mellan världsmarknadspriserna och priserna inom gemenskapen täckas av ett exportbidrag.
2. Exportbidraget skall vara detsamma för hela gemenskapen. Det får variera beroende på användning och bestämmande.
Exportbidraget skall beviljas på ansökan av berörd part.
Vid fastställande av exportbidraget skall särskild hänsyn tas till behovet av att skapa en balans mellan användningen av gemenskapens basvaror vid framställningen av bearbetade varor för export till tredje land och användningen av produkter från tredje land som förts in enligt bestämmelserna för aktiv förädling.
På förslag av kommissionen skall rådet med kvalificerad majoritet fastställa allmänna bestämmelser om beviljande av och förutfastställelse av exportbidrag och kriterier för fastställande av dessa belopp.
Exportbidrag skall fastställas med jämna mellanrum i enlighet med förfarandet i artikel 17. Vid behov får kommissionen, på begäran av en medlemsstat eller på eget initiativ, ändra exportbidragen under mellanperioderna.
3. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 17.
Artikel 10
I den mån det är nödvändigt för att den gemensamma organisation av marknaden för fjäderfäkött skall fungera väl, får rådet, på förslag av kommissionen, med kvalificerad majoritet helt eller delvis förbjuda tillämpningen av bestämmelserna för aktiv förädling för produkter enligt artikel 1.1 som skall användas till framställningen av de produkter som anges i den punkten.
Artikel 11
1. De allmänna bestämmelserna om tolkningen av Gemensamma tulltaxan och de särskilda tillämpningsföreskrifterna skall gälla tullklassificeringen av produkter som omfattas av denna förordning. Tullnomenklaturen som skapas genom tillämpningen av denna förordning skall ingå som del i Gemensamma tulltaxan.
2. Såvida inte annat föreskrivs i denna förordning eller rådet, på förslag av kommissionen, med kvalificerad majoritet fattar beslut om undantag från denna förordning, skall följande vara förbjudet:
- Införande av tullar eller avgifter med motsvarande verkan.
- Tillämpning av någon kvantitativ restriktion eller åtgärd med motsvarande verkan. Varje åtgärd som begränsar utfärdandet av import- eller exportlicenser till en angiven personkategori skall betraktas som en åtgärd som har samma verkan som en kvantitativ restriktion.
Artikel 12
1. Om gemenskapsmarknaden för en eller flera av de produkter som anges i artikel 1.1, till följd av import eller export är utsatt för eller hotas av allvarliga störningar som kan äventyra de mål som fastställs i artikel 39 i fördraget, får lämpliga åtgärder avseende handeln med tredje land vidtas till dess att störningen eller hotet om störning har upphört.
På förslag av kommissionen skall rådet med kvalificerad majoritet fastställa närmare tillämpningsföreskrifter för denna punkt samt närmare ange under vilka omständigheter och inom vilka gränser medlemsstaterna får vidta skyddsåtgärder.
2. Om den situation som avses i punkt 1 uppstår skall kommissionen, på begäran av en medlemsstat eller på eget initiativ, fatta beslut om nödvändiga åtgärder. Medlemsstaterna skall underrättas om beslutet som skall gälla med omedelbar verkan. Om kommissionen mottar en begäran från en medlemsstat, skall den fatta beslut om denna begäran inom 24 timmar efter det att den mottagits.
3. En medlemsstat får hänskjuta kommissionens beslut om åtgärder till rådet inom tre arbetsdagar efter det att beslutet meddelades. Rådet skall sammanträda utan dröjsmål och får med kvalificerad majoritet ändra eller upphäva åtgärderna i fråga.
Artikel 13
De produkter som anges i artikel 1.1 och som framställs av eller utvinns ur produkter som inte är angivna i artikel 9.2 och 10.1 i fördraget skall inte få omsättas fritt inom gemenskapen.
Artikel 14
För att ta hänsyn till eventuella begränsningar av den fria omsättningen till följd av åtgärder för att förhindra spridning av djursjukdomar, får extraordinära åtgärder för att stödja marknader som påverkas av sådana begränsningar vidtas i enlighet med det förfarande som föreskrivs i artikel 17. Sådana åtgärder får endast vidtas i den mån och under den tid som det är absolut nödvändigt för att stödja denna marknad.
Artikel 15
Medlemsstaterna och kommissionen skall till varandra överlämna sådana uppgifter som är nödvändiga för att tillämpa denna förordning. Bestämmelser om överlämnande och spridning av sådana uppgifter skall fastställas i enlighet med det förfarande som föreskrivs i artikel 17.
Artikel 16
1. Härmed inrättas en förvaltningskommitté för fjäderfäkött och ägg (nedan kallad "kommittén"). Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
2. Inom kommittén skall medlemsstaternas röster vägas enligt artikel 148.2 i fördraget. Ordföranden får inte rösta.
Artikel 17
1. När förfarandet som föreskrivs i denna artikel skall tillämpas, skall ordföranden hänskjuta ärendet till kommittén, antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med en majoritet av 41 röster.
3. Kommissionen skall besluta med omedelbar verkan. Om beslutet inte är förenligt med kommitténs yttrande skall kommissionen emellertid genast underrätta rådet. I sådana fall får kommissionen uppskjuta verkställandet av de beslutade åtgärderna under en tid som inte överstiger en månad från dagen då rådet underrättats.
Rådet får inom en månad fatta ett annat beslut med kvalificerad majoritet.
Artikel 18
Kommittén får överväga varje annan fråga som dess ordförande hänskjuter till kommittén på eget initiativ eller på begäran av en medlemsstats företrädare.
Artikel 19
Om inte annat följer av denna förordning, skall artikel 92 94 i fördraget gälla för produktionen av och handeln med de produkter som anges i artikel 1.1.
Artikel 20
Denna förordning skall tillämpas så att hänsyn tas samtidigt och på lämpligt sätt till de mål som fastställs i artiklarna 39 och 110 i fördraget.
Artikel 21
Om Italien åberopar bestämmelserna i artikel 23 i rådets förordning (EEG) nr 2727/75(4) av den 29 oktober 1975 om den gemensamma organisationen av marknaden för spannmål, skall rådet, på förslag av kommissionen, med kvalificerad majoritet besluta om de åtgärder som krävs för att undvika en snedvridning av konkurrensen.
Artikel 22
1. Rådets förordning nr 123/67/EEG(5) av den 13 juni 1967 om den gemensamma organisationen av marknaden för fjäderfäkött, senast ändrad genom rådets beslut av den 1 januari 1973(6) om anpassning av dokumenten avseende de nya medlemsstaternas anslutning till Europeiska gemenskaperna, upphävs härmed.
2. Alla hänvisningar till den förordning som upphävs i punkt 1 skall betraktas som hänvisningar till den här förordningen.
Hänvisningar till artiklar i den upphävda förordningen skall läsas enligt den jämförelsetabell som finns i bilagan.
Artikel 23
Denna förordning träder i kraft den 1 november 1975.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: De tekniska krav som motorfordon måste uppfylla enligt nationell lagstiftning gäller bl.a. föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt.
Dessa krav skiljer sig åt från en medlemsstat till en annan. Det är därför nödvändigt att alla medlemsstater antar samma krav, antingen som tillägg till eller i stället för sina nuvarande regler, för att därmed för alla fordonstyper medge det förfarande för EEG-typgodkännande som behandlats i rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(3).
Tillnärmningen av den nationella lagstiftningen om motorfordon innefattar medlemsstaternas ömsesidiga erkännande av de kontroller som utförs av var och en av dem på grundval av gemensamma bestämmelser. För att ett sådant system skall bli framgångsrikt måste dessa bestämmelser tillämpas av alla medlemsstater från samma datum.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I detta direktiv avses med fordon varje motorfordon som är avsett att användas på väg, med eller utan karosseri, med minst fyra hjul och som är konstruerade för en högsta hastighet som överstiger 25 km/tim och släpvagnar till dessa fordon, dock med undantag av spårbundna fordon, traktorer och maskiner för jordbruk eller skogsbruk samt andra motorredskap.
Artikel 2
Ingen medlemsstat får vägra att bevilja EEG-typgodkännande eller nationellt typgodkännande för ett fordon av skäl som hänför sig till de föreskrivna skyltarna och märkningarna eller deras placering och fastsättningsmetod om de uppfyller kraven i bilagan.
Artikel 3
Ingen medlemsstat får vägra att registrera ett fordon eller förbjuda att det säljs, tas i bruk eller används av skäl som hänför sig till de föreskrivna skyltarna och märkningarna eller deras placering och fastsättningsmetod om de uppfyller kraven i bilagan till detta direktiv.
Artikel 4
De ändringar som är nödvändiga för att anpassa kraven i bilagan till den tekniska utvecklingen skall antas enligt det förfarande som beskrivs i artikel 13 i direktiv 70/156/EEG.
Artikel 5
2. Efter anmälan av detta direktiv skall medlemsstaterna underrätta kommissionen om alla förslag till lagar och andra författningar som de avser att anta inom det område som omfattas av detta direktiv; underrättelsen skall lämnas i så god tid att kommissionen hinner lämna synpunkter på förslaget.
Artikel 6
RÅDETS DIREKTIV av den 8 december 1975 om kvaliteten på badvatten (76/160/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 100 och 235 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: För att skydda miljön och människors hälsa är det nödvändigt att minska föroreningen av badvatten och att skydda sådant vatten mot ytterligare försämring.
Kontroll av badvatten är nödvändig för att inom ramen för den gemensamma marknaden uppnå gemenskapens mål vad avser en förbättring av levnadsvillkoren, en harmonisk utveckling av ekonomiska verksamheter inom gemenskapen som helhet och en fortgående och balanserad tillväxt.
Inom detta område finns det vissa lagar och andra författningar i medlemsstaterna som direkt påverkar den gemensammamarknadens funktion. Fördraget ger dock inte alla de befogenheter som är nödvändiga för att vidta åtgärder.
Enligt Europeiska gemenskapernas åtgärdsprogram för miljön(3) skall gemensamma kvalitetsmål uppställas med avseende på miljökvaliteten, bl.a. angivande av parametervärden för vatten, inklusive badvatten.
För att uppnå dessa kvalitetsmål måste medlemsstaterna fastställa gränsvärden enligt vissa parametrar. Badvatten måste överensstämma med dessa värden inom tio år efter anmälan av detta direktiv.
Det bör föreskrivas att badvatten under vissa förhållanden skall anses uppfylla de relevanta parametervärdena, även om en viss procent av proven som tagits under badsäsongen inte överensstämmer med de gränsvärden som anges i bilagan.
För att uppnå ett visst mått av flexibilitet vid tillämpningen av detta direktiv måste medlemsstaterna ha befogenhet att föreskriva undantag. Sådana undantag får emellertid inte bortse från krav som är väsentliga för skyddet av människors hälsa.
Den tekniska utvecklingen gör det nödvändigt med en snabb anpassning av de tekniska krav som fastställs i bilagan. För att underlätta beslut om de åtgärder som krävs för detta ändamål, bör ett förfarande fastställas genom vilket ett nära samarbete upprättas mellan medlemsstaterna och kommissionen inom en kommitté för anpassning till den tekniska utvecklingen.
Allmänhetens intresse för miljön och en förbättrad miljökvalitet ökar. Allmänheten bör därför få objektiv information om kvaliteten på badvatten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) "badvatten": allt rinnande eller stillastående sötvatten och havsvatten, i vilket - badning är uttryckligen tillåten av de behöriga myndigheterna i varje medlemsstat, eller
- badning inte är förbjuden och traditionellt utövas av ett stort antal badare,
b) "badplats": varje plats där badvatten finns,
c) "badsäsong": den period under vilken ett stort antal badare kan förutses med hänsyn till lokalt bruk, inbegripet eventuella lokala regler för badning och väderleksförhållanden.
Artikel 2
Fysikaliska, kemiska och mikrobiologiska parametrar som gäller för badvatten anges i bilagan, som utgör en integrerad del av detta direktiv.
Artikel 3
1. Medlemsstaterna skall för alla badplatser eller för varje enskild badplats fastställa de värden som skall gälla för badvatten i fråga om de parametrar som anges i bilagan.
Artikel 4
Kommissionen får delta i dessa överläggningar.
Artikel 5
- i 90 % av proverna i alla andra fall med undantag av parametrarna för "kolibakterier, totalt" och "fekala kolibakterier" där procentsatsen får vara 80 %,
och om, i fråga om de 5, 10 eller 20 % av proven som inte överensstämmer med värdena
- vattnet inte avviker från de relevanta parametervärdena med mer än 50 % utom för mikrobiologiska parametrar, pH och löst syre,
Artikel 6
Artikel 7
Artikel 8
Bestämmelserna i detta direktiv får åsidosättas a) i fråga om vissa parametrar märkta (0) i bilagan vid exceptionella meteorologiska eller geografiska förhållanden,
b) om badvatten berikas på naturlig väg med vissa ämnen och detta orsakar avvikelse från de värden som föreskrivs i bilagan.
Naturlig berikning avser den process genom vilken en viss vattenmassa, utan mänsklig påverkan, tillförs vissa ämnen ur marken.
De undantag som föreskrivs i denna artikel får inte i något fall medföra att krav som är väsentliga för att skydda människors hälsa åsidosätts.
Om en medlemsstat åsidosätter bestämmelserna i detta direktiv skall den omedelbart meddela kommissionen detta med uppgift om skälen och den förväntade tidsperioden.
Artikel 9
Sådana ändringar som är nödvändiga för att anpassa detta direktiv till den tekniska utvecklingen skall avse - analysmetoderna,
- de G- och I-parametervärden som anges i bilagan.
De skall antas i enlighet med det förfarande som fastställs i artikel 11.
Artikel 10
Artikel 11
3. a) Kommissionen skall själv anta förslaget om det är förenligt med kommitténs yttrande.
b) Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
c) Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 12
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv inom två år efter dagen för anmälan. De skall genast underrätta kommissionen om detta.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 13
Medlemsstaterna skall fyra år efter anmälan av detta direktiv och därefter regelbundet till kommissionen överlämna en utförlig rapport om sitt badvatten och dess mest betydelsefulla egenskaper.
Kommissionen kan offentliggöra den erhållna informationen efter det att den berörda medlemsstaten har gett sitt tillstånd.
Artikel 14
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 27 juli 1976 om tillnärmning av medlemsstaternas lagstiftning om alkoholmätare och alkoholaerometrar (76/765/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: Definition, konstruktion och metoder för godkännande och provning av alkoholmätare och alkoholaerometrar är i medlemsstaterna underkastade tvingande bestämmelser som skiljer sig mellan medlemsstaterna och därmed utgör hinder för rörligheten av och handeln med dessa mätdon inom gemenskapen. Dessa bestämmelser måste därför närmas till varandra.
Harmonisering av lagar och andra författningar som avser dessa mätdon är också väsentlig som ett komplement till gällande bestämmelser om metoder att bestämma alkoholhalt utgående från mätresultat, så att alla risker avlägsnas för flertydighet i eller ifrågasättande av resultaten av sådana mätningar.
Rådets direktiv 71/316/EEG av den 26 juli 1971 om tillnärmning av medlemsstaternas lagstiftning om gemensamma föreskrifter för både mätdon och metrologiska kontrollmetoder(3) har fastställt förfaranden för EEG-typgodkännande och första EEG-verifikation. Enligt det direktivet är det nödvändigt att fastställa de tekniska krav som skall gälla för konstruktion och funktion av alkoholmätare och alkoholaerometrar för att de efter föreskriven kontroll och märkning fritt skall få importeras, marknadsföras och användas.
I sin resolution av den 17 december 1973(4) om industripolitik uppmanade rådet kommissionen att före den 1 december 1974 till rådet lämna ett förslag till ett direktiv om alkoholmätning och alkoholmätare.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Detta direktiv fastställer egenskaper hos alkoholmätare och alkoholaerometrar som används för att bestämma alkoholhalten i blandningar av vatten och etanol.
Artikel 2
Artikel 3
Ingen medlemsstat får begränsa, vägra eller förbjuda att någon alkoholmätare eller alkoholaerometer släpps ut på marknaden eller tas i drift, under åberopande av dess metrologiska egenskaper, om den försetts med märkning för EEG-typgodkännande eller första EEG-verifikation.
Artikel 4
Bestämmelserna skall börja tillämpas senast den 1 januari 1980.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 16 december 1976 om minimikrav på utbildning av vissa förare av vägfordon (76/914/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 75 i detta,
med beaktande av rådets förordning (EEG) nr 543/69 av den 25 mars 1969 om harmonisering av viss social lagstiftning rörande transporter på väg(), senast ändrad genom förordning (EEG) nr 515/72(), och särskilt artikel 5.1 b andra strecksatsen och artikel 2 c i denna,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(),
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
med beaktande av följande: I artikel 5.1 b andra strecksatsen i förordning (EEG) nr 543/69 föreskrivs att förare av ett fordon som är avsett för transport av gods med en högsta tillåtna vikt över 7,5 metriska ton och som omfattas av förordningen, måste, om vederbörande inte har fyllt 21 år, inneha ett intyg om yrkeskompetens som är erkänt i en av medlemsstaterna. Intyget skall styrka att föraren har genomgått utbildning för förare av fordon som är avsedda för godstransporter på väg.
Vid fastställande av miniminivån för sådan utbildning bör man särskilt ta hänsyn till de olika förutsättningar som råder för gods- respektive persontransporter på väg.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Den som innehar gällande nationellt körkort och som har genomgått yrkesutbildning som omfattar åtminstone de ämnen som är uppräknade i bilagan till detta direktiv, skall anses ha uppfyllt minimikravet på utbildning för förare av fordon avsedda för godstransporter på väg enligt artikel 5.1 b andra strecksatsen i förordning (EEG) nr 543/69 eller för förare av fordon avsedda för persontransporter på väg enligt punkt 2 c av nämnda artikel.
2. Kursinnehåll och uppläggning i fråga om den yrkesutbildning som avses i punkt 1 skall fastställas av medlemsstaten. Att sådan utbildning har genomgåtts skall styrkas genom examen eller kunskapskontroll som ombesörjs av staten eller av de organ som staten har utsett att utföra kontrollen under direkt överinseende av staten.
3. Varje medlemsstat får kräva att förare som utför inrikestransporter på dess territorium och förare som utför internationella transporter med fordon registrerade i denna stat skall genomgå en mer omfattande utbildning än den som beskrivs i bilagan. Denna utbildning kan utgöras av utbildning som redan finns eller av utbildning som en medlemsstat beslutar införa i framtiden.
Artikel 2
1. Det intyg om yrkeskompetens som avses i andra strecksatsen i artikel 5.1 b och artikel 5.2 c i förordning (EEG) nr 543/69 skall utfärdas till de personer som uppfyller de villkor som föreskrivs i artikel 1 i detta direktiv av den stat eller av de organ som staten utsett att ombesörja utfärdandet under direkt överinseende av staten.
2. Rättigheter som förvärvats med stöd av de föreskrifter som avses i punkt 1 innan de nationella lagar och andra författningar som har antagits till följd av detta direktiv träder i kraft, skall förbli giltiga på samma sätt som utbildningsintyg, som utfärdats enligt detta direktiv.
Artikel 3
1. Efter samråd med kommissionen skall medlemsstaterna inom två år efter anmälan av detta direktiv genomföra de åtgärder som är nödvändiga för att följa direktivet.
2. Varje medlemsstat skall tillställa kommissionen prov på de utbildningsintyg eller likvärdiga dokument som staten inför för tillämpning av artikel 2.1. Kommissionen skall snarast vidarebefordra dessa underlag till de övriga medlemsstaterna.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EEG) nr 2566/76 av den 20 juli 1976 om godkännande av avtalet i form av skriftväxling rörande ändringar i tabell I och II i bilaga till protokoll 2 till avtalet mellan Europeiska ekonomiska gemenskapen och Schweiz
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 113 i detta,
med beaktande av kommissionens rekommendation, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Härmed godkänns på gemenskapens vägnar avtalet i form av skriftväxling om ändringar i tabell I och II i bilaga till protokoll 2 till avtalet mellan Europeiska ekonomiska gemenskapen och Schweiz.
Avtalets text ingår i bilaga till denna förordning.
Artikel 2
Rådets ordförande bemyndigas att utse den person som är behörig att med bindande verkan för gemenskapen underteckna avtalet.
Artikel 3
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS ANDRA DIREKTIV av den 13 december 1976 om samordning av de skyddsåtgärder som krävs i medlemsstaterna av de i artikel 58 andra stycket i fördraget avsedda bolagen i bolagsmännens och tredje mans intressen när det gäller att bilda ett aktiebolag samt att bevara och ändra dettas kapital, i syfte att göra skyddsåtgärderna likvärdiga (77/91/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 54.3 g i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
med beaktande av följande: Eftersom aktiebolagen spelar en framträdande roll i medlemsstaternas näringsliv och deras verksamhet ofta sträcker sig utöver de nationella gränserna, är det i fråga om dessa bolag särskilt viktigt att fortsätta den samordning som föreskrivs i artikel 54.3 g i fördraget och i Allmänna handlingsprogrammet för upphävande av begränsningar av etableringsfriheten och som inleddes med direktiv 68/151/EEG (3).
För att aktieägarna och borgenärerna skall kunna garanteras ett minimum av likvärdigt skydd är det särskilt viktigt att samordna de nationella bestämmelserna om att bilda ett aktiebolag samt om att bevara, öka och sätta ned dess kapital.
Inom gemenskapen måste ett aktiebolags bolagsordning eller stiftelseurkund utformas på ett sådant sätt att varje intressent ur dessa handlingar kan inhämta grundläggande uppgifter om bolaget, däribland en detaljerad redovisning av kapitalets sammansättning.
Sådana gemenskapsregler om att bevara det kapital som utgör borgenärernas säkerhet skall antas, som särskilt förbjuder en minskning av kapitalet genom utdelning till aktieägarna och begränsar bolagens möjligheter att förvärva egna aktier.
Med hänsyn till ändamålet med artikel 54.3 i fördraget måste medlemsstaternas lagstiftning om ökning och nedsättning av kapitalet säkerställa att de principer beaktas och harmoniseras som syftar till en lika behandling av aktieägare med samma ställning och till ett skydd för borgenärer med fordringar som har uppkommit före en kapitalnedsättning,
HÄRIGENOM FÖRESKRIVS FÖLJANDE
Artikel 1
1. De samordningsåtgärder som detta direktiv föreskriver skall vidtas i fråga om bestämmelserna i medlemsstaternas lagar eller andra författningar om följande bolagsformer: - I Belgien: la société anonyme/de naamloze vennootschap.
- I Danmark: aktieselskabet.
- I Italien: la società per azioni.
2. Medlemsstaterna behöver inte tillämpa detta direktiv på förvaltningsbolag med rörligt kapital eller på kooperativa företag som är organiserade i någon av de i punkt 1 angivna bolagsformerna. Om lagstiftningen i en medlemsstat utnyttjar denna möjlighet, skall den föreskriva att dessa bolag skall ta in orden "förvaltningsbolag med rörligt kapital" eller "kooperativt företag" i samtliga de handlingar som nämns i artikel 4 i direktiv 68/151/EEG.
Med "förvaltningsbolag med rörligt kapital" avses i detta direktiv endast bolag - som uteslutande har till föremål för sin verksamhet att placera sina medel i olika värdepapper, fastigheter eller andra tillgångar med enda syfte att sprida investeringsriskerna och fördela resultatet av kapitalförvaltningen mellan aktieägarna,
- som inbjuder allmänheten att förvärva aktier i bolaget, och
- vars bolagsordning anger att bolaget inom gränserna för ett minimikapital och ett maximikapital alltid får ge ut, lösa in eller avyttra sina aktier.
Artikel 2
Bolagsordningen eller stiftelseurkunden skall alltid innehålla minst följande uppgifter: a) bolagsform och firma;
b) föremålet för bolagets verksamhet;
c) - om bolaget inte har något "auktoriserat" kapital, det tecknade kapitalets storlek;
- om bolaget har ett "auktoriserat" kapital, storleken av detta och det tecknade kapitalet vid bolagsbildningen eller då bolaget får tillstånd att börja sin verksamhet och vid varje ändring av det "auktoriserade" kapitalet, dock med förbehåll för vad som gäller enligt artikel 2.1 e i direktiv 68/151/EEG;
d) bestämmelser som anger antalet ledamöter och hur dessa skall utses i de organ som företräder bolaget mot tredje man och svarar för förvaltning, ledning, övervakning eller kontroll av bolaget samt bestämmelser om kompetensfördelningen mellan organen, allt i den mån föreskrifter inte finns i lag eller annan författning;
e) tiden för bolagets bestånd om inte denna tid är obestämd.
Artikel 3
Minst följande uppgifter skall finnas antingen i bolagsordningen eller stiftelseurkunden eller i en särskild handling som skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG: a) bolagets säte;
b) de tecknade aktiernas nominella belopp och, minst en gång om året, deras antal;
c) antalet tecknade aktier utan nominellt belopp, om den nationella lagstiftningen tillåter att sådana aktier ges ut;
d) i förekommande fall de särskilda villkor som begränsar aktiernas överlåtbarhet;
e) om det finns aktier av olika slag, uppgifter enligt b, c och d för varje aktieslag med uppgift om de rättigheter som är förenade med varje aktieslag;
f) huruvida aktierna är ställda till viss man eller till innehavaren, om den nationella lagstiftningen tillåter båda formerna, och bestämmelser om hur aktierna omvandlas från den ena formen till den andra, om inte förfarandet är reglerat i lag eller annan författning;
g) hur stor del av det tecknade kapitalet som är betalt då bolaget bildas eller då det får tillstånd att börja sin verksamhet;
h) det nominella värdet av de aktier eller, i avsaknad av sådant värde, det antal aktier som ges ut mot tillskott av annan egendom än pengar (apportegendom) samt beskrivning av denna egendom och namnet på den som tillskjuter egendomen;
i) identiteten hos de fysiska eller juridiska personer eller bolag av vilka eller i vilkas namn bolagsordningen eller stiftelseurkunden eller, om bolagsbildningen inte sker i ett sammanhang, utkasten till dessa handlingar har undertecknats;
j) åtminstone uppskattningsvis summan av alla kostnader som har uppkommit för bolaget eller påförts detta med anledning av bolagsbildningen och, i förekommande fall, innan bolaget får tillstånd att börja sin verksamhet;
k) särskilda förmåner som vid bolagsbildningen eller före tillståndet att börja verksamheten har tillerkänts någon som har deltagit i bolagsbildningen eller i åtgärder som har lett fram till tillståndet.
Artikel 4
1. Om enligt lagstiftningen i en medlemsstat ett bolag inte får börja sin verksamhet utan tillstånd, skall denna lagstiftning även innehålla bestämmelser om ansvaret för förbindelser som har ingåtts av bolaget eller för dettas räkning innan ansökningen om tillstånd beviljades eller avslogs.
2. Punkt 1 tillämpas inte på förbindelser med anledning av avtal som bolaget har ingått på villkor att det får tillstånd att börja sin verksamhet.
Artikel 5
1. Om lagstiftningen i en medlemsstat kräver att ett bolag skall bildas av flera bolagsmän, medför inte det förhållandet att därefter alla aktierna förenas på en hand eller antalet bolagsmän sjunker under det i lagstiftningen föreskrivna minimiantalet att bolaget utan vidare upplöses.
2. Om enligt lagstiftningen i en medlemsstat ett bolag i fall som avses i punkt 1 kan upplösas genom förordnande av rätten, får behörig domstol ge bolaget den frist som detta behöver för att vidta rättelse.
3. När förordnandet om upplösning har meddelats, skall bolaget träda i likvidation.
Artikel 6
1. Medlemsstaternas lagstiftning skall föreskriva att ett kapital på minst 25 000 europeiska beräkningsenheter måste tecknas för att bolaget skall få bildas eller få tillstånd att börja sin verksamhet.
Med en europeisk beräkningsenhet avses en sådan enhet som har bestämts genom kommissionens beslut nr 3289/75/EKSG (4). Som motvärde i nationell valuta gäller första gången motvärdet den dag då detta direktiv antas.
3. Med hänsyn till den ekonomiska och monetära utvecklingen inom gemenskapen och till tendensen att tillåta endast större och medelstora företag att välja de i artikel 1.1 angivna bolagsformerna, skall rådet vart femte år på förslag av kommissionen överväga och vid behov ändra de i denna artikel i europeiska beräkningsenheter uttryckta beloppen.
Artikel 7
Det tecknade kapitalet får endast bestå av tillgångar som kan värderas ekonomiskt. I dessa tillgångar får dock inte inräknas åtaganden att utföra arbete eller att tillhandahålla tjänster.
Artikel 8
1. Aktierna får inte ges ut mot vederlag som understiger det nominella beloppet eller, om sådant saknas, det bokförda parivärdet.
2. Medlemsstaterna kan dock tillåta att de som yrkesmässigt åtar sig att placera aktier får betala mindre än fullt belopp för de aktier som de tecknar i ett sådant sammanhang.
Artikel 9
1. Aktier som ges ut mot vederlag måste då bolaget bildas eller får tillstånd att börja sin verksamhet vara betalda till minst 25 procent av det nominella beloppet eller, om sådant saknas, av det bokförda parivärdet.
2. Aktier som har getts ut mot apportegendom innan bolaget bildas eller får tillstånd att börja sin verksamhet skall vara fullt betalda inom fem år från bolagsbildningen eller tillståndet att börja verksamheten.
Artikel 10
1. En eller flera av bolaget oberoende sakkunniga, som utses eller godkänns av en förvaltningsmyndighet eller en domstol, skall avge ett utlåtande om apportegendomen innan bolaget bildas eller får tillstånd att börja sin verksamhet. Beroende på varje medlemsstats lagstiftning kan de sakkunniga vara fysiska eller juridiska personer eller bolag.
2. Sakkunnigutlåtandet skall minst beskriva apportegendomen samt ange vilka värderingsmetoder de sakkunniga har använt och huruvida de därvid beräknade värdena åtminstone motsvarar antal, nominellt värde eller, i avsaknad av sådant värde, bokfört parivärde och i förekommande fall överkurs i fråga om de aktier för vilka apportegendomen utgör vederlag.
3. Sakkunnigutlåtandet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
4. En medlemsstat får underlåta att tillämpa denna artikel om samtliga aktier till 90 procent av sitt nominella värde eller, i avsaknad av sådant värde, av sitt bokförda parivärde utges mot apportegendom från ett eller flera bolag och följande villkor är uppfyllda: a) de i artikel 3 i avsedda personerna eller bolagen med anknytning till det bolag som tar emot apportegendomen har avstått från att kräva sakkunnigutlåtande;
b) avståendet har offentliggjorts enligt punkt 3;
c) de bolag som lämnar apportegendomen har reserver som enligt lag eller bolagsordning inte får delas ut och som uppgår till minst det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet hos de aktier som ges ut mot apportegendom;
d) de bolag som lämnar apportegendomen förklarar, att de med belopp som motsvarar det vid c angivna värdet åtar sig ansvar för skulder som kan uppkomma för det mottagande bolaget från det att detta bolag har gett ut aktierna mot apportegendom till dess att ett år har förflutit från bolagets offentliggörande av årsredovisningen för det räkenskapsår under vilket apportegendomen lämnades; överlåtelse av aktierna får inte ske under denna tid;
e) det vid d angivna ansvaret har offentliggjorts enligt punkt 3;
f) de bolag som lämnar apportegendomen för över ett belopp som motsvarar det vid c angivna värdet till en reserv som får delas ut först tre år efter det att det mottagande bolagets årsredovisning har offentliggjorts för det räkenskapsår under vilket apportegendomen lämnades eller, i förekommande fall, först vid den senare tidpunkt då alla fordringar som omfattas av det vid d angivna ansvaret och som görs gällande under den nu angivna treårsperioden har tillgodosetts.
Artikel 11
1. Om ett bolag inom en tid som av den nationella lagstiftningen skall bestämmas till minst två år från det att bolagets bildades eller tilläts att börja sin verksamhet förvärvar tillgångar från en person eller ett bolag som avses i artikel 3 i mot ett vederlag som motsvarar minst en tiondel av det tecknade kapitalet, skall förvärvet granskas och offentliggöras enligt artikel 10 samt underställas bolagsstämman för godkännande.
Medlemsstaterna får föreskriva att dessa bestämmelser även skall tillämpas när tillgångarna tillhör en aktieägare eller någon annan.
2. Punkt 1 tillämpas inte i fråga om förvärv som sker inom ramen för bolagets löpande verksamhet, på begäran eller under kontroll av en förvaltningsmyndighet eller en domstol eller på en fondbörs.
Artikel 12
Aktieägarna får inte befrias från sin skyldighet att betala aktierna i andra fall än som kan följa av bestämmelserna om nedsättning av det tecknade kapitalet.
Artikel 13
Om ett bolag av annat slag ombildas till aktiebolag skall medlemsstaterna, i avvaktan på en senare samordning av den nationella lagstiftningen, se till att minst de skyddsåtgärder som föreskrivs i artiklarna 2-12 iakttas.
Artikel 14
Artiklarna 2-13 skall inte inverka på medlemsstaternas föreskrifter om kompetens och tillvägagångssätt vid ändring av en bolagsordning eller en stiftelseurkund.
Artikel 15
1. a) Med undantag för det fallet att det tecknade kapitalet sätts ned får någon utdelning inte ske till aktieägarna, om enligt bolagets årsredovisning nettotillgångarna på bokslutsdagen för det senaste räkenskapsåret understiger eller till följd av utdelningen skulle komma att understiga det tecknade kapitalet och de reserver som enligt lag eller bolagsordning inte får delas ut.
b) Det vid a angivna tecknade beloppet skall minskas med sådan icke inbetald del därav som inte redovisas på balansräkningens aktivsida.
c) Det belopp som delas ut till aktieägarna får inte överstiga vinsten för det senast avslutade räkenskapsåret med tillägg för balanserad vinst och belopp från reserver som får användas för detta ändamål samt med avdrag för balanserad förlust och belopp som enligt lag eller bolagsordning har avsatts till reserver.
d) Med "utdelning" avses i a och c särskilt utbetalning av vinst eller ränta som hänför sig till aktierna.
2. Om lagstiftningen i en medlemsstat tillåter förskottsutdelning av vinst skall minst följande villkor iakttas: a) ett delårsbokslut skall upprättas som visar att tillräckliga medel finns tillgängliga för utdelningen;
b) det belopp som skall delas ut får inte överstiga den vinst som har uppkommit efter det senaste räkenskapsår för vilket årsbokslut har upprättats, med tillägg för balanserad vinst och belopp från reserver som får användas för detta ändamål samt med avdrag för balanserad förlust och belopp som enligt lag eller bolagsordning skall föras över till reserver.
3. Punkterna 1 och 2 inkräktar inte på medlemsstaternas bestämmelser om ökning av det tecknade kapitalet genom överföring av reserver till detta.
4. Lagstiftningen i en medlemsstat får föreskriva undantag från punkt 1 a i fråga om förvaltningsbolag med fast kapital.
I denna punkt anses som förvaltningsbolag med fast kapital endast bolag: - som uteslutande har till föremål för sin verksamhet att placera sina medel i olika värdepapper, olika fastigheter eller andra tillgångar i det enda syftet att sprida investeringsriskerna och låta resultatet av kapitalförvaltningen komma aktieägarna till godo, och
- som vänder sig till allmänheten för att placera sina egna aktier.
I den omfattning den nu angivna möjligheten används i medlemsstaternas lagstiftning a) skall denna ålägga bolagen ifråga att föra in ordet "förvaltningsbolag" i alla dokument som anges i artikel 4 i direktiv 68/151/EEG;
b) får denna inte tillåta ett bolag som nu avses och vars nettotillgångar understiger det i punkt 1 a nämnda beloppet att dela ut medel till aktieägarna, om enligt årsredovisningen för det senaste räkenskapsåret summan av bolagets samtliga tillgångar på bokslutsdagen understiger eller till följd av utdelningen skulle komma att understiga en och en halv gånger beloppet av bolagets samtliga skulder enligt årsredovisningen;
c) skall denna föreskriva att ett nu avsett bolag, som delar ut medel till aktieägarna när nettotillgångarna understiger det i punkt 1 a angivna beloppet, skall upplysa om utdelningen i en not till årsredovisningen.
Artikel 16
En utdelning i strid med artikel 15 skall återbetalas av de aktieägare som har mottagit denna, om bolaget visar att aktieägarna kände till att utdelningen var olaglig eller att de med hänsyn till omständigheterna inte kunde vara okunniga om det.
Artikel 17
1. Vid betydande förlust av det tecknade kapitalet skall kallelse inom den tid som anges i medlemsstaternas lagstiftning ske till en bolagstämma, som skall pröva om bolaget skall upplösas eller om andra åtgärder skall vidtas.
2. Gränsen för betydande förlust enligt punkt 1 får i medlemsstaternas lagstiftning inte sättas högre än till hälften av det tecknade kapitalet.
Artikel 18
1. Ett bolag får inte teckna sina egna aktier.
2. Om aktierna i ett bolag har tecknats av någon i eget namn men för bolagets räkning, skall denne anses ha tecknat aktierna för egen räkning.
3. Aktier som har tecknats i strid med denna artikel skall betalas av de i artikel 3 i angivna personerna eller bolagen eller, vid ökning av det tecknade kapitalet, av medlemmarna i styrelsen eller direktionen.
Lagstiftningen i en medlemsstat får dock bestämma att den skall befrias från betalningsansvar som kan visa att han inte har försummat något.
Artikel 19
1. Om lagstiftningen i en medlemsstat tillåter att ett bolag förvärvar egna aktier, antingen direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall enligt den lagstiftningen minst följande villkor gälla för ett sådant förvärv: a) Tillstånd till förvärvet skall lämnas av bolagsstämman som skall ange de närmare förutsättningarna för detta och särskilt det högsta antal aktier som får förvärvas, den tid inom vilken tillståndet gäller, vilken tid inte får överstiga 18 månader, samt vid förvärv mot vederlag det lägsta och högsta vederlaget. Medlemmarna av styrelsen eller direktionen skall se till att de vid b, c och d angivna villkoren iakttas när förvärvet äger rum.
b) Det nominella värdet eller, om sådant värde saknas, det bokförda parivärdet hos de förvärvade aktierna inräknat de aktier som bolaget tidigare har förvärvat och fortfarande innehar samt de aktier som har förvärvats av någon som handlat i eget namn men för bolagets räkning, får inte överstiga tio procent av det tecknade kapitalet.
c) Förvärvet får inte medföra att värdet av nettotillgångarna understiger det belopp som anges i artikel 15.1 a.
d) Förvärvet får endast omfatta helt betalda aktier.
2. Lagstiftningen i en medlemsstat får medge undantag från punkt 1 a första meningen, om ett förvärv av egna aktier är nödvändigt för att bolaget skall undgå en betydande och nära förestående skada. I ett sådant fall skall styrelsen eller direktionen informera den närmast följande bolagsstämman om grunden för förvärvet och syftet med detta, om de förvärvade aktiernas antal och nominella värde eller, i avsaknad av sådant värde, bokförda parivärde, om den andel av det tecknade kapitalet som de förvärvade aktierna utgör samt om vederlaget för aktierna.
3. Medlemsstaterna behöver inte tillämpa punkt 1 a första meningen på aktier som förvärvas av bolaget, direkt eller av någon som handlar i eget namn men för bolagets räkning, för att fördelas bland de anställda i bolaget eller ett detta närstående bolag. Sådana aktier skall fördelas inom 12 månader från förvärvet.
Artikel 20
1. Medlemsstaterna behöver inte tillämpa artikel 19 på: a) aktier som förvärvas för att genomföra ett beslut om nedsättning av kapitalet eller i fall som avses i artikel 39;
b) aktier som förvärvas som ett led i en allmän förmögenhetsövergång;
c) helt betalda aktier som förvärvas utan vederlag eller som utgör inköpsprovision för banker och andra finansinstitut;
d) aktier som förvärvas på grund av en lagstadgad skyldighet eller till följd av ett rättsligt avgörande till skydd för en aktieägarminoritet, särskilt vid fusion, ändring av föremålet för bolagets verksamhet eller av bolagets form, byte av säte till utlandet eller införandet av begränsningar i rätten att överlåta aktier;
e) aktier som förvärvas från en aktieägare på grund av bristande betalning av aktierna;
f) aktier som förvärvas för att hålla minoritetsaktieägare i närstående bolag skadeslösa;
g) helt betalda aktier som förvärvas vid en exekutiv aktion som äger rum för att infria en fordran som bolaget har mot en aktieägare;
h) helt betalda aktier som har getts ut av ett förvaltningsbolag med fast kapital enligt artikel 15.4 andra stycket och som på placerarnas begäran förvärvas av detta bolag eller av ett detta närstående bolag. Artikel 15.4 a skall därvid tillämpas. Ett sådant förvärv får inte medföra att nettotillgångarna understiger det tecknade kapitalet ökat med de reserver som enligt lag inte får delas ut.
2. Aktier som har förvärvats enligt 1 b-g skall dock avyttras inom högst tre år, med mindre det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet av de förvärvade aktierna inräknat de aktier som bolaget har förvärvat genom någon som handlat i eget namn men för bolagets räkning, inte överstiger tio procent av det tecknade kapitalet.
3. Om aktierna inte avyttras inom den tid som anges i punkt 2 skall de förklaras ogiltiga. Lagstiftningen i en medlemsstat kan bestämma att ogiltigförklaringen skall åtföljas av en motsvarande nedsättning av det tecknade kapitalet. En sådan nedsättning skall föreskrivas i den mån förvärvet av de aktier som skall förklaras ogiltiga har medfört att nettotillgångarna kommit att understiga det belopp som anges i artikel 15.1 a.
Artikel 21
Aktier som har förvärvats i strid med artiklarna 19 och 20 skall avyttras inom ett år från förvärvet. Om de inte avyttras inom denna tid tillämpas artikel 20.3.
Artikel 22
1. Om lagstiftningen i en medlemsstat tillåter ett aktiebolag att förvärva egna aktier, direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall lagstiftningen för det fortsatta innehavet av aktierna alltid kräva att minst följande villkor iakttas:
a) av de rättigheter som är knutna till aktier får rösträtt aldrig utövas för de egna aktierna; b) om dessa aktier tas upp som en tillgång i balansräkningen skall ett motsvarande belopp, som bolaget inte får förfoga över, tas upp som en reserv bland skulderna;
2. Om lagstiftningen i en medlemsstat tillåter ett bolag att förvärva egna aktier, direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall lagstiftningen kräva att förvaltningsberättelsen innehåller minst följande uppgifter: a) skälen för de förvärv som har skett under räkenskapsåret;
b) antal och nominellt värde eller, i avsaknad av sådant värde, bokfört parivärde beträffande de aktier som har förvärvats och avyttrats under räkenskapsåret samt den andel av det tecknade kapitalet som dessa aktier utgör;
c) vid förvärv eller avyttring mot vederlag, uppgift om vederlaget för aktierna;
d) antal och nominellt värde eller, i avsaknad av sådant värde, bokfört parivärde beträffande samtliga aktier som har förvärvats och som innehas av bolaget samt den andel av det tecknade kapitalet som dessa aktier utgör.
Artikel 23
1. Ett bolag får inte ge förskott, lämna lån eller ställa säkerhet i syfte att tredje man skall förvärva aktier i bolaget.
2. Punkt 1 tillämpas inte på åtgärder som utgör led i en banks eller något annat finansinstituts löpande verksamhet eller som vidtas i syfte att aktier skall förvärvas av eller till förmån för de anställda i bolaget eller ett detta närstående bolag. Sådana åtgärder får dock inte leda till att nettotillgångarna understiger det belopp som anges i artikel 15.1 a.
3. Punkt 1 tillämpas inte på åtgärder som vidtas för att aktier skall förvärvas enligt artikel 20.1 h.
Artikel 24
1. Om ett bolag direkt eller genom någon som handlar i eget namn men för bolagets räkning tar emot egna aktier som säkerhet, jämställs detta med förvärv som avses i artiklarna 19 och 20.1 samt artiklarna 22 och 23.
2. Medlemsstaterna behöver inte tillämpa punkt 1 på åtgärder i en banks eller något annat finansinstituts löpande verksamhet.
Artikel 25
1. Alla kapitalökningar skall beslutas av bolagsstämman. Ett sådant beslut, liksom genomförandet av kapitalökningen, skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
2. Bolagsordningen, stiftelseurkunden eller bolagsstämman, vilken senares beslut skall offentliggöras enligt punkt 1, får dock ge bemyndigande om att öka det tecknade kapitalet upp till ett högsta belopp som fastställs med hänsyn till eventuella lagregler om sådant högsta belopp. Inom ramen för det fastställda beloppet beslutar det bemyndigade bolagsorganet i förekommande fall om ökning av det tecknade kapitalet. Bemyndigandet gäller i högst fem år och kan förlängas av bolagsstämman en eller flera gånger med högst fem år varje gång.
3. Om det finns flera slag av aktier, skall bolagsstämmans beslut om kapitalökning enligt punkt 1 eller om bemyndigande att öka kapitalet enligt punkt 2 bli föremål för en särskild omröstning minst för varje kategori av aktieägare vilkas rätt berörs av beslutet.
4. Denna artikel tillämpas vid emission av alla värdepapper som kan bytas ut mot aktier eller som är förenade med teckningsrätt till aktier, men inte vid själva utbytet av värdepapperen eller vid utnyttjandet av teckningsrätten.
Artikel 26
Om aktier ges ut mot vederlag som ett led i ökningen av det tecknade kapitalet, skall de betalas med minst 25 procent av aktiernas nominella värde eller, i avsaknad av sådant värde, av det bokförda parivärdet. Om en överkurs fastställs, skall denna betalas helt.
Artikel 27
1. Om aktier ges ut mot apportegendom som ett led i ökningen av det tecknade kapitalet, skall aktierna vara helt betalda inom fem år från beslutet om ökning av det tecknade kapitalet.
3. Medlemsstaterna behöver inte tillämpa punkt 2, om ökningen av det tecknade kapitalet sker för att genomföra en fusion eller ett offentligt erbjudande om köp eller byte och i syfte att ersätta aktieägarna i ett bolag som upplöses genom fusionen eller är föremål för det offentliga erbjudandet om köp eller byte.
4. Medlemsstaterna behöver inte tillämpa punkt 2 när alla aktier som emitteras som ett led i ökningen av det tecknade kapitalet ges ut mot apportegendom från ett eller flera bolag, om alla aktieägare i det bolag som tar emot apportegendomen har avstått från sakkunnigutlåtande samt villkoren i artikel 10.4b-f är uppfyllda.
Artikel 28
Om en kapitalökning inte fulltecknas, skall kapitalet ökas med det tecknade beloppet endast om emissionsvillkoren uttryckligen har föreskrivit det.
Artikel 29
1. Vid varje ökning av det tecknade kapitalet, som skall betalas med pengar, skall aktierna med företrädesrätt erbjudas aktieägarna i förhållande till den andel av kapitalet som deras aktier representerar.
2. Medlemsstaterna a) behöver inte tillämpa punkt 1 på aktier med en begränsad rätt till utdelning enligt artikel 15 och/eller vid utskiftning av bolagets förmögenhet i samband med likvidation; eller
b) får - om i ett bolag med aktier av olika slag i fråga om rösträtt eller rätt till utdelning enligt artikel 15 eller vid utskiftning i samband med likvidation, det tecknade kapitalet ökas genom att nya aktier av endast ett av dessa aktieslag ges ut - tillåta att ägarna till aktier av annat slag får utöva sin företrädesrätt att teckna nya aktier först efter ägarna till aktier av det slag som emissionen avser.
3. Erbjudandet om företrädesrätt och den tid inom vilken denna rätt får utnyttjas skall offentliggöras i den nationella tidning som har utsetts i överensstämmelse med direktiv 68/151/EEG. Lagstiftningen i en medlemsstat behöver dock inte föreskriva ett offentliggörande, om alla bolagets aktier är ställda till viss man. I sådant fall skall samtliga aktieägare underrättas skriftligen. Den tid inom vilken företrädesrätten skall utnyttjas får inte understiga 14 dagar från det att erbjudandet offentliggörs eller den skriftliga underrättelsen avsänds.
4. Företrädesrätten får inte begränsas eller upphävas i bolagsordningen eller stiftelseurkunden. Detta får däremot ske genom ett beslut av bolagsstämman. Direktionen eller styrelsen skall i så fall lämna bolagsstämman en skriftlig redogörelse som anger skälen för att begränsa eller upphäva företrädesrätten och grunderna för den föreslagna emissionskursen. Bolagsstämmans beslut skall fattas enligt bestämmelserna i artikel 40 om beslutförhet och majoritet. Beslutet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
5. Lagstiftningen i en medlemsstat får bestämma att bolagsordningen, stiftelseurkunden eller bolagsstämman, den senare med iakttagande av bestämmelserna i punkt 4 angående beslutförhet, majoritet och offentliggörande, kan bemyndiga det bolagsorgan att begränsa eller upphäva företrädesrätten som har rätt att besluta om ökning av aktiekapitalet inom gränserna för det "auktoriserade" kapitalet. Ett sådant bemyndigande får inte gälla för längre tid än ett bemyndigande enligt artikel 25.2.
6. Punkterna 1-5 tillämpas vid emission av alla värdepapper som kan bytas ut mot aktier eller som är förenade med teckningsrätt till aktier, men inte vid själva utbytet av värdepapperen eller vid utnyttjandet av teckningsrätten.
7. Företrädesrätten anses inte utesluten enligt punkt 4 eller 5, om aktierna på grund av beslutet om ökning av det tecknade kapitalet ges ut till banker eller andra finansinstitut för att dessa skall erbjuda aktierna till bolagets aktieägare enligt punkterna 1 och 3.
Artikel 30
Artikel 31
Om det finns flera slag av aktier, skall bolagsstämmans beslut om nedsättning av det tecknade kapitalet bli föremål för en särskild omröstning minst för varje kategori av aktieägare vilkas rätt berörs av beslutet.
Artikel 32
1. Om det tecknade kapitalet sätts ned har åtminstone de borgenärer, vilkas fordringar har uppkommit före offentliggörandet av beslutet om nedsättningen, rätt att minst få säkerhet för de fordringar som inte är förfallna till betalning vid offentliggörandet. Lagstiftningen i medlemsstaterna bestämmer under vilka förutsättningar denna rätt får utövas. Lagstiftningen får utesluta rätten endast om en borgenär har tillfredsställande säkerhet eller sådan inte behövs med hänsyn till bolagets ställning.
2. Medlemsstaternas lagstiftning skall vidare minst föreskriva att nedsättningen inte gäller eller att någon utbetalning inte får ske till förmån för aktieägarna, förrän borgenärerna har fått gottgörelse eller en domstol har beslutat att deras framställning därom inte behöver efterkommas.
3. Denna artikel tillämpas även när nedsättningen av det tecknade kapitalet sker genom att bolaget helt eller delvis avstår från betalning av aktieägarnas insatser.
Artikel 33
1. Medlemsstaterna behöver inte tillämpa artikel 32 vid en nedsättning av det tecknade kapitalet som sker för att täcka en inträffad förlust eller för att föra över vissa belopp till en reserv, om reserven därefter inte överstiger tio procent av det nedsatta tecknade kapitalet. Utom vid nedsättning av det tecknade kapitalet får denna reserv inte delas ut till aktieägarna; den får endast användas för att täcka en inträffad förlust eller för att öka det tecknade kapitalet genom överföring av reserver, i den mån medlemsstaterna tillåter en sådan åtgärd.
2. I de fall som avses i punkt 1 skall medlemsstaternas lagstiftning minst föreskriva de åtgärder som behövs för att belopp som härrör från nedsättningen av det tecknade kapitalet inte skall kunna användas för utbetalningar till aktieägarna eller för att befria dessa från skyldigheten att betala sina insatser.
Artikel 34
Det tecknade kapitalet får inte sättas ned under det minimikapital som har fastställts i överensstämmelse med artikel 6. Medlemsstaterna får dock tillåta en sådan nedsättning, om de även föreskriver att beslutet om nedsättning får verkställas först sedan det tecknade kapitalet har ökats till minst det fastställda minimikapitalet.
Artikel 35
Om lagstiftningen i en medlemsstat tillåter att det tecknade kapitalet helt eller delvis löses in utan att kapitalet sätts ned, skall lagstiftningen minst kräva att följande villkor är uppfyllda: a) Om bolagsordningen eller stiftelseurkunden ger möjlighet till inlösen skall beslut om inlösen fattas av bolagstämman, som minst skall iaktta de allmänna villkoren för beslutförhet och majoritet. Om bolagsordningen eller stiftelseurkunden inte ger möjlighet till inlösen skall beslut om inlösen fattas av bolagstämman, som i så fall minst skall iaktta villkoren för beslutförhet och majoritet enligt artikel 40. Beslutet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
b) Endast belopp som får delas ut enligt artikel 15.1 får användas för inlösen.
c) De aktieägare som har fått sina aktier inlösta har kvar sina rättigheter i bolaget med undantag för rätten att återfå insatserna och rätten att delta i en första vinstutdelning avseende icke inlösta aktier.
Artikel 36
1. Om lagstiftningen i en medlemsstat tillåter bolagen att sätta ned det tecknade kapitalet genom att tvångsvis dra in aktier, skall lagstiftningen minst kräva att följande villkor är uppfyllda:
a) Tvångsindragningen skall föreskrivas eller tillåtas i bolagsordningen eller stiftelseurkunden innan teckning sker av de aktier som skall dras in. b) I det fallet att tvångsindragningen endast tillåts i bolagsordningen eller stiftelseurkunden skall den beslutas av bolagstämman, om inte samtliga berörda aktieägare har godkänt indragningen.
c) Det bolagsorgan som beslutar om tvångsindragningen skall bestämma villkor och sätt för denna, om inte det har skett redan i bolagsordningen eller stiftelseurkunden.
d) Artikel 32 tillämpas utom i fråga om helt betalda aktier som ställs till bolagets förfogande utan vederlag eller som dras in med utnyttjande av medel som får delas ut enligt artikel 15.1; i dessa fall skall ett belopp som motsvarar det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet för samtliga indragna aktier föras över till en reserv. Utom vid nedsättning av det tecknade kapitalet får denna reserv inte delas ut till aktieägarna; den får endast användas för att täcka en inträffad förlust eller för att öka det tecknade kapitalet genom överföring av reserver, i den mån medlemsstaterna tillåter en sådan åtgärd.
e) Beslutet om tvångsindragning skall offentliggöras enligt varje lands lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
2. Artikel 30 första stycket samt artiklarna 31, 33 och 40 tillämpas inte i de fall som avses i punkt 1.
Artikel 37
1. Om det tecknade kapitalet sätts ned genom indragning av aktier som bolaget har förvärvat direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall bolagsstämman alltid besluta om indragningen.
2. Artikel 32 tillämpas utom i fråga om helt betalda aktier som har förvärvats utan vederlag eller med medel som får delas ut enligt artikel 15.1; i dessa fall skall ett belopp som motsvarar det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet för samtliga indragna aktier föras över till en reserv. Utom vid nedsättning av det tecknade kapitalet får denna reserv inte delas ut till aktieägarna; den får endast användas för att täcka en inträffad förlust eller för att öka det tecknade kapitalet genom överföring av reserver, i den mån medlemsstaterna tillåter en sådan åtgärd.
3. Artiklarna 31, 33 och 40 tillämpas inte i de fall som avses i punkt 1.
Artikel 38
Om det finns flera slag av aktier skall i de fall som avses i artikel 35, artikel 36.1 b och artikel 37.1 bolagsstämmans beslut om inlösen av det tecknade kapitalet eller nedsättning av detta genom indragning av aktier bli föremål för en särskild omröstning minst för varje kategori av aktieägare vilkas rätt berörs av åtgärden.
Artikel 39
Om lagstiftningen i en medlemsstat tillåter bolagen att ge ut aktier som kan återköpas, skall lagstiftningen för återköp av aktierna minst kräva att följande villkor är uppfyllda: a) återköpet skall tillåtas i bolagsordningen eller stiftelseurkunden innan teckning sker av de aktier som kan återköpas;
b) aktierna skall vara helt betalda;
c) villkoren och sättet för återköpet skall vara bestämda i bolagsordningen eller stiftelseurkunden;
d) återköpet får endast ske med medel som kan delas ut enligt artikel 15.1 eller med intäkter från en nyemission som sker i och för återköpet;
e) ett belopp som motsvarar det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet av alla återköpta aktier skall föras över till en reserv som inte får delas ut till aktieägarna i annat fall än då det tecknade kapitalet sätts ned; denna reserv får endast användas för att öka det tecknade kapitalet genom överföring av reserver;
f) punkt e tillämpas inte, om återköpet har skett med intäkter från en nyemission som har ägt rum i och för återköpet;
g) om det har beslutats att en överkurs skall betalas till aktieägarna med anledning av återköpet, får överkursen endast erläggas med medel som får delas ut enligt artikel 15.1 eller med medel ur en reserv, annan än den som avses i e, som inte får delas ut till aktieägarna i annat fall än då det tecknade kapitalet sätts ned; denna reserv får endast användas för att öka det tecknade kapitalet genom överföring av reserver, för att täcka kostnader som avses i artikel 3 j eller emissionskostnader för aktier eller obligationer eller för att betala en överkurs till innehavare av aktier eller obligationer som skall återköpas;
h) återköpet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
Artikel 40
1. Medlemsstaternas lagstiftning skall föreskriva att de beslut som avses i artikel 29.4 och 5 samt artiklarna 30, 31, 35 och 38 skall kräva minst en majoritet som inte får understiga två tredjedelar av de röster som är förenade med de företrädda värdepapperen eller det företrädda tecknade kapitalet.
2. Medlemsstaternas lagstiftning får dock föreskriva att enkel majoritet av rösterna enligt punkt 1 är tillräcklig, om minst hälften av det tecknade kapitalet är företrätt.
Artikel 41
1. Medlemsstaterna får frångå artikel 9.1, artikel 19.1 a första ledet och b samt artiklarna 25, 26 och 29 i den mån det behövs för att bestämmelser skall kunna antas eller tillämpas som har till ändamål att underlätta för anställda och andra i den nationella lagstiftningen angivna personkategorier att få del i företagens kapital.
2. Medlemsstaterna får underlåta att tillämpa artikel 19.1 a första ledet samt artiklarna 30, 31 och 36-39 på bolag som bildas enligt särskild lagstiftning och som vid sidan av "kapitalaktier" ger ut "arbetsaktier" till förmån för de anställda som ett kollektiv, vilket på bolagsstämman företräds av fullmäktige med rösträtt.
Artikel 42
För att detta direktiv skall kunna genomföras måste medlemsstaternas lagstiftning behandla de aktieägare lika som befinner sig i samma ställning.
Artikel 43
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som behövs för att följa detta direktiv inom två år efter dagen för anmälan. De skall genast underrätta kommissionen om detta.
RÅDETS DIREKTIV av den 25 juli 1977 om renrasiga avelsdjur av nötkreatur (77/504/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 43 och 100 i detta,
med beaktande av Europaparlamentets yttrande(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
med beaktande av följande: Produktionen av nötkreatur upptar en mycket viktig plats i gemenskapens jordbruk. Tillfredsställande resultat är till stor del beroende av användningen av renrasiga avelsdjur.
De flesta medlemsstater har hittills strävat efter att som ett led i den nationella avelspolitiken främja produktionen av husdjur av ett begränsat antal raser som uppfyller särskilda avelsmässiga normer. Raser och normer skiljer sig åt från en medlemsstat till en annan och dessa skillnader hindrar handeln inom gemenskapen.
Om dessa skillnader skall kunna avlägsnas, vilket skulle leda till en ökning av jordbrukets produktivitet på området, måste handeln med alla renrasiga avelsdjur inom gemenskapen gradvis göras fri. En fullständig frihet i handeln förutsätter en ytterligare harmonisering, särskilt i fråga om godkännande för avel.
Medlemsstaterna måste få möjlighet att kräva att härstamningsintyg som är utformade enligt ett gemenskapsförfarande skall uppvisas.
Inom vissa tekniska områden bör åtgärder för genomförande vidtas. För att besluta om sådana åtgärder bör ett förfarande fastställas som leder till ett nära samarbete mellan medlemsstaterna och kommissionen inom Ständiga kommittén för husdjursavel. Till dess att beslut fattas om dessa åtgärder för genomförande skall nu gällande bestämmelser på de områden det är fråga om förbli oförändrade.
Det måste säkerställas att import av renrasiga avelsdjur av nötkreatur från icke-medlemsländer inte får ske på villkor som är mindre stränga än de som tillämpas inom gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I detta direktiv används följande beteckningar med de betydelser som här anges: a) renrasigt avelsdjur av nötkreatur: varje nötkreatur vars föräldrar samt far- och morföräldrar är införda eller registrerade i en stambok för samma ras och som självt är infört i eller är registrerat och berättigat till införande i en sådan stambok. b) stambok: varje bok, förteckning eller dataregister
- som förs av en avelsorganisation eller avelsförening som är officiellt godkänd av den medlemsstat där organisationen eller föreningen bildats, och
- där renrasiga avelsdjur av en viss ras av nötkreatur är införda eller registrerade med uppgifter om deras härstamning.
Artikel 2
Medlemsstaterna skall se till att följande inte får förbjudas, begränsas eller hindras på avelsmässiga grunder: - Handel med renrasiga avelsdjur av nötkreatur inom gemenskapen.
- Handel med sperma och embryon från renrasiga avelsdjur av nötkreatur inom gemenskapen.
- Upprättande av stamböcker förutsatt att de uppfyller kraven enligt artikel 6.
- Godkännande av organisationer eller föreningar som för stamböcker enligt artikel 6.
- Handel inom gemenskapen med tjurar som används för artificiell insemination, om inte annat följer av artikel 3.
Artikel 3
Rådet skall på förslag från kommissionen före den 1 juli 1980 anta gemenskapsbestämmelser för godkännande av renrasiga avelsdjur av nötkreatur för avelsändamål.
Till dess att sådana bestämmelser träder i kraft skall godkännande av renrasiga djur av nötkreatur för avelsändamål, godkännande av tjurar för artificiell insemination samt användning av sperma och embryon lyda under nationell rätt, förutsatt att denna inte är mer restriktiv än den lagstiftning som är tillämplig på renrasiga avelsdjur av nötkreatur, sperma och embryon i den medlemsstat som är destinationsland.
Artikel 4
Avelsorganisationer eller avelsföreningar som är officiellt godkända av en medlemsstat får inte motsätta sig att renrasiga avelsdjur av nötkreatur från andra medlemsstater införs i deras stamböcker, förutsatt att djuren uppfyller de krav som fastställs enligt artikel 6.
Artikel 5
Medlemsstaterna får kräva att renrasiga avelsdjur av nötkreatur samt sperma och embryon från sådana djur vid handel inom gemenskapen skall åtföljas av ett härstamningsintyg som har utformats enligt det förfarande som fastställs i artikel 8, särskilt då det gäller resultat från husdjurskontroll och avelsprövningar.
Artikel 6
1. Följande skall bestämmas enligt det förfarande som fastställs i artikel 8:
- Metoder för husdjurskontroll och avelsprövningar samt metoder för beräkning av djurens avelsvärde.
- Villkor för upprättande av stamböcker.
- Villkor för införande i stamböcker.
- Vilka uppgifter som skall anges i härstamningsintyget.
2. Till dess att bestämmelserna i punkt 1 första, andra och tredje strecksatserna träder i kraft a) skall de officiella kontroller som avses i punkt 1 första strecksatsen och som utförs i varje medlemsstat, samt de stamböcker som för närvarande finns, erkännas av övriga medlemsstater,
b) skall godkännandet av avelsorganisationer eller avelsföreningar även fortsättningsvis regleras av de föreskrifter som för närvarande gäller i varje medlemsstat,
c) skall upprättandet av nya stamböcker även fortsättningsvis uppfylla de villkor som för närvarande gäller i varje medlemsstat.
Artikel 7
Till dess att gemenskapsregler införs på området får de villkor som gäller import av renrasiga avelsdjur av nötkreatur från icke-medlemsländer inte vara mer gynnsamma än de som gäller för handeln inom gemenskapen.
Medlemsstaterna får inte tillåta import av renrasiga avelsdjur av nötkreatur från icke-medlemsländer om inte djuren åtföljs av ett härstamningsbevis som intygar att de är införda eller registrerade i en stambok i det exporterande icke-medlemslandet. Bevis måste framläggas på att djuren är införda i eller registrerade och berättigade till införande i en stambok i gemenskapen.
Artikel 8
1. När det förfarande som fastställs i denna artikel skall tillämpas skall ordföranden utan dröjsmål hänskjuta ärendet till Ständiga kommittén för husdjursavel (i det följande kallad "kommittén"), upprättad genom rådets beslut 77/505/EEG, antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
2. Inom kommittén skall medlemsstaternas röster vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
3. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med en majoritet av 41 röster.
4. Kommissionen skall själv anta förslaget och genomföra det omedelbart om det har tillstyrkts av kommittén. Om förslaget inte har tillstyrkts av kommittén eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas och tillämpa dem omedelbart såvida inte rådet med enkel majoritet har avvisat förslaget.
Artikel 9
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 1979 och skall genast underrätta kommissionen om detta.
Artikel 10
Detta direktiv riktar sig till medlemsstaterna.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(1), senast ändrad genom förordning (EEG) nr 1707/73(2),
med beaktande av rådets förordning nr 162/66/EEG av den 27 oktober 1966 om handeln med oljor och fetter mellan gemenskapen och Grekland(3),
med beaktande av rådets förordning nr 171/67/EEG av den 27 juni 1967 om exportbidrag och avgifter på olivolja(4), senast ändrad genom förordning (EEG) nr 2429/72(5), särskilt artikel 11 i denna, och
med beaktande av följande: I artikel 2 i kommissionens förordning (EEG) nr 616/72 av den 27 mars 1972 om tillämpningsföreskrifter för exportbidrag och avgifter på olivolja(6), senast ändrad genom förordning (EEG) nr 503/76(7), föreskrivs att den rätt att importera med befrielse från avgift som anges i artikel 9 i förordning nr 171/67/EEG, skall beviljas för de kvaliteter av olivolja för vilka det finns ett kontantbidrag.
Kontantbidraget beviljas endast för vissa kvaliteter av olivolja och vissa presentationsformer av oljan. För att förhindra vissa uppgörelser som inte svarar mot sedvanliga exportmönster, bör det föreskrivas att rätten att importera med befrielse från avgift bör medges endast när exporten omfattar varor och presentationsformer för vilka ett kontantbidrag verkligen kan beviljas.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för oljor och fetter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 2 i förordning (EEG) nr 616/72 skall ändras på följande sätt:
"Den rätt till avgiftsfri import som anges i artikel 9.1 i förordning nr 171/67/EEG, skall vara beroende av att exporten omfattar kvaliteter på olivoljan och i förekommande fall presentationsformer, för vilka ett kontantbidrag gäller den dag då ansökan om detta tillstånd lämnas in."
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRSTA DIREKTIV av den 18 april 1978 om ändring av bilagorna till direktiv 66/402/EEG om saluföring av utsäde av stråsäd (78/387/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 66/402/EEG av den 14 juni 1966 om saluföring av utsäde av stråsäd(1), senast ändrat genom rådets direktiv 78/55/EEG(2), särskilt artikel 21a i detta, och
med beaktande av följande: Mot bakgrund av den tekniska och vetenskapliga kunskapsutvecklingen bör bilagorna 1, 2 och 3 till ovannämnda direktiv ändras av de skäl som anges nedan.
Villkoren för certifiering av majsutsäde bör anpassas till befintliga internationella program för sortcertifiering av utsäde.
I syfte att förbättra kvaliteten på utsäde bör bestämmelser antas om villkoren för föregående skörd.
I syfte att höja det genetiska värdet på utsäde bör bestämmelser om standarder för sortrenhet som måste uppfyllas av grödan antas för ytterligare ett antal arter.
Vissa standarder som skall uppfyllas av utsäde av ris bör anpassas till den utsädeskvalitet som normalt uppnås.
För att uppfylla villkoren för officiella undersökningar av utsäde som utförs i enlighet med gällande internationella metoder är det nödvändigt att ändra vissa bestämmelser.
I den situation som för närvarande råder har det inte varit möjligt att uppnå fullständig harmonisering inom gemenskapen av de villkor som gäller för förekomst a
KOMMISSIONENS DIREKTIV av den 19 maj 1978 om anpassning till teknisk utveckling av rådets direktiv 76/114/EEG om tillnärmning av medlemsstaternas lagstiftning om föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt på motorfordon och släpvagnar till dessa fordon (78/507/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(1), i dess lydelse enligt anslutningsakten och särskilt artiklarna 11, 12 och 13 i denna,
med beaktande av rådets direktiv 76/114/EEG av den 18 december 1975 om tillnärmning av medlemsstaternas lagstiftning om föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt på motorfordon och släpvagnar till dessa fordon(2), och
med beaktande av följande: Den internationella standardiseringsorganisationen ISO har nu antagit två internationella standarder om ett världstäckande klassificeringssystem, som gör det möjligt att identifiera tillverkaren av ett fordon(3) och även fordonet(4). Det är därför lämpligt att införa i direktiv 76/114/EEG detta system för identifiering av tillverkare, och samtidigt anpassa kraven om identifiering av fordon i direktivet med ISO-standarden.
Bestämmelserna i detta direktiv har tillstyrkts av Kommittén för anpassning till teknisk utveckling av direktiv om avskaffande av tekniska handelshinder inom motorfordonssektorn.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till direktiv 76/114/EEG ändras enligt bilagan till detta direktiv.
Artikel 2
1. Från den 1 oktober 1978 får ingen medlemsstat, av skäl som hänför sig till föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt, - vägra att bevilja EEG-typgodkännande för en fordonstyp, vägra att utfärda det dokument som anges i artikel 10.1 sista strecksatsen i direktiv 70/156/EEG, eller vägra att bevilja nationellt typgodkännande, eller
- förbjuda att fordon tas i bruk
om föreskrivna skyltar och märkningar samt deras placering och fastsättning på fordonstypen eller fordonet överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
2. Från den 1 oktober 1981 gäller följande: - Medlemsstaterna får inte längre utfärda den handling som anges i artikel 10.1 sista strecksatsen i direktiv 70/156/EEG för en typ av fordon för vilka föreskrivna skyltar och märkningar samt deras placering och fastsättning inte överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
- Medlemsstaterna får vägra att bevilja nationellt typgodkännande för en typ av fordon för vilken föreskrivna skyltar och märkningar samt deras placering och fastsättning inte överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
3. Från den 1 oktober 1981 får medlemsstaterna förbjuda att fordon tas i bruk om deras föreskrivna skyltar och märkningar samt placering och fastsättning inte överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
Artikel 3
Medlemsstaterna skall senast den 1 oktober 1978 sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv och skall genast underrätta kommissionen om detta.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EEG) nr 1883/78 av den 2 augusti 1978 om allmänna bestämmelser för finansiering av interventioner genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 729/70 av den 21 april 1970 om finansiering av den gemensamma jordbrukspolitiken(1), senast ändrad genom förordning (EEG) nr 2788/72(2), särskilt artikel 3.2 i denna,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(3), och
med beaktande av följande: I enlighet med artikel 3.2 i förordning (EEG) nr 729/70 bör allmänna bestämmelser för gemenskapsfinansiering av interventioner fastställas.
För detta ändamål bör en förteckning utarbetas över de åtgärder som motsvarar begreppet intervention för stabilisering av marknaderna.
Det bör fastställas att utgifter i samband med interventionsåtgärder för vilka ett belopp per enhet bestäms inom ramen för en gemensam organisation av marknaderna helt skall täckas av gemenskapsmedel.
För de interventionsåtgärder för vilka ett belopp per enhet inte bestäms inom ramen för den gemensamma organisationen av marknaderna, bör grundläggande regler fastställas särskilt vad avser metoden för bestämning av de belopp som skall finansieras, finansieringen av utgifter som följer av att nödvändiga medel binds upp för interventionsköp av produkter, värderingen av lager som skall överföras från ett räkenskapsår till nästföljande och finansieringen av utgifter i samband med lagring och vid behov i samband med bearbetning.
De olika utgifts- och intäktsslagen för varje sektor på grundval av dessa regler bör bli föremål för närmare bestämmelser. Under tiden bör finansieringsförordningarna för varje sektor fortsätta att gälla.
De allmänna bestämmelserna för gemenskapsfinansiering av interventioner bör samlas i en enda förordning. Rådets förordning (EEG) nr 2824/72 av den 28 december 1972 om allmänna bestämmelser för finansiering av interventioner genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket(4) bör därför upphävas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De åtgärder som förtecknas i bilagan motsvarar begreppet intervention för stabilisering av jordbruksmarknaderna enligt artikel 3.1 i förordning (EEG) nr 729/70.
Artikel 2
När, inom ramen för den gemensamma organisationen av marknaden, ett belopp fastställs per enhet för en interventionsåtgärd skall utgifterna i samband med detta helt täckas av gemenskapsmedel.
Artikel 3
När det inom ramen för den gemensamma organisationen av marknaden inte fastställs ett belopp per enhet för en interventionsåtgärd, skall denna finansieras av garantisektionen vid EUGFJ i enlighet med de bestämmelser som anges i artikel 4 8.
Artikel 4
2. För övriga interventionsåtgärder som anges i artikel 3 skall finansieringen vara lika med utgifterna med avdrag för eventuella intäkter som interventionsåtgärden medför.
Artikel 5
I fråga om medel som har sitt ursprung i medlemsstaterna och som används till interventionsköp av produkter, skall de räntekostnader som skall finansieras av garantisektionen vid EUGFJ beräknas enligt en metod och en räntesats som är enhetlig inom hela gemenskapen och som skall fastställas enligt det förfarande som avses i enlighet med artikel 13 i förordning (EEG) nr 729/70. Räntesatsen skall vara representativ för de faktiska räntesatser som tillämpas.
Artikel 6
Materiella åtgärder i samband med lagring och, i förekommande fall, bearbetning av interventionsprodukter, skall finansieras av garantisektionen vid EUGFJ med hjälp av schablonbelopp som är enhetliga inom hela gemenskapen och som skall fastställas enligt förfarandet i artikel 13 i förordning (EEG) nr 729/70, vid behov efter granskning av ärendet i den berörda förvaltningskommittén.
Artikel 7
Om de aktuella produkterna till följd av lagringen minskar i värde, skall den finansiella effekten av denna värdeminskning fastställas och bokföras när produkten övergår i intervention. För detta ändamål skall värdeminskningskoefficienterna och de priser för vilka de skall tillämpas bestämmas enligt förfarandet i artikel 26 i rådets förordning (EEG) nr 2727/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för spannmål(14), senast ändrad genom förordning (EEG) nr 1254/78(15), eller motsvarande artikel i övriga förordningar om den gemensamma organisationen av jordbruksmarknaderna, och vid behov efter granskning i EUGFJ-kommittén.
Artikel 8
I de årsräkenskaper som anges i artikel 4.1 skall de kvantiteter lagrade produkter som skall överföras till påföljande räkenskapsår som regel värderas till sina inköpspriser. För detta ändamål skall det pris som skall tillämpas för kvantiteter som överförs till påföljande räkenskapsår fastställas för de olika produkterna enligt förfarandet i artikel 13 i förordning (EEG) nr 729/70, på grundval av de inköpspriser som betalats av interventionsorganen under en referensperiod och med beaktande av den värdeminskning som anges i artikel 7.
Om det beräknade priset för en given produkt när interventionen upphör är väsentligt lägre än värdet av de lager som skall överföras, värderade enligt det förfarande som anges i första stycket, får dock beslut fattas om att ersätta det inköpspris som interventionsorganen betalat med ett annat pris. Detta pris skall fastställas enligt förfarandet i artikel 13 i förordning (EEG) nr 729/70, vid behov efter granskning i den berörda förvaltningskommittén. Det får inte vara lägre än de genomsnittliga inköpspriserna och de priser som erhålls vid avyttring av interventionslager.
Artikel 9
Vid behov skall tillämpningsföreskrifter för denna förordning antas i enlighet med förfarandet i artikel 13 i förordning (EEG) nr 729/70.
Artikel 10
Förordning (EEG) nr 2824/72 upphör att gälla.
Artikel 11
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(1), senast ändrad genom direktiv 78/547/EEG(2), och särskilt artiklarna 11, 12 och 13 i detta,
med beaktande av rådets direktiv 71/320/EEG av den 26 juli 1971 om tillnärmning av medlemsstaternas lagstiftning om bromsutrustning på vissa kategorier av motorfordon och släpvagnar till dessa fordon(3), i dess lydelse enligt kommissionens direktiv 75/524/EEG(4), och med beaktande av följande:
Med hänsyn till vunna erfarenheter och den tekniska utvecklingen är det nu möjligt att göra kraven strängare och att anpassa dem bättre till faktiska provningsförhållanden.
Bestämmelserna i detta direktiv är i överenstämmelse med yttrandet från Kommittén för anpassning till teknisk utveckling av direktiv om avskaffande av tekniska handelshinder inom motorfordonssektorn.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Bilagorna 1, 2, 3, 4, 5, 6 och 9 till direktiv 71/320/EEG ändras härmed enligt bilagan till detta direktiv.
2. I väntan på att särskilda bestämmelser angående låsningsfria bromssystem skall träda i kraft, skall fordon i kategorierna M1, M2, M3, N1, N2, N3, O3 och O4 som är utrustade med sådana system underkastas bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
Artikel 2
1. Från den 1 januari 1980 får ingen medlemsstat, av skäl som hänför sig till bromsutrustningen,
- vägra att bevilja EEG-typgodkännande eller att utfärda det exemplar av det intyg som anges i sista strecksatsen i artikel 10.1 i direktiv 70/156/EEG eller att bevilja ett nationellt typgodkännande med avseende på en fordonstyp, eller
- förbjuda att fordon tas i bruk,
om bromsutrustningen på fordonstypen eller fordonen överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
2. Från den 1 oktober 1980 skall medlemsstaterna
- inte längre utfärda det exemplar av det intyg som anges i sista strecksatsen i artikel 10.1 i direktiv 70/156/EEG med avseende på en fordonstyp vars bromsutrustning inte överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv,
- vägra att bevilja ett nationellt typgodkännande för en fordonstyp vars bromsutrustning inte överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
3. Från den 1 oktober 1981 får medlemsstaterna förbjuda ibruktagande av fordon vars bromsutrustning inte överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
4. Utan hinder av punkterna 1-3 skall medlemsstaterna tillämpa bestämmelserna i punkt 1.2.1 i bilaga 4 till direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv, endast från den 1 oktober 1983.
5. Före den 1 januari 1980 skall medlemsstaterna sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv och genast underrätta kommissionen om detta.
Artikel 3
KOMMISSIONENS FÖRORDNING (EEG) nr 883/79 av den 3 maj 1979 om ändring av förordning (EEG) nr 2960/77 om närmare bestämmelser för försäljning av olivolja som innehas av interventionsorgan
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(1), senast ändrad genom förordning (EEG) nr 590/79(2), särskilt artikel 12.4 i denna, och
med beaktande av följande: I artikel 6 i kommissionens förordning (EEG) nr 2960/77(3) föreskrivs att eventuella köpare får ta ett prov på de oljor som säljs av interventionsorganen.
För att säkerställa att den olja som anbudet gäller och den olja som tilldelats är identiska, bör det vara möjligt att ta ytterligare ett prov innan det tilldelade partiet plomberas.
För att underlätta avhämtningen av de sålda oljorna bör avhämtningstidens längd ändras genom att den anpassas efter det tilldelade partiets storlek.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för oljor och fetter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 2960/77 skall ändras på följande sätt: 1. Artikel 5.3 skall ersättas med följande:
"3. Under perioden från och med den 1 januari till och med 31 december 1979 skall minimipriset vara exklusive skatt och hänföra sig till 100 kg olivolja som levereras fritt lager, antingen i köparens egna fat och lastad på ett fordon som tillhandahållits av honom, eller i köparens tankfordon."
2. Artikel 6 andra stycket skall ersättas med följande:
"Detta prov skall placeras i två etiketterade flaskor, som skall plomberas i närvaro av både den som är ansvarig för lagret och den eventuelle köparen eller dennes vederbörligen bemyndigade företrädare. En flaska skall lämnas till den eventuelle köparen och den andra till den som är ansvarig för lagret."
"Artikel 10Interventionsorganet skall genast meddela varje anbudsgivare med rekommenderat brev med mottagningsbevis om resultatet av hans deltagande i anbudsförfarandet."
4. Följande stycke skall läggas till i artikel 11.1:
"Innan plomberingen utförs får den vars anbud antagits begära ett prov på denna olja. Detta prov skall placeras i två etiketterade flaskor, som skall plomberas i närvaro av både den som är ansvarig för lagret och den vars anbud antagits eller dennes vederbörligen bemyndigade företrädare. En flaska skall lämnas till anbudsgivaren och den andra till den som är ansvarig för lagret så att det vid behov kan kontrolleras att den vara som ett prov togs på enligt artikel 6 och den vara som tilldelats stämmer överens."
1. Köparen skall, innan han avhämtar oljan, betala det preliminära försäljningspriset till interventionsorganet. Detta skall beräknas genom att multiplicera den kvantitet som enligt uppgift fanns i partiet med det pris som erbjudits för partiet.
2. Om det preliminära beloppet inte betalas inom den tid som anges i artikel 13.1, skall köpet automatiskt upphävas. I sådana fall skall den säkerhet som avses i artikel 8 förverkas.
2. Den kvantitet olja som levererats till köparen får avvika från den kvantitet för vilken anbudet lämnades, beroende på den faktiska kvantiteten i behållaren vid leveranstillfället."
8. Artikel 21 andra stycket skall utgå.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS ELFTE DIREKTIV av den 26 mars 1980 om harmonisering av medlemsstaternas lagstiftning om omsättningsskatt - uteslutning av de franska utomeuropeiska departementen från tillämpningsområdet för direktiv 77/388/EEG (80/368/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 99 och 100 i detta,
med beaktande av kommissionens förslag, och
med beaktande av följande: Enligt artikel 227.2 tredje stycket i fördraget skall gemenskapens institutioner inom ramen för den ordning som anges i fördraget sörja för att den ekonomiska och sociala utvecklingen i de franska utomeuropeiska departementen möjliggörs.
I överensstämmelse med domstolens dom av den 10 oktober 1978 i mål 148-77 tillämpas fördraget och härledd lagstifting på de franska utomeuropeiska departementen, såvida inte gemenskapens institutioner beslutar om särskilda åtgärder som är anpassade till de ekonomiska och sociala villkoren i dessa departement.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande strecksats skall läggas till i artikel 3.2 i direktiv 77/388/EEG"- Frankrike:
de utomeuropeiska departementen."
Artikel 2
Detta direktiv skall tillämpas från och med den 1 januari 1979.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EEG) nr 1698/80 av den 30 juni 1980 om tillägg till förordning (EEG) nr 797/80 om justering av förutfastställda exportavgifter och exportbidrag för socker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3330/74 av den 19 december 1974 om den gemensamma organisationen av marknaden för socker(), senast ändrad genom förordning (EEG) nr 1396/78(), särskilt artiklarna 17.5, 19.2 och 19.4 i denna, och
med beaktande av följande: Enligt kommissionens förordning (EEG) nr 797/80 av den 31 mars 1980 om justering av förutfastställda exportavgifter och exportbidrag för socker() skall exportbidragen höjas och exportavgifterna sänkas i fråga om exportlicenser som utfärdats före den 1 juli 1980 men som utnyttjas först efter detta datum.
När det gäller exportavgifterna kan det förekomma att avgiftsbeloppet är lägre än det belopp med vilket justeringen skall göras. För att undvika att företagen blir olika behandlade måste därför ett tillägg göras till den aktuella förordningen, enligt vilket skillnaden skall betraktas som ett exportbidrag som ges till den berörda parten i stället för utkrävandet av exportavgiften.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för socker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 1 i förordning (EEG) nr 797/80 skall ändras på följande sätt: 1. I punkt 1 skall "på begäran av berörd part" utgå.
2. I punkt 2 skall följande läggas till som ett tredje stycke:
"Om exportavgiften är lägre än det belopp med vilket den skall justeras, skall skillnaden mellan de två beloppen betraktas som ett exportbidrag som skall ges till den berörda parten. I sådana fall skall exportavgiften inte betalas."
Artikel 2
Denna förordning träder i kraft den 1 juli 1980.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS DIREKTIV av den 20 juli 1981 om ändring av rådets direktiv 77/541/EEG om tillnärmning av medlemsstaternas lagstiftning om bilbälten och fasthållningsanordningar i motorfordon (81/576/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Rådets direktiv 77/541/EEG av den 28 juni 1977 om tillnärmning av medlemsstaternas lagstiftning om bilbälten och fasthållningsanordningar i motorfordon(4) uppställer bl.a. i bilaga 1 krav på montering av bilbälten och fasthållningsanordningar i fordon i kategori M1 enligt definition i bilaga 1 i rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(5), senast ändrat genom direktiv 80/1267/EEG(6).
Av trafiksäkerhetsskäl bör hädanefter montering av bilbälten och fasthållningsanordningar som överensstämmer med direktiv 77/541/EEG krävas i fordon i vissa M- och N-kategorier, och monteringen av dessa tillåtas och främjas i fordon i de övriga M- och N-kategorierna genom en utvidgning av räckvidden för detta direktiv. En sådan utvidgning har möjliggjorts av den tekniska utvecklingen i fråga om konstruktion av motorfordon.
Av detta skäl bör direktiv 77/541/EEG ändras.
Ändring av detta direktiv innebär anpassning till den tekniska utvecklingen av vissa krav i bilagorna till direktiv 77/541/EEG. Ikraftträdandet av bestämmelserna i det nuvarande direktivet bör fås att sammanfalla med ikraftträdandet av bestämmelserna som efter antagande av det nuvarande direktivet kommer att antas för anpassning av kraven i bilagorna till direktiv 77/541/EEG till den tekniska utvecklingen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"Artikel 9
I detta direktiv avses med "fordon" varje motorfordon i kategorierna M och N enligt definition i bilaga 1 till direktiv 70/156/EEG som är avsett att användas på väg, som har minst fyra hjul och som är konstruerat för en högsta hastighet som överstiger 25 km/tim."
2. I bilaga 1: a) Avsnitt 3.1 skall ersättas med följande:
"3.1 Fordonsutrustning
Varje fordon som omfattas av artikel 9 och tillhör kategorierna M1 eller N1 eller kategori M2 (utom fordon med en tillåten största vikt som överstiger 3 500 kg och fordon med utrymmen särskilt utformade för stående passagerare) skall vara utrustade med bilbälten eller fasthållningsanordningar som uppfyller kraven i detta direktiv och har följande bältesarrangemang (som varken medger att låsningsfria upprullningsdon [1.8.1] eller upprullningsdon med manuell upplåsning [1.8.2] kan användas).
I de fall där andra fordon som omfattas av artikel 9 är utrustade med bilbälten eller fasthållningsanordningar skall dessa uppfylla alla krav i detta direktiv med undantag av avsnitten 3.1.1-3.1.3."
b) Avsnitt 3.1.1 skall ersättas med följande:
"3.1.1 För främre yttre sittplatser, trepunktsbilbälte med nödlåsande upprullningsdon med flerfunktion (1.8.4). Följande skall dock gälla: 3.1.1.1 För passagerarsätet är automatiskt låsande upprullningsdon (1.8.3) tillåtna.
3.1.1.2 För passagerarsätet i fordon i kategori M2 anses höftbälten, med eller utan upprullningsdon, som tillräckliga om vindrutan befinner sig utanför den referenszon som definieras i bilaga 2 till direktiv 74/60/EEG.
Med avseende på bilbältena skall vindrutan anses vara en del av referenszonen när den kan komma i statisk kontakt med provningsutrustningen enligt den metod som beskrivs i bilaga 2 till direktiv 74/60/EEG."
c) Avsnitt 3.1.3 skall ersättas med följande:
"3.1.3 På bakre sittplatser i fordon i kategori M1, höftbälten eller trepunktsbälten antingen de är försedda med upprullningsdon eller inte."
d) Lägg till ett nytt avsnitt 3.1.5 enligt följande:
"3.1.5 Oavsett föregående bestämmelser får ett nödlåsande upprullningsdon av typ 4 N (1.8.5) tillåtas i stället för ett upprullningsdon av typ 4 (1.8.4) i fordon i kategorierna N1 och M2, där det på ett tillfredsställande sätt har visats för provningsorganet som ansvarar för provningarna att montering av ett upprullningsdon av typ 4 skulle besvära föraren."
Artikel 2
Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv på samma dag som planerats för ikraftträdandet av bestämmelserna som krävs för att följa det direktiv som skall antas efter detta direktiv enligt artikel 10 i direktiv 77/541/EEG så att kraven i bilagorna till det sistnämnda direktivet kan anpassas till den tekniska utvecklingen. De skall genast underrätta kommissionen om detta.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 19 oktober 1981 om ändring med anledning av Greklands anslutning av direktiv 79/869/EEG om mätmetoder samt provtagnings- och analysfrekvenser avseende ytvatten för dricksvattenframställning i medlemsstaterna (81/855/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 och 235 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1), och
med beaktande av följande: Artikel 11.2 i rådets direktiv 79/869/EEG av den 9 oktober 1979 om mätmetoder samt provtagnings- och analysfrekvenser avseende ytvatten för dricksvattenframställning i medlemsstaterna(2) bör ändras av hänsyn till Greklands anslutning till Europeiska gemenskaperna.
I enlighet med artikel 198 första stycket i fördraget har rådet samrått med Ekonomiska och sociala kommittén om kommissionens förslag. Kommittén hade inte möjlighet att avge sitt yttrande inom den tidsgräns som rådet hade fastställt. Enligt artikel 198 andra stycket i fördraget skall avsaknaden av ett yttrande inte hindra rådet från att vidta åtgärder. Eftersom det är önskvärt att de nödvändiga ändringarna antas snabbt finner rådet det angeläget att utnyttja denna möjlighet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 11.2 i direktiv 79/869/EEG skall "41" ersättas med "45".
Artikel 2
Detta direktiv träder i kraft den 1 januari 1981.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EEG) nr 654/81 av den 10 mars 1981 om ändring av rådets förordning (EEG) nr 3179/78 om Europeiska ekonomiska gemenskapens antagande av konventionen om framtida multilateralt samarbete om fisket i Nordvästatlanten
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(), och
med beaktande av följande: Genom rådets förordning (EEG) nr 3179/78() antog gemenskapen konventionen om framtida multilateralt samarbete om fisket i Nordvästatlanten.
Den 7 juni 1979 antog Nordvästatlantiska fiskeriorganisationens allmänna råd, i enlighet med artikel 20 punkt 2 i den konventionen, med ikraftträdande den 1 januari 1980 sådana ändringar i bilaga 3 till konventionen om framtida multilateralt samarbete om fisket i Nordvästatlanten som rör avgränsningen mellan de statistiska delområdena i farvattnen mellan Grönlands västkust och Kanadas kust.
Konventionens lydelse ändrades därför genom förordning (EEG) nr 653/80() men tillämpningen av ändringen var begränsad till och med den 31 december 1980 eftersom den var avsedd som en interimsåtgärd i enlighet med artikel 103 i fördraget.
Det är därför nödvändigt att förordning 3179/78 slutgiltigt ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag (),
med beaktande av Europaparlamentets yttrande (),
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
med beaktande av följande: Genom förordning nr 79/65/EEG (), senast ändrad genom förordning (EEG) nr 2910/73 () inrättade rådet ett informationssystem för jordbruksföretagens redovisningsuppgifter för att belysa inkomstförhållanden och andra ekonomiska förhållanden i jordbruksföretag i Europeiska ekonomiska gemenskapen.
Informationssystemets undersökningsområde måste bestå av alla jordbruksföretag av en viss ekonomisk storlek, oberoende av om jordbrukaren åtar sig annat arbete utanför företaget.
För att få redovisningsresultat som är tillräckligt enhetliga på gemenskapsnivå bör de rapporterande företagen fördelas efter områden och de olika företagskategorierna genom att undersökningsområdet delas in enligt gemenskapens typologi för jordbruksföretag, fastställd genom beslut 78/463/EEG ().
Alla rapporterande företag som undersöks i medlemsstaterna för registrering av inkomster i jordbruket som underlag för jordbrukspolitiken bör tillhöra gemenskapens informationssystem och antalet rapporterande företag bör därför ökas. Detta antal bör kunna variera inom vissa gränser och beroende på utvecklingen inom jordbruket och kraven på uppgifter från den gemensamma jordbrukspolitiken.
Det nationella samordningsorganet måste ha en nyckelroll i handhavandet av informationssystemet. I detta syfte bör det förses med nya uppgifter.
Erfarenheten visar att det inte längre är önskvärt att införa tilläggsvillkor i det avtal som skall slutas mellan medlemsstaten och bokföringsbyråerna.
Informationssystemets områden skall i största möjliga mån vara identiska med dem som används för att redovisa andra regionala uppgifter som är väsentliga för att skapa riktlinjer för den gemensamma jordbrukspolitiken. I detta avseende bör bilagan till förordning nr 79/65/EEG ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Följande fotnot skall läggas till längst ner på sidan:
"b) " () EGT nr L 148, 5.6.1978, s. 1."
2) Artikel 4 skall ersättas med följande:
"Artikel 4
1. Det undersökningsområde som avses i artikel 1.2 a skall omfatta de jordbruksföretag som är av en storlek som i ekonomiskt avseende är lika med eller större än det tröskelvärde, uttryckt i europeiska storleksenheter (ESE) som definieras genom beslut 78/463/EEG.
2. För att bli behörigt som rapporterande företag skall ett jordbruksföretag
a) ha en storlek som i ekonomiskt avseende är lika med eller större än ett tröskelvärde som fastställs enligt punkt 1,
b) drivas av en jordbrukare som vill och kan sköta redovisningen för jordbruket och är beredd att ställa redovisningsuppgifter från sitt företag till kommissionens förfogande,
c) tillsammans med de övriga företagen och på områdesnivå vara representativt för undersökningsområdet.
3. Det högsta antalet rapporterande företag skall vara 45 000.
4. Tillämpningsföreskrifter till denna artikel, särskilt tröskelvärdet för företagens ekonomiska storlek och antalet rapporterande företag per område, skall fastställas enligt förfarandet i artikel 19."
3) Artikel 5 skall ersättas med följande:
"Artikel 5
1. Varje medlemsstat skall före den 1 februari 1982 inrätta en nationell kommitté för informationssystemet, nedan kallad "den nationella kommittén".
2. Den nationella kommittén skall ha ansvaret för valet av rapporterande företag. För detta ändamål skall dess uppgifter framför allt omfatta godkännandet av
a) planen för val av rapporterande företag, särskilt hur de rapporterande företagen skall fördelas per företagskategori och tillämpningsföreskrifterna för val av företag,
b) rapporten om tillämpningen av planen för val av rapporterande företag.
3. Ordföranden i den nationella kommittén skall utses av medlemsstaten bland medlemmarna i denna kommitté.
Den nationella kommitténs beslut skall vara enhälliga. Om enighet inte kan uppnås skall beslut fattas av en myndighet som medlemsstaten utser.
4. Medlemsstater som har flera områden får för varje område under sin jurisdiktion upprätta en regional kommitté för informationssystemet; nedan kallad "den regionala kommittén".
Den regionala kommittén skall särskilt ha som uppgift att arbeta med det samordningsorgan som anges i artikel 6 för att välja ut rapporterande företag.
5. Tillämpningsföreskrifterna till denna artikel skall antas enligt förfarandet i artikel 19."
4) Artikel 6 skall ersättas med följande:
"Artikel 6
1. Varje medlemsstat skall tillsätta ett samordningsorgan, vars uppgifter skall vara
a) att underrätta den nationella kommittén, de regionala kommittéerna och bokföringsbyråerna om de gällande tillämpningsföreskrifterna och att säkerställa att dessa föreskrifter tillämpas korrekt,
b) att utarbeta och till den nationella kommittén överlämna för godkännande och därefter till kommissionen överlämna
P planen för val av rapporterande företag, vilken skall utarbetas med de senaste statistikuppgifterna som underlag, sammanställd enligt gemenskapens typologi för jordbruksföretag,
P rapporten om genomförandet av planen för val av rapporterande företag,
c) att sammanställa
P förteckningen över rapporterande företag,
P förteckningen över bokföringsbyråer som vill och kan upprätta företagsredovisningar, enligt de avtalsvillkor som anges i artiklarna 9 och 14, d) att sammanställa de företagsredovisningar som bokföringsbyråerna översänt och med hjälp av ett gemensamt kontrollprogram kontrollera att de är korrekt ifyllda,
e) att överlämna de ifyllda företagsredovisningarna till kommissionen omedelbart efter kontrollen,
f) att till den nationella kommittén, de regionala kommittéerna och bokföringsbyråerna överlämna alla förfrågningar om information som avses i artikel 16 och att överlämna svaren på dessa till kommissionen.
2. Tillämpningsföreskrifterna till denna artikel skall utarbetas enligt förfarandet i artikel 19."
5) Artikel 9.2 andra stycket skall upphöra att gälla.
6) Artikel 16.1 skall ersättas med följande:
"1. Den nationella kommittén, de regionala kommittéerna, samordningsorganet och bokföringsbyråerna skall vara skyldiga att, inom sina respektive ansvarsområden, ge kommissionen alla uppgifter som den begär av dem om hur de utför sina arbetsuppgifter vid tillämpningen av denna förordning.
Denna begäran om uppgifter till den nationella kommittén, de regionala kommittéerna eller bokföringsbyråerna och svaren på dessa skall meddelas skriftligen genom samordningsorganet."
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 75 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande (), och
med beaktande av följande: Rådet har samrått med Ekonomiska och sociala kommittén om kommissionens förslag med stöd av artikel 198 första stycket i fördraget. Kommittén har inte kunnat inkomma med sitt yttrande inom den av rådet utsatta tiden. Artikel 198 andra stycket i fördraget tillåter rådet att vidta fortsatta åtgärder även utan sådant yttrande. Rådet anser att denna möjlighet måste utnyttjas med tanke på vikten av att erforderliga ändringar snabbt antas.
Förordning (EEG) nr 1108/70 (), i dess lydelse enligt förordning nr 1384/79 () skall ändras på så sätt att Greklands järnvägsnät tas in i bilagan till sistnämnda förordning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande tillägg skall göras till förteckningen i bilaga 2 till förordning (EEG) nr 1108/70 under punkt "A.1.JÄRNVÄG - Huvudnät" efter rubriken "Förbundsrepubliken Tyskland":
"Grekland
P ¼ñãáíéóðüò Óéäçñïäñüìùí ¸ëëÜäïò A.E. (ÏÓÅ)."
Artikel 2
Denna förordning träder i kraft dagen efter dess offentliggörande i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 66/401/EEG av den 14 juni 1966 om saluföring av utsäde av foderväxter(), senast ändrat genom direktiv 81/126/EEG(), särskilt artikel 21 a i detta,
med beaktande av rådets direktiv 69/208/EEG av den 30 juni 1969 om saluföring av utsäde av olje- och spånadsväxter(), senast ändrat genom direktiv 81/126/EEG, särskilt artikel 20 a i detta, och
med beaktande av följande: Mot bakgrund av den vetenskapliga och tekniska kunskapsutvecklingen bör bilaga 1 och 2 till direktiv 66/401/EEG och 69/208/EEG ändras av nedan angivna skäl.
De villkor som skall uppfyllas för gröda och utsäde, även standarder för sortrenhet, bör ändras så att de överensstämmer med de system för certifiering av utsäde avsett för internationell handel som fastställts av Organisationen för europeiskt ekonomiskt samarbete (OECD). De datum för genomförandet som fastställts i artikel 2, andra strecksatsen, i kommissionens direktiv 78/386/EEG av den 18 april 1978 om ändring av bilagorna till direktiv 66/401/EEG om saluföring av utsäde av foderväxter(), senast ändrat genom direktiv 81/126/EEG, samt i artikel 2.1 första strecksatsen i kommissionens direktiv 78/388/EEG av den 18 april 1978 om ändring av bilagorna till direktiv 69/208/EEG om saluföring av utsäde av olje- och spånadsväxter(), senast ändrat genom direktiv 81/126/EEG, bör följaktligen anpassas till den aktuella situationen.
Det har i det nuvarande läget inte varit möjligt att, i fråga om solroshybrider, föreskriva om en harmonisering inom gemenskapen av de minimistandarder för sortrenhet som grödor och utsäde måste motsvara. Ett försök skall dock göras före den 1 juli 1983 att upprätta sådana standarder i syfte att uppnå en harmonisering.
De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga kommittén för utsäde och uppförökningsmaterial för jordbruk, trädgårdsnäring och skogsbruk.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga 1 till direktiv 66/401/EEG ändras på följande sätt:
1. I andra och tredje meningen i punkt 4 skall orden "Vicia faba" tilläggas efter "Pisum sativum".
2. I andra och tredje meningen i punkt 4 skall orden "Raphanus sativus ssp. oleifera" utgå.
Artikel 2
Bilaga 2 till direktiv 66/401/EEG ändras på följande sätt:
1. Punkt 1 i avsnitt I skall ersättas med följande:
Lägsta sortrenhet skall främst undersökas vid fältbesiktningar som utförs enligt de villkor som fastställts i bilaga 1."
Artikel 3
Bilaga 1 till direktiv 69/208/EEG ändras på följande sätt:
Punkt 3 skall ersättas med följande:
- en per 30 m² vid produktion av basutsäde,
- en per 10 m² vid produktion av certifikatutsäde."
Artikel 4
Bilaga 2 till direktiv 69/208/EEG ändras på följande sätt:
Punkt 1 i avsnitt I skall ersättas med följande:
"Utsädet skall ha tillräcklig sortäkthet och sortrenhet. I synnerhet skall utsäde av nedan angivna arter motsvara följande standarder eller andra villkor:
>Plats för tabell>
Lägsta sortrenhet skall främst undersökas vid fältbesiktningar som utförs enligt de villkor som fastställts i bilaga 1."
Artikel 5
I artikel 2.1 andra strecksatsen i direktiv 78/386/EEG skall "den 1 januari 1982" ersättas med "vid ett datum som kommer att fastställas senare".
Artikel 6 I artikel 2.1 första strecksatsen i direktiv 78/388/EEG skall "den 1 januari 1982" ersättas med "vid ett datum som kommer att fastställas senare".
Artikel 7
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa:
- bestämmelserna i artikel 5 och 6, med verkan från och med den 1 januari 1982,
- bestämmelserna i artikel 2 i fråga om Poa spp., med verkan från och med den 1 januari 1983,
- de övriga bestämmelserna i detta direktiv, senast den 1 januari 1983.
2. Medlemsstaterna skall se till att utsäde inte underkastas några begränsningar av saluföringen till följd av olika datum för genomförandet av detta direktiv i enlighet med punkt 1, tredje strecksatsen.
Artikel 8
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av protokollet om immunitet och privilegier för Europeiska gemenskaperna, särskilt artikel 13 i detta,
med beaktande av kommissionens förslag, och
RÅDETS BESLUT av den 26 oktober 1983 om motåtgärder inom den internationella handelssjöfarten (83/573/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 84.2 i detta, och
med beaktande av följande: Utfallet av det informationssystem för sjöfarten som inrättades genom föreskrifterna i besluten 78/774/EEG (), 79/4/EEG (), 80/1181/EEG (), 81/189/EEG () och 82/870/EEG () samt vissa medlemsstaters erfarenhet visar att det skulle vara välbetänkt att inom gemenskapen inrätta ett lämpligt förfarande för motåtgärder inom den internationella handelssjöfarten som berörda medlemsstater kan vidta gentemot tredje länder.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 3
Vid samrådsförfarande enligt artikel 1 bör medlemsstaterna om så är lämpligt i största möjliga utsträckning ange a) den utveckling som har orsakat att motåtgärder vidtagits,
b) det område där motåtgärden skall tillämpas,
c) den typ av sjöfartstjänst som berörs (t.ex. linjefart),
d) den typ av motåtgärder som har vidtagits eller skall vidtas,
e) den tid under vilken motåtgärden skall tillämpas,
f) motåtgärdens rimlighet i förhållande till skadan.
Artikel 4
Det står medlemsstaterna fritt att ensidigt tillämpa nationella motåtgärder.
Artikel 5
Beslutet riktar sig till medlemsstaterna.
RÅDETS ÅTTONDE DIREKTIV av den 10 april 1984 grundat på artikel 54.3 g i fördraget, om godkännande av personer som har ansvar för lagstadgad revision av räkenskaper (84/253/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 54.3 g i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
med beaktande av följande: Enligt direktiv 78/660/EEG (4) skall årsbokslutet i vissa företagsformer revideras av en eller flera personer som är behöriga att företa sådan revision. Endast företag som anges i artikel 11 i det direktivet får undantas från revisionen.
Direktivet har kompletterats med direktiv 83/349/EEG (5) om sammanställd redovisning.
Kvalifikationskraven måste harmoniseras i fråga om de personer som är behöriga att genomföra lagstadgad revision av räkenskaper. Det bör säkerställas att sådana personer är oberoende och har ett gott anseende.
Genom en yrkesexamen måste en hög nivå garanteras när det gäller de teoretiska kunskaper och den förmåga att praktiskt tillämpa kunskaperna som behövs för en lagstadgad revision av räkenskaper.
Medlemsstaterna måste ges rätt att godkänna personer som, utan att uppfylla alla de krav som ställs på teoretisk utbildning, ändå under lång tid genom yrkesmässig verksamhet har fått tillräcklig erfarenhet inom områdena ekonomi, juridik och redovisning samt har godkänts vid yrkesexamen.
Medlemsstaterna måste även ges rätt att besluta om övergångsbestämmelser till förmån för yrkesmässigt verksamma personer.
Medlemsstaterna får godkänna såväl fysiska personer som revisionsbolag, vilka kan vara juridiska personer eller andra former av bolag eller sammanslutningar.
Fysiska personer som utför lagstadgad revision av räkenskaper på ett sådant revisionsbolags vägnar måste uppfylla villkoren i detta direktiv.
En medlemsstat får godkänna personer som utanför den staten har förvärvat kvalifikationer som är likvärdiga med dem som föreskrivs i detta direktiv.
Om en medlemsstat då detta direktiv antas erkänner som revisorer vissa kategorier av fysiska personer vilka uppfyller i direktivet uppställda krav men vilkas yrkesexamen ligger på en lägre nivå än avslutad högskoleutbildning, bör denna medlemsstat i fortsättningen på vissa villkor och till dess ytterligare samordning sker få särskilt godkänna sådana personer att utföra lagstadgad revision i bolag och företagsgrupper av begränsad storlek. En förutsättning bör vara att medlemsstaten inte har utnyttjat de möjligheter till undantag från kravet på lagstadgad revision som lämnas i gemenskapsdirektiven om årsbokslut och sammanställt bokslut.
Detta direktiv berör varken den etableringsfrihet eller den rätt att fritt tillhandahålla tjänster som tillkommer personer med uppgift att utföra lagstadgad revision av räkenskaper.
Frågan om att erkänna ett sådant godkännande att utföra revision som har meddelats en medborgare i en annan medlemsstat kommer att regleras särskilt i direktiv om etablering och utövande av verksamhet inom områdena företagsekonomi, nationalekonomi och redovisning samt i direktiv om frihet att tillhandahålla tjänster inom dessa områden.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
AVSNITT I
Artikel 1
1. De samordningsåtgärder som föreskrivs i detta direktiv skall vidtas i fråga om sådana lagar och andra författningar i medlemsstaterna som avser personer, vilka skall: a) utföra lagstadgad granskning av bolags och andra företags årsbokslut samt verifiera att innehållet i förvaltningsberättelserna är förenligt med årsboksluten, förutsatt att sådan granskning och verifiering föreskrivs i gemenskapsrätten,
b) utföra lagstadgad granskning av sammanställda bokslut och verifiera att innehållet i de sammanställda förvaltningsberättelserna är förenligt med de sammanställda boksluten, förutsatt att sådan granskning och verifiering föreskrivs i gemenskapsrätten.
2. Beroende på varje medlemsstats lagstiftning kan de i punkt 1 angivna personerna vara fysiska personer eller juridiska personer eller andra former av bolag eller sammanslutningar (revisionsbolag enligt definitionen i detta direktiv).
AVSNITT II Regler om godkännande
Artikel 2
1. Lagstadgad revision av de i artikel 1.1 angivna handlingarna får endast utföras av godkända personer. Medlemsstaternas myndigheter får endast godkänna: a) Fysiska personer som uppfyller minst de villkor som anges i artikel 3-19.
b) Revisionsbolag som uppfyller minst följande villkor: i) De fysiska personer som på revisionsbolagets vägnar utför lagstadgad revision av de i artikel 1 angivna handlingarna skall uppfylla minst de i artikel 3-19 angivna villkoren; medlemsstaterna får föreskriva att sådana fysiska personer även skall vara godkända.
ii) En majoritet av röstetalet skall tillkomma fysiska personer eller revisionsbolag som uppfyller minst de i artikel 3-19 uppställda villkoren, med undantag för artikel 11.1 b; medlemsstaterna får föreskriva att sådana fysiska personer och revisionsbolag även skall vara godkända. De medlemsstater som då detta direktiv antas inte kräver nu angiven majoritet behöver dock inte föreskriva sådan, förutsatt att alla aktier eller andra andelar i revisionsbolaget är ställda till viss man och kan överlåtas endast med samtycke av revisionsbolaget och/eller, om medlemsstaten föreskriver det, med godkännande av behörig myndighet.
iii) En majoritet av ledamöterna i revisionsbolagets förvaltnings- eller ledningsorgan måste vara fysiska personer eller revisionsbolag som uppfyller minst de i artikel 3-19 uppställda villkoren; medlemsstaterna får föreskriva att sådana personer eller revisionsbolag även skall vara godkända. Om ett organ inte har fler än två ledamöter, måste en av dessa minst uppfylla de angivna villkoren.
Med förbehåll för vad som gäller enligt artikel 14.2 skall godkännandet av ett revisionsbolag återkallas när något av kraven i b inte längre är uppfyllt. Medlemsstaterna får dock förordna om en frist på högst två år för att uppfylla kraven i b ii och iii.
2. Då bestämmelserna i detta direktiv tillämpas, får de uppgifter som ankommer på medlemsstaternas myndigheter utövas av yrkesföreningar, om dessa enligt nationell lagstiftning har befogenhet att lämna sådant godkännande som avses i direktivet.
Artikel 3
Myndigheterna i en medlemsstat skall godkänna endast personer som har ett gott anseende och inte utövar någon form av verksamhet som enligt medlemsstatens lagar är oförenlig med lagstadgad revision av de i artikel 1.1 angivna handlingarna.
Artikel 4
En fysisk person får godkännas att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna, endast om han efter att ha kvalificerat sig för tillträde till universitetsstudier har genomgått en teoretisk och praktisk utbildning samt avlagt en statligt organiserad eller godkänd yrkesexamen som är jämförbar med slutexamen från ett universitet.
Artikel 5
Det i examen ingående teoretiska kunskapsprovet måste särskilt omfatta följande ämnesområden: a) - räkenskapsrevision,
- balansanalys,
- extern redovisning,
- sammanställd redovisning,
- kostnadsbokföring och internredovisning,
- intern revision och kontroll,
- föreskrifter om upprättande av års- och sammanställt bokslut samt föreskrifter om metoder för värdering av balansposter och beräkning av resultatposter,
- rättsliga och yrkesmässiga normer för lagstadgad revision och för dem som utför sådan revision,
b) i den utsträckning det har betydelse för revisionen: - associationsrätt,
- lagstiftning om konkurs och liknande förfaranden,
- beskattningsrätt,
- civil- och handelsrätt,
- lagstiftning om social trygghet och arbetsrätt,
- informations- och databehandling,
- företagsekonomi, nationalekonomi och finansiering,
- matematik och statistik,
- grundläggande principer för ekonomisk styrning av företag.
Artikel 7
1. Med avvikelse från bestämmelserna i artikel 5 och 6 får en medlemsstat föreskriva att personer med universitetsexamen eller annan likvärdig examen eller med likvärdiga betyg i ett eller flera av de i artikel 6 angivna ämnena, får befrias från att avlägga teoretiska kunskapsprov i de ämnen som täcks av denna examen eller dessa betyg.
2. Med avvikelse från bestämmelserna i artikel 5 får en medlemsstat föreskriva att den som har en akademisk examen eller motsvarande kompetens i ett eller flera av de i artikel 6 angivna ämnena får befrias från att avlägga prov som avser hans förmåga att praktiskt tillämpa kunskaperna i dessa ämnen, om han har fått en praktisk utbildning i ämnena som dokumenteras genom av staten erkända examen eller betyg.
Artikel 8
1. För att garantera förmågan att praktiskt tillämpa de teoretiska kunskaperna, vilken förmåga även prövas i examen, skall under minst tre år en praktisk utbildning äga rum som bl.a. skall omfatta revision av årsbokslut och sammanställda bokslut eller liknande redovisningshandlingar. Denna praktiska utbildning måste till minst två tredjedelar fullgöras hos någon som enligt medlemsstatens lagstiftning är godkänd i överensstämmelse med detta direktiv; medlemsstaten får dock tillåta att den praktiska utbildningen fullgörs hos någon som enligt en annan medlemsstats lagstiftning är godkänd i överensstämmelse med detta direktiv.
2. Medlemsstaterna skall säkerställa att hela den praktiska utbildningen fullgörs hos personer som erbjuder tillräckliga garantier med avseende på utbildningen.
Artikel 9
Medlemsstaterna får tillåta personer att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna även om de inte uppfyller villkoren enligt artikel 4, under förutsättning att de kan visa a) att de under 15 år har utövat yrkesmässig verksamhet som har gett dem möjligheter att förvärva tillräcklig erfarenhet på ekonomi-, juridik- och redovisningsområdena samt har godkänts vid en sådan yrkesexamen som avses i artikel 4, eller
b) att de under sju år har utövat yrkesmässig verksamhet inom de angivna områdena och dessutom har erhållit praktisk utbildning enligt artikel 8 samt har godkänts vid en sådan yrkesexamen som avses i artikel 4.
Artikel 10
1. Medlemsstaterna får från de i artikel 9 angivna åren för yrkesmässig verksamhet räkna av tid för teoretisk utbildning inom de ämnesområden som anges i artikel 6, förutsatt att denna utbildning har avslutats med en statligt erkänd examen. Utbildningen får inte understiga ett år och får inte heller med mer än fyra år räknas av från tiden för yrkesmässig verksamhet.
2. Tiden för den yrkesmässiga verksamheten och den praktiska utbildningen får inte understiga tiden för den teoretiska och praktiska yrkesutbildning som har föreskrivits enligt artikel 4.
Artikel 11
1. Myndigheterna i en medlemsstat får godkänna personer som helt eller delvis har förvärvat sina kvalifikationer i någon annan stat, om dessa personer uppfyller följande två villkor: a) en behörig myndighet skall finna att deras kompetens är likvärdig med den som krävs enligt medlemsstatens lagstiftning i överensstämmelse med detta direktiv, och
b) de skall ha styrkt att de har sådana juridiska kunskaper som i medlemsstaten krävs för lagstadgad revision av de i artikel 1.1 angivna handlingarna. Myndigheterna i medlemsstaten behöver dock inte fordra att sådana kunskaper styrks, om myndigheterna finner att de juridiska kunskaper som har förvärvats i en annan stat är tillräckliga.
2. Artikel 3 skall tillämpas.
Artikel 12
1. En medlemsstat får anse sådana yrkesutövare som godkända enligt detta direktiv, vilka har godkänts genom ett förvaltningsbeslut av en behörig myndighet i den medlemsstaten innan de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas.
2. Inträder en fysisk person i en av staten erkänd yrkesförening får detta anses som ett godkännande genom förvaltningsbeslut av behörig myndighet enligt punkt 1, om inträdet enligt lagstiftningen i den staten ger föreningsmedlemmen rätt att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna.
Artikel 13
Till dess att de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas får en medlemsstat anse sådana yrkesutövare som godkända enligt detta direktiv, vilka visserligen inte har godkänts genom förvaltningsbeslut av en behörig myndighet men som dels har samma kvalifikationer i medlemsstaten som de personer vilka har godkänts genom sådana beslut och dels vid tidpunkten för dessa godkännanden utför lagstadgad revision av de i artikel 1.1 angivna handlingarna på de godkända personernas vägnar.
Artikel 14
1. En medlemsstat får anse sådana revisionsbolag som godkända enligt detta direktiv, vilka har godkänts genom förvaltningsbeslut av en behörig myndighet i den medlemsstaten innan de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas.
2. Villkoren enligt artikel 2.1 b ii och iii måste uppfyllas senast inom en tidsfrist som inte får överstiga fem år räknat från den tidpunkt då de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas.
3. Fysiska personer som till dess de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas utför lagstadgad revision av de i artikel 1.1 angivna handlingarna för ett revisionsbolags räkning, får därefter meddelas tillstånd att fortsätta att utföra sådan revision även om de inte uppfyller alla villkor i detta direktiv.
Artikel 15
Intill ett år efter den tidpunkt då de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas får de yrkesutövare som inte har godkänts genom förvaltningsbeslut av en behörig myndighet, men som i en medlemsstat ändå har rätt att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna och som faktiskt har utfört sådan revision fram till den nämnda tidpunkten, godkännas av medlemsstaten enligt detta direktiv.
Artikel 16
Artikel 18
1. I sex år räknat från den tidpunkt då de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas får medlemsstaterna vidta övergångsåtgärder för att reglera förhållandena för sådana personer som vid nämnda tidpunkt är i färd med sin teoretiska eller praktiska utbildning, men som då utbildningen avslutas inte skulle uppfylla de villkor som detta direktiv ställer upp och därför inte skulle få utföra den lagstadgade revision av de i artikel 1.1 angivna handlingarna för vilken de har utbildats.
2. Artikel 3 skall tillämpas.
Artikel 19
De i artikel 15 och 16 nämnda yrkesutövarna och de i artikel 18 nämnda personerna får med avvikelse från artikel 4 godkännas, endast om de enligt behöriga myndigheters uppfattning är lämpliga att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna och har kvalifikationer som är likvärdiga med dem som innehas av personer som godkänns enligt artikel 4.
Artikel 20
I avvaktan på en senare samordning av den lagstadgade revisionen av räkenskapshandlingar får en medlemsstat - som inte utnyttjar den i artikel 51.2 i direktiv 78/660/EEG angivna möjligheten och i vilken stat, då detta direktiv antas, flera kategorier fysiska personer enligt nationell lagstiftning är behöriga att utföra lagstadgad revision av de i artikel 1.1 a angivna handlingarna - särskilt godkänna fysiska personer som handlar i eget namn att utföra lagstadgad revision av de i artikel 1.1 a angivna handlingarna i bolag som inte överskrider gränserna för två av de tre kriterierna i artikel 27 i direktiv 78/660/EEG, om dessa personer: a) uppfyller de i artikel 3-19 i detta direktiv ställda villkoren, dock att nivån för yrkesexamen får vara lägre än vad som krävs enligt artikel 4, och
b) redan har utfört lagstadgad revision i det ifrågavarande bolaget, innan detta överskred gränserna för två av de tre kriterierna enligt artikel 11 i direktiv 78/660/EEG.
Om bolaget ingår i en grupp av företag vars räkenskaper skall sammanställas och som överskrider gränserna för två av de tre kriterierna i artikel 27 i direktiv 78/660/EEG, får dock inte sådana personer utföra lagstadgad revision i bolaget av de handlingar som anges i artikel 1.1 a i detta direktiv.
Artikel 21
I avvaktan på en senare samordning av den lagstadgade revisionen av räkenskapshandlingar får en medlemsstat - som inte utnyttjar den i artikel 6.1 i direktiv 83/349/EEG angivna möjligheten och i vilken stat, då detta direktiv antas, flera kategorier fysiska personer enligt nationell lagstiftning är behöriga att utföra lagstadgad revision av de i artikel 1.1 b angivna handlingarna - lämna särskilt tillstånd för en person som har godkänts enligt artikel 20 i detta direktiv att utföra lagstadgad revision av de i artikel 1.1 b angivna handlingarna, om på moderbolagets bokslutsdag den grupp av företag vars räkenskaper skall sammanställas sammanlagt enligt företagens senaste årsbokslut inte överskrider gränserna för två av de tre kriterierna i artikel 27 i direktiv 78/660/EEG, förutsatt att personen i fråga är behörig att utföra lagstadgad revision av de i artikel 1.1 a i detta direktiv angivna handlingarna i samtliga de företag som ingår i sammanställningen.
Artikel 22
En medlemsstat som tillämpar artikel 20 får i fråga om där avsedda personer tillåta att den i artikel 8 angivna praktiska utbildningen fullgörs hos någon som enligt den statens lagstiftning har godkänts att utföra sådan lagstadgad revision som avses i artikel 20.
AVSNITT III Yrkesmässig omsorg och oberoende
Artikel 23
Medlemsstaterna skall föreskriva att de personer som har godkänts att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna skall utföra revisionen med yrkesmässig omsorg.
Artikel 24
Medlemsstaterna skall föreskriva att dessa personer inte får utföra en lagstadgad revision, om de inte är oberoende enligt lagstiftningen i den medlemsstat som kräver revisionen.
Artikel 25
Artikel 23 och 24 skall även tillämpas på fysiska personer som uppfyller villkoren i artikel 3-19 och som utför lagstadgad revision av de i artikel 1.1 angivna handlingarna på ett revisionsbolags vägnar.
Artikel 26
Medlemsstaterna skall säkerställa att godkända personer blir föremål för lämpliga påföljder om de inte utför revisionen enligt artikel 23, 24 och 25.
Artikel 27
Medlemsstaterna skall säkerställa att i varje fall de aktieägare och andra delägare i godkända revisionsbolag samt de ledamöter i dessa bolags förvaltnings-, lednings- och övervakningsorgan, som i en medlemsstat inte personligen uppfyller villkoren enligt artikel 3-19, inte ingriper i revisionsarbetet på något sätt som äventyrar oberoendet hos de fysiska personer som på revisonsbolagens vägnar reviderar de i artikel 1.1 angivna handlingarna.
AVSNITT IV Offentliggörande
Artikel 28
1. Medlemsstaterna skall säkerställa att namn och adress för alla fysiska personer och revisionsbolag som av dem har godkänts att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna är offentligt tillgängliga.
2. Därutöver skall följande uppgifter om varje godkänt revisionsbolag vara offentligt tillgängliga: a) Namn och adress för de fysiska personer som anges i artikel 2.1 b i.
b) Namn och adress för aktieägare eller andra delägare i revisionsbolaget.
c) Namn och adress för ledamöter i revisionsbolagets företagsledning.
3. I de fall en fysisk person får utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna under de förutsättningar som anges i artikel 20, 21 och 22 skall punkt 1 i denna artikel tillämpas. Därvid skall emellertid anges i vilka kategorier av bolag och företagsgrupper som en sådan revision får utföras.
AVSNITT V Avslutande bestämmelser
Artikel 29
Den kontaktkommitté som har tillsatts enligt artikel 52 i direktiv 78/660/EEG skall även: a) med förbehåll för artikel 169 och 170 i Romfördraget underlätta en enhetlig tillämpning av detta direktiv genom regelbundet samråd, särskilt om praktiska problem i samband med tillämpningen,
b) vid behov ge kommissionen råd om tillägg till eller ändringar i detta direktiv.
Artikel 30
1. Medlemsstaterna skall före den 1 januari 1988 sätta i kraft de lagar och andra författningar som behövs för att följa detta direktiv. De skall genast underrätta kommissionen om det.
2. Medlemsstaterna får föreskriva att de i punkt 1 avsedda bestämmelserna skall tillämpas först från den 1 januari 1990.
3. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
4. Medlemsstaterna skall även till kommissionen överlämna förteckningar över examina som har anordnats eller erkänts i överensstämmelse med artikel 4.
Artikel 31
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(), senast ändrad genom förordning nr (EEG) nr 2260/84(), särskilt artikel 5.4 till denna,
med beaktande av kommissionens förslag, och
med beaktande av följande: Genom artikel 5 i förordning nr 136/66/EEG införs en form av produktionsstöd för olivolja. Detta stöd för områden som är planterade med olivträd på ett visst datum beviljas odlare som är medlemmar av de producentorganisationer som anges i artikel 20c.1 i förordning nr 136/66/EGG och vars genomsnittliga produktion är minst 100 kg olja per regleringsår och till andra odlare på grundval av antalet olivträd samt produktionspotentialen och avkastningen från dessa träd, fastställd enligt en standardmetod, och under förutsättning att de odlade oliverna verkligen har skördats.
I avvaktan på upprättandet av ett register för olivodling, bör stödet till de berörda odlarna beräknas på grundval av den genomsnittliga avkastningen av olivträd.
För att säkerställa att stödsystemet fungerar på rätt sätt är det nödvändigt att bestämma för vilka typer av olivolja stöd skall beviljas.
För att säkerställa att stödsystemet fungerar på rätt sätt bör rättigheterna och skyldigheterna för alla berörda parter, nämligen odlare, producentorganisationer och sammanslutningar av producentorganisationer samt de berörda medlemsstaterna, fastställas.
De sammanslutningar av organisationer för olivoljeproducenter som avses i artikel 20c.2 i den förordningen bör bestå av ett minimiantal av grupper eller representera en minsta procentuella andel av den inhemska produktionen. Dessa minsta antal eller andelar bör fastställas på en nivå som gör det möjligt att utföra det speciella samordnings- och kontrollarbete som dessa sammanslutningar är skyldiga att utföra på ett effektivt sätt.
I artikel 20c i den förordningen anges att producentorganisationer och sammanslutningar av producentorganisationer bör utföra vissa kontroll- och samordningsuppgifter. Dessa uppgifter bör därför exakt anges.
För att förvaltningen skall fungera på rätt sätt skall producentorganisationer och sammanslutningar av dessa hos de behöriga nationella myndigheterna ansöka om godkännande i god tid före regleringsårets början. Den behöriga medlemsstaten bör besluta om dessa ansökningar inom en skälig tid.
Enligt artikel 20d.1 i den förordningen får en del av stödbeloppet behållas för att täcka de utgifter som producentorganisationer och sammanslutningar av dessa ådrar sig för att utföra kontrollarbetet. Åtgärder bör vidtas för att säkerställa att dessa belopp endast används för att betala för de arbetsuppgifter som avses i artiklarna 20c.1 och 20c.2 i den förordningen.
Artikel 20d.2 i den förordningen fastställer att endast sammanslutningar skall vara berättigade till förskottsbetalning av stödbeloppet. För att förvaltningen skall skötas på ett riktigt sätt bör detta förskott inte överstiga en viss procentuell andel av stödet.
För att säkerställa att systemet med produktionsstöd till odlare som tillhör producentorganisationer fungerar på rätt sätt, bör bestämmelser införas om att stöd endast bör utbetalas för de kvantiteter som erhålls från godkända fabriker. För att bli godkända bör fabrikerna i fråga uppfylla flera villkor.
Ifrågavarande stöd är till stor fördel för oljeproducenterna och utgör en finansiell börda för gemenskapen. För att säkerställa att stödet endast beviljas för olja som är berättigad till det, bör bestämmelser fastställas om inrättandet av ett lämpligt system för administrativa kontroller.
För att stödsystemet skall fungera på rätt sätt, bör medlemsstaterna bestämma vilken kvantitet av olja som är berättigad till stöd i de fall då den verkliga produktionen av olivolja är oklar.
Erfarenheten har visat, att trots de många särskilda kontroller som införts är en noggrann och effektiv kontroll och verifiering svår att genomföra, på grund av det stora antalet odlare som skall kontrolleras. Dessa svårigheter måste lösas genom att ett dataregister upprättas i varje medlemsstat som innehåller all nödvändig information för att underlätta kontrollen och snabbt upptäcka oegentligheter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Från och med regleringsåret 1984/1985 skall de allmänna bestämmelser som fastställs i denna förordning tillämpas vid beviljande av produktionsstöd för olivolja enligt artikel 5 i förordning nr 136/66/EEG.
3. Stödet skall beviljas efter ansökan från de berörda parterna till den medlemsstat i vilken oljan har framställts.
4. För olivodlare som är medlemmar i en producentorganisation enligt artikel 20c.1 i förordning nr 136/66/EEG och vars normala produktion inte är mindre än 100 kg olivolja per regleringsår, skall stödet beviljas enligt artikel 5.2 första strecksatsen i den förordningen för den kvantitet olja som verkligen framställts vid en godkänd fabrik, om inte annat följer av artikel 7.
För andra olivodlare skall stödet beviljas enligt artikel 5.2 andra strecksatsen i förordning nr 136/66/EEG, och stödet skall motsvara det stöd som erhålls om avkastningen från oliver och olivolja, fastställd enligt den standardmetod enligt artikel 18, tillämpas för antalet olivträd i produktion.
5. För regleringsåren 1984/85 och 1985/86 skall de producerande medlemsstaterna bestämma vilka olivodlare, med en genomsnittlig produktion av minst 100 kg olja per regleringsår, som är berättigade att erhålla stöd, beviljat efter den kvantitet av olja som verkligen har framställts, genom användning av avkastningen av oliver och olivolja fastställd enligt artikel 18, i förhållande till antalet olivträd i produktionen.
6. Före den 31 mars 1986 skall rådet med kvalificerad majoritet på förslag av kommissionen fastställa de kriterier som skall tillämpas från och med regleringsåret 1986/87 vid bestämmande av de olivodlare som normalt framställer minst 100 kg olja per regleringsår.
Artikel 3
1. Varje olivodlare skall vid början av regleringsåret och före en fastställd dag till de behöriga myndigheterna i medlemsstaten i fråga inge en skördedeklaration, som vid första tillfället det inges skall innehålla:
- närmare uppgifter om de olivträd som odlas och var de finns,
- en kopia av den deklaration som lämnats för sammanställning av registret över olivodling. Denna deklaration får, när det gäller Grekland och till dess att registret över olivodling är sammanställt i den medlemsstaten, ersättas av den deklaration som anges i artikel 1.1 i förordning (EEG) nr 1590/83.
2. Under de följande regleringsåren skall varje olivodlare, före en dag som skall fastställas, inge en kompletterande deklaration, i vilken odlaren uppger alla förändringar som har skett eller att den tidigare lämnade skördedeklarationen fortfarande är tillämplig.
3. Olivodlare som är medlemmar i en producentorganisation skall, på en dag som skall fastställas, till den organisation som de tillhör lämna en ansökan om individuellt stöd med ett bevis på att oliverna är pressade eller bearbetade, eller en faktura för oliverna eller båda dokumenten.
4. De olivodlare som avses i punkt 3 skall lämna skördedeklarationen och ansökan om stöd via sin organisation.
Producentorganisationerna skall till den behöriga medlemsstaten anmäla namnen på de olivodlare som avses i andra stycket.
6. För de olivodlare som inte är medlemmar i en producentorganisation skall den inlämnade individuella skördedeklarationen anses som en ansökan om stöd, förutsatt att den före en dag som skall fastställas kompletteras med:
- en deklaration om att de har skördat sina oliver för regleringsåret i fråga, och
- upplysningar om den avsedda användningen av oliverna.
7. Olivodlare som försummar att uppfylla förpliktelserna i denna artikel skall inte beviljas stöd.
Artikel 4
1. Med beaktande av de andra kraven i artikel 20c.1 i förordning nr 136/66/EEG får en producentorganisation inte godkännas enligt den förordningen om den inte
a) i fråga om organisationer som producerar och ökar marknadsvärdet av oliver och olivolja, består av minst 700 olivodlare, eller
b) i övriga fall, består av minst 1 200 olivodlare. Skulle en eller flera organisationer som producerar och ökar marknadsvärdet av oliver och olivolja vara medlemmar i organisationen i fråga, skall de berörda odlarna beaktas individuellt vid beräkning av det minsta antalet odlare som fordras, eller
c) företräder minst 25 % av olivodlarna eller produktionen av olivolja i den ekonomiska region där den har upprättats.
2. Endast olivodlare med följande kännetecken får tillhöra en organisation: olivodlare som äger en olivodling som de brukar eller olivodlare som har brukat en olivodling under minst tre år.
För att uppnå detta skall olivodlare överlämna de upplysningar som behövs till de producentorganisationer som de tillhör för att fastställa att de brukar en olivodling samt uppgifter om alla förändringar som skett sedan de ansökte om medlemsskap.
3. I detta direktiv avses med ekonomisk region ett område som, enligt kännetecken som skall fastställas av den berörda medlemsstaten, har likartade produktionsvillkor med avseende på olivodling.
4. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att uppmuntra inrättandet av de producentgrupper som anges i förordning (EEG) nr 1360/78 () eller andra organisationer för att framställa och öka marknadsvärdet av oliver och olivolja, vilka kan godkännas som producentorganisationer enligt denna förordning.
Artikel 5
1. Producentorganisationer som önskar bli erkända från början av ett regleringsår skall ansöka hos den behöriga myndigheten i medlemsstaten i fråga senast den 30 juni under det föregående regleringsåret.
2. Senast den 15 oktober skall den behöriga myndigheten, efter att ha mottagit ansökan, fatta beslut om denna efter att ha kontrollerat, om organisationen uppfyller kraven enligt artikel 20c.1 i förordning nr 136/66/EEG och enligt artikel 4, och genast anmäla detta till den berörda organisationen och till kommissionen.
Tillståndet skall träda i kraft från början av det regleringsår som följer efter ansökningsåret.
3. Godkända producentorganisationer skall senast den 30 juni varje år anmäla alla ändringar som skett i deras organisationer efter deras godkännande eller sedan den sista årliga deklarationen inlämnades och anmäla alla mottagna återkallelser av eller ansökningar om medlemskap till den behöriga myndigheten.
Den behöriga myndigheten skall på grundval av denna anmälan och andra lämpliga undersökningar förvissa sig om att villkoren för godkännande fortfarande är uppfyllda.
Om villkoren inte längre uppfylls eller om organisationens struktur inte gör det möjligt att kontrollera medlemmarnas produktion, skall den behöriga myndigheten snarast och senast före det följande regleringsårets början återkalla godkännandet och anmäla sitt beslut om detta till kommissionen.
Artikel 6
1. Godkända producentorganisationer skall
- lämna in skördedeklarationer från alla sina medlemmar enligt artikel 3.1,
- utföra kontroller på plats av de upplysningar som lämnats, i en viss del av dessa deklarationer, vilken skall fastställas,
- en gång i månaden överlämna medlemmarnas ansökningar om stöd i ett standardformat som kan användas vid den databearbetning som anges i artikel 16. Stöd skall begäras för den kvantitet som framställts av de medlemmar som har avslutat sin oljeproduktion, förutsatt att de kontroller som anges i artikel 8 har utförts och att de skyldigheter som följer av dessa har uppfyllts.
Alla ansökningar som gäller produktionen från ett enda regleringsår skall, med risk för uteslutning, inlämnas före en fastställd dag.
2. Om en producentorganisation tillhör en sammanslutning av dessa organisationer, skall skördedeklarationerna och ansökningarna om stöd från de olivodlare som är medlemmar överlämnas av sammanslutningen.
Artikel 7
Den kvantitet av olja för vilken stöd erhålls får inte vara större än den kvantitet som fastställs genom standardmetoden enligt artikel 18, dvs. att den fastställda skörden av oliver och olja tillämpas för antalet olivträd i produktionen, om en olivodlare som är medlem i en producentorganisation
- även har arrenderat olivodlingar för mindre än tre år,
- har sålt antingen delar av eller hela sin produktion av olja, och
- har blivit medlem i organisationen under regleringsåret.
Artikel 8
1. Varje producentorganisation skall, före överlämnandet av ansökningan om stöd, kontrollera den kvantitet av olivolja för vilken stöd söks för var och en av dess medlemmar. Organisationen skall särskilt kontrollera:
- att den produktion av oliver, av varje odlare deklarerad som pressad i en godkänd fabrik, stämmer överens med de uppgifter som lämnats i hans skördedeklaration, på grundval av kännetecken som skall fastställas,
- att de uppgifter som lämnats av varje odlare i fråga om de kvantiteter av oliver som pressats och de kvantiteter av olja som erhållits stämmer överens med de kvantiteter av oliver och olja som uppgivits i bokföringen hos de godkända fabrikerna.
2. Producentorganisationer skall överlämna sina medlemsregister till de behöriga myndigheterna i den berörda medlemsstaten i följande fall:
- Om de upplysningar som anges i punkt 1 första strecksatsen inte förefaller att stämma överens, efter det att organisationen har erhållit alla stöddokument och alla upplysningar som kan användas för att fastställa den kvantitet som verkligen producerats.
- Om de upplysningar som anges i punkt 1 andra strecksatsen inte förefaller att stämma överens.
- Om upplysningarna i skördedeklarationen inte stämmer med vad som framkommit vid kontrollerna.
Artikel 9
1. Med beaktande av kraven i artikel 20c.2 i förordning nr 136/66/EEG får en sammanslutning inte godkännas om den inte består av minst 10 producentorganisationer, godkända enligt artikel 5, eller ett antal organisationer som svarar för minst 5 % av den olivolja som framställs i den berörda medlemsstaten.
De producentorganisationerna som innefattas i en sammanslutning skall dock komma från minst två ekonomiska regioner.
2. Bestämmelserna om godkännande och återkallande av godkännande enligt vad som anges i artikel 5 skall även tillämpas för sammanslutningar. Artikel 10
De sammanslutningar som avses i artikel 20c.2 i förordning nr 136/66/EEG
- skall samordna arbetet i de organisationer som de består av och säkerställa att detta arbete är förenligt med bestämmelserna i denna förordning och skall framförallt snarast kontrollera, enligt ett procenttal som skall bestämmas, på vilket sätt de kontroller som anges i artiklarna 6 och 8 har genomförts,
- skall överlämna de skördedeklarationer och ansökningar om stöd som inlämnats till dem av de organisationer som de består av till de behöriga myndigheterna,
- skall ta emot förskott av produktionsstödet, såsom anges i artikel 12, och saldot på stödbeloppen från den berörda medlemsstaten och skall snarast dela upp dem mellan de producenter som är medlemmar i de organisationer som tillhör dem.
Artikel 11
1. Det belopp som innehållits enligt artikel 20d.1 i förordning nr 136/66/EEG skall användas på följande sätt:
a) Ett belopp som skall fastställas skall utbetalas till varje sammanslutning på grundval av antalet medlemmar i de producentorganisationer som tillhör den.
b) Saldot skall utbetalas till alla producentorganisationer på grundval av
- antalet individuella ansökningar om stöd som inges till varje organisation av dess medlemmar,
- kontroller som utförts enligt förfarandet för erhållande av stöd.
2. De medlemsstater i vilka olivolja framställs skall garantera att de summor som överlämnats till sammanslutningarna och producentorganisationerna vid tillämpningen av punkt 1 endast används av dem för att finansiera den verksamhet som de är ansvariga för enligt denna förordning.
3. Om beloppen inte används, helt eller delvis, såsom anges i punkt 2 skall de återbetalas till den behöriga medlemsstaten och avräknas från de utgifter som finansieras av EUGFJ.
4. För att underlätta verksamheten i sammanslutningar och producentorganisationer är medlemsstaterna behöriga att i början av varje regleringsår betala dem ett förskott, som skall beräknas på grundval av en enhetstaxa för antalet medlemmar.
5. De producerande medlemsstaterna skall fastställa bestämmelser om tilldelningen av stödbelopp och tidsbegränsningar för betalning till olivodlare.
Artikel 12
1. De producerande medlemsstaterna skall ha rätt att till sammanslutningar av producentorganisationer utbetala ett förskott på de yrkade stödbeloppen.
2. Under regleringsåren 1984/1985, 1985/1986 samt 1986/1987 skall det förskott som avses i punkt 1 till varje odlare inte överstiga
- det belopp som erhålls genom tillämpning av skörden av oliver och olja, fastställd enligt artikel 18, för antalet olivträd i produktion enligt skördedeklarationen eller det belopp som erhålls för den uppgivna kvantiteten i ansökan, om den kvantiteten är mindre än den som anges ovan, eller
- 50 % av det belopp som erhålls vid beräkning av ett genomsnitt av de stödbelopp som betalats under de två föregående regleringsåren.
Artikel 13
1. Medlemsstaterna skall endast godkänna fabriker vars ägare
a) till medlemsstaten i fråga, enligt bestämmelser som skall fastställas, har överlämnat fullständiga upplysningar om fabrikens tekniska utrustning och nuvarande pressningskapacitet samt alla ändringar av dessa uppgifter,
b) har samtyckt till att genomgå alla kontroller som föreskrivs enligt stödförfarandet och till att godkänna alla kontroller som anses nödvändiga i sina lokaler samt att tillåta alla kontroller av deras bokföring,
c) under det föregående regleringsåret inte blivit föremål för åtgärder beroende på oriktigheter som upptäckts vid kontroller enligt artikel 14 och denna artikel, beträffande godkännande för regleringsåret 1984/1985,
- inte blivit föremål för åtgärder rörande oriktigheter som upptäckts vid kontroller gjorda för regleringsåret 1983/1984 enligt artikel 7 och 9 i förordning (EEG) nr 2959/82(), och
- inte har fått sitt godkännade indraget för en tid som sträcker sig efter den 31 oktober 1984 enligt den förordningen,
d) samtycka till att föra en standardiserad lagerredovisning enligt kriterier som skall fastställas.
2. Medlemsstaterna skall innan de beviljar ett godkännande kontrollera om villkoren för ett godkännande är uppfyllda och skall särskilt på platsen kontrollera den tekniska utrustningen och den faktiska pressningskapaciteten i fabrikerna.
3. Under regleringsåren 1984/1985 och 1985/1986 får de berörda medlemsstaterna bevilja tillfälligt godkännande till den berörda fabriken, så snart en ansökan om godkännande innehållande de upplysningar som anges i punkt 1 har överlämnats.
Detta tillfälliga godkännande skall bli definitivt så snart den berörda medlemsstaten har förvissat sig om att de villkor för godkännande som fastställs i punkt 1 är uppfyllda.
Om det visar sig att ett av de villkor som anges i punkt 1 inte är uppfyllt, skall det tillfälliga godkännandet återkallas.
4. I de fall då ett av villkoren för godkännande enligt punkt 1 inte längre är uppfyllt skall godkännandet återkallas för den tid som är beroende av hur allvarlig överträdelsen är.
5. I de fall godkännandet återkallas i enlighet med punkt 3 eller 4 får ingen ny ansökan om godkännande under den tid då godkännandet är återkallat beviljas.
- samma fysiska eller juridiska person som förestår fabriken i fråga,
eller - någon fysisk eller juridisk person som önskar förestå fabriken i fråga, om inte den personen tillfredsställande kan bevisa för den berörda medlemsstaten att ansökan om nytt godkännande inte är ämnad att kringgå den påförda sanktionen.
Artikel 14
1. Varje producerande medlemsstat skall tillämpa ett kontrollsystem för att säkerställa att den produkt för vilken stöd beviljas är berättigad till detta stöd.
2. Producerande medlemsstater skall kontrollera verksamheten i varje producentorganisation och sammanslutning och framförallt kontrollera att kontrollförfarandena har genomförts av dessa organ.
3. Under varje regleringsår och framför allt under den tid då oljan pressas, skall de producerande medlemsstaterna på plats kontrollera verksamheten och bokföringen hos en viss procent av de godkända fabrikerna, vilken skall fastställas.
De utvalda fabrikerna skall vara representativa för pressningskapaciteten i ett produktionsområde.
4. Om den olivolja som anges i punkt 1 i bilagan till förordning nr 136/66/EEG framställts av odlare som inte är medlemmar i en producentorganisation, skall kontrollen innebära provtagning på plats som skall bekräfta
- att skördedeklarationerna är riktiga,
- att de skördade oliverna skall användas för att framställa olja och, om möjligt, att de faktiskt har bearbetats till olja.
Kontrollerna skall ske hos en procentuell andel av odlarna och denna andel skall fastställas på grundval av framför allt företagens storlek.
5. Medlemsstaterna skall bl. a. använda de dataregister som föreskrivs i artikel 16 för dessa kontroller och verifieringar.
Dessa register skall användas som stöd i den kontrollverksamhet som skall förekomma enligt punkt 1 4.
Artikel 15
1. Medlemsstaterna skall besluta vilken kvantitet av olja är berättigad till stöd på grundval av de ansökningar som överlämnas enligt artiklarna 3 och 6, med hänsyn tagen till alla dithörande fakta och särskilt till alla kontroller och godkännanden som föreskrivs i denna förordning.
Den kvantitet olivolja som avses i punkt 4 i bilagan till förordning nr 136/66/EEG för vilken stöd får medges skall bestämmas på grundval av den typ av olja som anges i punkt 1 i den bilagan.
2. För producenter vars bokföringsuppgifter har överlämnats till medlemsstaten av deras organisationer enligt artikel 8.2 skall medlemsstaten besluta för vilken kvantitet av olja stödet skall ges. 3. Om resultaten av de kontroller som anges i artiklarna 13 och 14 inte överensstämmer med uppgifterna i lagerbokföringen i en godkänd fabrik, skall den ifrågavarande medlemsstaten, med beaktande av alla sanktioner som får åläggas fabriken, fastställa den kvantitet olja för vilken stöd får beviljas för varje producent som är medlem i en organisation som har pressat sin olivskörd i fabriken i fråga.
4. Som underlag för bestämmandet av den kvantitet som är berättigad till stöd, i de fall som omfattas av punkt 2 och 3, skall medlemsstaten framför allt använda skörden av oliver och olja, fastställd enligt den standardmetod som anges i artikel 18.
Artikel 16
1. Varje producerande medlemsstat skall upprätta och underhålla permanenta dataregister innehållande uppgifter om produktionen av oliver och olivolja.
2. Dessa register skall innehålla minst följande information:
a) För varje olivodlare och för varje regleringsår som en ansökan om stöd har inlämnats
- de upplysningar som finns i den skördedeklaration som föreskrivs i artikel 3.
- de kvantiteter av producerad olja, för vilka en ansökan om produktionsstöd har inlämnats samt den kvantiteten för vilken stöd har utbetalats,
- uppgifter som erhållits vid de kontroller på plats som gjorts hos olivodlaren.
b) För producentorganisationer och sammanslutningar av dessa: all information som behövs för att kontrollera deras verksamhet i samband med det nuvarande stödsystemet samt även resultaten av de kontroller som utförts av medlemsstaterna.
c) För fabriker som framställer olivolja och för varje regleringsår: de uppgifter som finns i lagerbokföringen, information om den tekniska utrustningen och pressningskapaciteten samt resultaten av de kontroller som utförts enligt denna förordning.
d) De förväntade årliga skördarna för varje enhetligt produktionsområde.
Artikel 17
1. De register som anges i artikel 16 skall vara konfidentiella.
Följande organ skall ha tillgång till dem:
- De nationella myndigheter som är bemyndigade av medlemsstaten.
- Kommissionens tjänstemän i samarbete med de behöriga tjänstemännen i medlemsstaterna och enligt förordning (EEG) nr 729/70(), senast ändrad genom förordning (EEG) nr 3509/80(), särskilt med tanke på de fastställda förfarandena.
- Producentorganisationer och sammanslutningar av dessa, i fråga om de aspekter som medlemsstaterna anser vara nödvändiga för att effektivt kontrollera sina respektive medlemmar.
2. De dataregister som upprättas och de program som används för att hantera dem skall vara kompatibla med de datasystem som används för registrering av olivodlingen i varje producerande medlemsstat.
Artikel 18
De skördar av oliver och olja som anges i artikel 5.2 första stycket andra strecksatsen i förordning nr 136/66/EEG skall fastställas för enhetliga produktionsområden, senast den 31 maj varje år på grundval av uppgifter som de producerande medlemsstaterna lämnar senast den 30 april varje år.
Artikel 19
Tillämpningsföreskrifter för denna förordning skall antas enligt förfarandet i artikel 38 i förordning nr 136/66/EEG.
Följande uppgifter skall fastställas enligt samma förfarande:
- De skördar som anges i artikel 18.
- De belopp som anges i artikel 11.1 a.
Artikel 20
För att möjliggöra en smidig övergång från den gällande ordningen till den som fastställs enligt denna förordning, får kommissionen besluta om nödvändiga åtgärder för regleringsåret 1984/85, enligt förfarandet i artikel 38 i förordning nr 136/66/EEG.
Artikel 21
Före slutet av det tredje året under vilket denna förordning tillämpas skall kommissionen överlämna en rapport till rådet om den verksamhet som fastställs i denna förordning tillsammans med förslag om hur rådet skall ändra verksamheten.
Artikel 22
Medlemsstaterna skall anmäla de åtgärder som genomförs enligt denna förordning till kommissionen.
Artikel 23
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag(),
med beaktande av Europaparlamentets yttrande(),
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
med beaktande av följande: I syfte att göra hälsoskyddsåtgärderna enhetliga för konsumenterna fastställs bestämmelser i direktiv 64/433/EEG(), senast ändrat genom direktiv 83/90/EEG() om hygienundersökningar och kontroller av färskt kött som kan komma att införas i handeln inom gemenskapen.
För att skydda människors och djurs hälsa inom gemenskapen har man i direktiv 72/462/EEG(), senast ändrat genom direktiv 83/91/EEG(), fastställt att medlemsstaternas behöriga myndigheter skall utföra hygienundersökningar vid import av färskt kött och att veterinära experter från medlemsstaterna och kommissionen skall genomföra inspektioner inom det exporterande tredje landet.
Bestämmelserna i direktiv 64/433/EEG omfattar endast färskt kött som kan komma att föras i handel inom gemenskapen. Medlemsstaternas myndigheter har dock infört nationella kontroller av färskt kött som enbart är avsett för den nationella marknaden.
Rådets direktiv 71/118/EEG(), senast ändrat genom direktiv 84/642/EEG() föreskriver att hälsoundersökningar och kontroller skall ske av färskt fjäderfäkött.
I samband med dessa hälsoundersökningar och kontroller debiteras avgifter som för närvarande finansieras på olika sätt i de skilda medlemsstaterna. Dessa skillnader kan påverka de konkurrensvillkor som råder för produkter som till största delen omfattas av en gemensam marknadsordning.
För att undanröja sådana skillnader bör harmoniserade regler fastställas för finansieringen av dessa hygienundersökningar och kontroller.
Med hänsyn till nationella förvaltnings- och finansieringsbestämmelser och -förfaranden bör en ytterligare frist på två år beviljas för att göra det möjligt för Grekland att införa det nödvändiga systemet för att ta ut avgifter i samband med undersökningar och kontroller.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Medlemsstaterna skall säkerställa att man från och med den 1 januari 1986
P tar ut avgifter för att täcka kostnaderna för hygienundersökningar och kontroller när ett djur enligt punkt 2 slaktas,
P för att dels säkerställa lika behandling enligt artikel 15 i direktiv 71/118/EEG och dels täcka de omkostnader som avses i direktiv 72/462/EEG tar ut en avgift för det kött som avses i dessa direktiv och som importeras från tredje land,
P förbjuder varje form av direkt eller indirekt återbetalning av avgifter.
1. Rådet skall på förslag av kommissionen och med kvalificerad majoritet före den 1 januari 1986, fatta beslut om den eller de avgiftsbelopp som avses i artikel 1.1 de första två strecksatserna och om principer och tillämpningsföreskrifter för detta direktiv, samt om möjliga undantag. De avgiftsbelopp som skall debiteras för kött som kommer från slakterier som inte har godkänts enligt direktiv 64/433/EEG skall däremot inte fastställas förrän i samband med att rådet före detta datum har antagit bestämmelser om undersökning av detta kött.
2. Medlemsstaterna kan debitera en summa som överstiger den eller de belopp som avses i punkt 1, under förutsättning att den sammanlagda avgift som uttas i varje medlemsstat är lägre än eller lika med de faktiska kostnaderna för undersökningarna.
Artikel 3
Kommissionen skall före den 1 januari 1990 överlämna en rapport om vunna erfarenheter tillsammans med eventuella förslag till ändringar av de ovannämnda artiklarna.
Artikel 4
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 1986. De skall genast underätta kommissionen om detta.
Grekland skall dock ha en ytterligare tidsfrist på två år för att följa det.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av kommissionens förslag(),
med beaktande av Europaparlamentets yttrande(),
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
med beaktande av följande: Enligt fördraget är all särbehandling som grundar sig på nationalitet när det gäller etablering och tillhandahållande av tjänster förbjuden fr.o.m. övergångsperiodens utgång. Principen om sådan behandling som grundar sig på nationalitet förekommer särskilt vid beviljande av de tillstånd som krävs för att utöva vissa former av verksamhet samt inregistrering eller medlemskap i yrkesorganisationer eller motsvarande organ.
Det förefaller ändå önskvärt att vissa bestämmelser införs för att underlätta det faktiska utövandet av etableringsrätten.
Enligt artikel 54.3 h i fördraget får medlemsstaterna inte bevilja någon form av stödåtgärder som skulle kunna snedvrida etableringsvillkoren.
Som villkor för att få utöva viss farmaceutisk verksamhet krävs i några medlemsstater förutom utbildnings-, examens- och andra behörighetsbevis en kompletterande yrkeserfarenhet; då det ännu inte föreligger någon överensstämmelse mellan medlemsstaterna inom detta område bör, för att undvika svårigheter, lämplig praktisk yrkeserfarenhet av samma längd som förvärvats i en annan medlemsstat erkännas som tillräcklig.
Inom ramen för ländernas hälso- och sjukvårdspolitik, som bl.a. går ut på att garantera en tillfredsställande utlämning av läkemedel överallt inom respektive lands territorium, begränsar vissa medlemsstater antalet nya apotek som får inrättas medan det i andra länder inte finns några bestämmelser av detta slag; under dessa omständigheter är det för tidigt att bestämma att följderna av ett erkännande av utbildnings-, examens- och andra behörighetsbevis i farmaci även skall omfatta utövandet av apotekarverksamhet som innehavare av ett apotek som varit öppet för allmänheten mindre än tre år; detta problem skall inom en viss bestämd tidsfrist utredas på nytt av kommissionen och rådet.
Då ett direktiv om ömsesidigt erkännande av examensbevis inte nödvändigtvis innebär likvärdighet när det gäller den utbildning som dessa examensbevis avser, bör rätten att använda yrkestitlar på grundval av utbildningen endast vara tillåten på språket i ursprungslandet eller det senaste hemvistlandet.
För att underlätta tillämpningen av detta direktiv för de nationella myndigheterna får en medlemsstat föreskriva att den person som uppfyller utbildningsvillkoren enligt detta direktiv samtidigt med de formella utbildningsbevisen skall förete ett intyg från de behöriga myndigheterna i ursprungslandet eller det senaste hemvistlandet som visar att dessa bevis är de som avses i direktivet.
Detta direktiv påverkar inte medlemsstaternas lagar eller författningar med bestämmelser som förbjuder bolag att utöva vissa former av verksamhet eller ålägger dem vissa villkor för detta.
Det är svårt att bedöma i vad mån föreskrifter i syfte att underlätta farmaceuters frihet att tillhandahålla tjänster f.n. kan vara till nytta; under nuvarande omständigheter bör några föreskrifter därför inte antas.
När det gäller kraven på god vandel och gott anseende bör skillnad göras mellan de krav som ställs för att påbörja verksamhet inom yrket och de krav som ställs för att få utöva yrket.
När det gäller verksamhet som anställd fastslås inte några särskilda bestämmelser i rådets förordning (EEG) nr 1612/68 av den 15 oktober 1968 om arbetskraftens fria rörlighet inom gemenskapen som hänför sig till god vandel eller gott anseende, yrkesansvar eller användningen av yrkestitlar(); beroende på den enskilda medlemsstaten tillämpas eller får dessa regler tillämpas på såväl anställda som självständigt verksamma yrkesutövare; sådan verksamhet för vilken det i alla medlemsstater krävs innehav av utbildnings-, examens- eller andra behörighetsbevis i farmaci utövas av såväl anställda som självständigt verksamma yrkesutövare eller av samma personer omväxlande som anställd eller som självständigt verksam yrkesutövare under deras yrkeskarriär; för att i möjligaste mån uppmuntra dessa yrkesutövares fria rörlighet inom gemenskapen förefaller det nödvändigt att utvidga detta direktiv till att även omfatta anställda.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 2
1. Varje medlemsstat skall erkänna de utbildnings-, examens- och andra behörighetsbevis som tilldelas medborgare i medlemsstaterna av övriga medlemsstater i enlighet med artikel 2 i direktiv 85/432/EEG och som finns uppräknade i artikel 4 genom att ge dessa bevis, när det gäller rätten att påbörja och utöva sådan verksamhet som avses i artikel 1, samma innebörd inom sitt territorium som dem som medlemsstaten själv utfärdar.
2. Medlemsstaterna är emellertid inte skyldiga att låta de utbildnings-, examens- och andra behörighetsbevis som avses i punkt 1 träda i kraft när det gäller att inrätta nya apotek som är öppna för allmänheten. Vid tillämpningen av detta direktiv skall apotek som varit i drift kortare tid än tre år betraktas som nyinrättade.
Fem år efter utgången av den tidsfrist som fastställts i artikel 19.1 skall kommissionen lägga fram en rapport för rådet om det sätt på vilket medlemsstaterna har tillämpat föregående stycke och om möjligheten att utvidga verkningarna av ett ömsesidigt erkännande av de utbildnings-, examens- och andra behörighetsbevis som avses i punkt 1. Den skall föreslå lämpliga åtgärder.
Artikel 3
1. Utan hinder av artikel 2 och utan att det påverkar tillämpningen av artikel 45 i 1979 års anslutningsakt skall Grekland endast åläggas att tillämpa bestämmelserna i artikel 2 om de utbildnings-, examens- och andra behörighetsbevis som utfärdas av de övriga medlemsstaterna, såvida det gäller utövande av de former av verksamhet som avses i artikel 1 som anställd i enlighet med förordning (EEG) nr 1612/68.
Så länge som Grekland använder denna undantagsbestämmelse och utan att det påverkar tillämpningen av artikel 45 i 1979 års anslutningsakt skall de övriga medlemsstaterna endast åläggas att tillämpa bestämmelserna i artikel 2 om de examensbevis som avses i artikel 4 d, såvida det gäller utövande av de former av verksamhet som avses i artikel 1 som anställd i enlighet med förordning (EEG) nr 1612/68.
2. Tio år efter utgången av den tidsfrist som fastställts i artikel 19 skall kommissionen föreslå rådet lämpliga åtgärder för att utvidga verkningarna av ett ömsesidigt erkännande av utbildnings-, examens- och andra behörighetsbevis i syfte att underlätta det faktiska utövandet av etableringsrätten mellan Grekland och de övriga medlemsstaterna. Rådet skall vidta åtgärder med anledning av dessa förslag i enlighet med det förfarande som fastställts i fördraget.
Artikel 4
De utbildnings-, examens- och andra behörighetsbevis som avses i artikel 2 är följande:
a) I Belgien:
Le diplôme légal de pharmacien/het wettelijk diploma van apoteker (det lagstadgade examensbeviset i farmaci) som utfärdas av universitetens medicinska och farmaceutiska fakulteter, av centrala examensnämnden eller av de statliga examensnämnderna för universitetsutbildningen.
b) I Danmark:
Bevis for bestået farmaceutisk kandidateksamen (intyg över genomgången farmaceutisk universitetsexamen).
c) I Tyskland:
1) Zeugnis über die staatliche Pharmazeutische Prüfung (statligt examensbevis för farmaceuter) som utfärdas av de behöriga myndigheterna,
2) Intyg från de behöriga myndigheterna i Tyskland som visar att de examensbevis som utfärdats efter den 8 maj 1945 av de behöriga myndigheterna i Tyska Demokratiska Republiken erkänns som likvärdiga med dem som avses i punkt 1 ovan.
d) I Grekland:
Ðéáôïðïéçôéêü ôùí áñìïäßùí áñ÷þí, éêáíüôçôáò Üóêçóçò ôçò öáñìáêåõôéêÞò, ÷ïñçãïýìåíï ìåôÜ êñáôéêÞ åîÝôáóç (det intyg som visar att innehavaren av detta är behörig att utöva verksamhet som farmaceut) som utfärdas av de behöriga myndigheterna efter statsexamen;
e) I Frankrike:
Statligt examensbevis som utfärdas av universiteten eller statligt examensbevis som farmacie doktor som utfärdas av universiteten.
f) I Irland:
Intyg som Registered Pharmaceutical Chemist.
g) I Italien:
Examensbevis eller intyg som innebär rätt att utöva verksamhet som farmaceut och som förvärvas efter statsexamen.
h) I Luxemburg:
Statligt examensbevis som farmaceut som utfärdas av statens examensnämnd och undertecknas av utbildningsministern.
i) I Nederländerna:
Het getuigschrift van med goed gevolg afgelegd apothekersexamen (bevis över genomgången farmaceutexamen).
j) I Storbritannien:
Intyg som Registered Pharmaceutical Chemist.
Artikel 5
Om det i en medlemsstat inte bara krävs ett utbildnings-, examens- eller annat behörighetsbevis för att påbörja eller utöva någon form av verksamhet som avses i artikel 1 utan även kompletterande yrkeserfarenhet, skall det landet som tillräckligt bevis godta ett intyg utfärdat av de behöriga myndigheterna i ursprungslandet eller det senaste hemvistlandet som visar att personen i fråga har utövat nämnda former av verksamhet under motsvarande period i ursprungslandet eller det senaste hemvistlandet.
Detta godkännande skall emellertid inte tillämpas på den tvååriga yrkeserfarenhet som krävs i Luxemburg för att tilldelas ett statligt tillstånd att driva ett apotek som är öppet för allmänheten.
Artikel 6
De utbildnings-, examens- och andra behörighetsbevis i farmaci som medlemsstaterna utfärdat till medborgare i medlemsstaterna och som inte uppfyller de minimivillkor för utbildningen som fastställts i artikel 2 i direktiv 85/432/EEG skall jämställas med de examensbevis som uppfyller dessa krav,
och i båda fallen,
- om de åtföljs av ett intyg som visar att innehavarna av dessa examensbevis i en medlemsstat faktiskt på föreskrivet sätt har utövat någon av de former av verksamhet som avses i artikel 1.2 i direktiv 85/432/EEG i minst tre år i följd under en femårsperiod före dagen för utfärdandet av intyget, förutsatt att det landet utfärdat bestämmelser som reglerar denna verksamhet.
KAPITEL IV Användning av akademisk titel
Artikel 7
1. Utan att det påverkar tillämpningen av artikel 14 skall värdlandet se till att medborgare i medlemsstaterna som uppfyller villkoren i artikel 2, 5 och 6 får rätt att använda den erkända akademiska titeln eller en eventuell förkortning av denna i ursprungslandet eller det senaste hemvistlandet på det landets språk. Värdlandet får kräva att denna titel åtföljs av namnet på och platsen för den institution eller examensnämnd som utfärdat den.
2. Om den akademiska titel som används i ursprungslandet eller det senaste hemvistlandet kan förväxlas med en titel som i värdlandet kräver kompletterande utbildning, som personen i fråga inte har genomgått, får värdlandet kräva att denne använder den först nämnda titeln i en lämplig form som värdlandet anger.
Artikel 8
1. Ett värdland som kräver bevis om god vandel eller bevis om gott anseende av de egna medborgare som vill påbörja sådan verksamhet som avses i artikel 1 skall när det gäller medborgare från andra medlemsstater som tillräckligt bevis godta ett intyg utfärdat av en behörig myndighet i ursprungslandet eller det senaste hemvistlandet, som visar att det landets krav på god vandel eller gott anseende för att påbörja verksamheten i fråga är uppfyllda.
2. Om det i ursprungslandet eller det senaste hemvistlandet inte krävs bevis om god vandel eller bevis om gott anseende för att påbörja verksamheten i fråga, får värdlandet kräva att personen i fråga företer utdrag ur kriminalregistret eller eventuellt motsvarande handling utfärdad av en behörig myndighet i ursprungslandet eller det senaste hemvistlandet.
4. Medlemsstaterna skall garantera de lämnade upplysningarnas konfidentiella natur.
Artikel 9
1. Om det i värdlandet finns bestämmelser i lagar och andra författningar om krav på god vandel eller gott anseende samt bestämmelser om disciplinpåföljd i händelse av allvarligt fel i yrkesutövningen eller fällande dom på grund av lagöverträdelser i samband med den yrkesutövning som avses i artikel 1, skall ursprungslandet eller det senaste hemvistlandet till värdlandet överlämna alla upplysningar som behövs om de åtgärder eller disciplinpåföljder av yrkesmässig eller administrativ karaktär som vidtagits mot personen i fråga eller om de straffrättsliga påföljder på grund av lagöverträdelser som ådömts denne under yrkesutövningen i ursprungslandet eller det senaste hemvistlandet.
2. Om värdlandet har ingående kunskap om ett allvarligt sakförhållande som har uppstått utanför dess territorium, innan personen i fråga etablerade sig i det landet, och som sannolikt kommer att påverka rätten att inom dess territorium utöva verksamheten i fråga, får det landet underrätta ursprungslandet eller det senaste hemvistlandet om detta.
Ursprungslandet eller det senaste hemvistlandet skall kontrollera riktigheten av sakförhållandena, om de sannolikt kommer att påverka rätten att i den medlemsstaten utöva verksamheten i fråga. Myndigheterna i det landet skall avgöra vilket slags utredningar som skall göras och i vilken omfattning och skall underrätta värdlandet om eventuella åtgärder som de vidtar med avseende på de upplysningar som överlämnats i enlighet med punkt 1.
3. Medlemsstaterna skall garantera de lämnade upplysningarnas konfidentiella natur. Artikel 10
Om värdlandet kräver intyg om den fysiska och psykiska hälsan av de egna medborgare som vill påbörja eller utöva sådan verksamhet som avses i artikel 1, skall det landet som tillräckligt bevis godta den handling som krävs i ursprungslandet eller det senaste hemvistlandet.
Om det i ursprungslandet eller det senaste hemvistlandet inte ställs några krav av detta slag för att påbörja eller utöva verksamheten i fråga, skall värdlandet godta intyg som utfärdats av behörig myndighet i det andra landet och som motsvarar de intyg som utfärdas i värdlandet.
Artikel 11
Handlingar som utfärdats i enlighet med artikel 8, 9 och 10 får när de företes inte vara äldre än tre månader.
Artikel 12
1. Det förfarande som genomförs enligt artikel 8, 9 och 10 för att personen i fråga skall beviljas tillstånd att utöva sådan verksamhet som avses i artikel 1 avslutas snarast möjligt och senast tre månader efter det att samtliga handlingar som rör denna person inlämnats med beaktande av de förseningar som kan uppstå på grund av eventuella överklaganden efter det att detta förfarande genomförts.
2. I de fall som avses i artikel 8.3 och 9.2 skall en begäran om utredning medföra att den tidsfrist som fastställts i punkt 1 förlängs.
Det ursprungsland eller senaste hemvistland som rådfrågats skall avge svar inom tre månader.
Efter att ha mottagit svaret eller efter tidsfristens utgång skall värdlandet fortsätta det förfarande som avses i punkt 1.
Artikel 13
Om ett värdland kräver att de egna medborgare som vill påbörja eller utöva den verksamhet som avses i artikel 1 avlägger ed eller avger en högtidlig försäkran och om formen för en sådan ed eller försäkran inte kan användas av medborgare i andra medlemsstater, skall värdlandet se till att en lämplig och likvärdig form av ed eller försäkran erbjuds personen i fråga.
Artikel 14
Om användningen av yrkestiteln för sådan verksamhet som avses i artikel 1 är reglerad i ett värdland, skall medborgare från andra medlemsstater som uppfyller villkoren i artikel 2, 5 och 6 använda den titel i värdlandet, som i det landet motsvarar denna utbildningsnivå, även i titelns förkortade form.
Artikel 15
1. Medlemsstaterna skall vidta nödvändiga åtgärder för att göra det möjligt för personerna i fråga att erhålla upplysningar om hälso- och socialförsäkringslagstiftningen och, där så är tillämpligt, om de yrkesetiska reglerna i värdlandet.
För detta ändamål får medlemsstaterna upprätta informationskontor där dessa personer kan få de upplysningar som behövs. Vid etablering får värdlandet kräva att personerna i fråga kontaktar dessa kontor.
2. Medlemsstaterna får upprätta de kontor som avses i punkt 1 vid de behöriga myndigheterna och organen, som de måste utse inom den tidsfrist som fastställts i artikel 19.1.
3. Medlemsstaterna skall se till att, där så är lämpligt, personerna i fråga i deras eget och deras patienters intresse förvärvar de språkkunskaper som krävs för att utöva yrket i värdlandet.
Artikel 16
Om det finns skälig grund till tvivel får värdlandet kräva att de behöriga myndigheterna i en annan medlemsstat styrker äktheten av utbildnings-, examens- och andra behörighetsbevis som utfärdats i den andra medlemsstaten och som avses i kapitel II och III samt styrker att personen i fråga har uppfyllt utbildningsvillkoren i direktiv 85/432/EEG.
Artikel 17
Inom den tidsfrist som fastställts i artikel 19.1 skall medlemsstaterna utse de myndigheter och organ som är behöriga att utfärda eller motta utbildnings-, examens- och andra behörighetsbevis samt de handlingar och upplysningar som avses i detta direktiv. De skall genast underrätta övriga medlemsstater och kommissionen om detta.
Artikel 18
Detta direktiv skall även tillämpas på de medborgare i medlemsstaterna som i enlighet med förordning (EEG) nr 1612/68 i egenskap av anställda utövar eller kommer att utöva sådan verksamhet som avses i artikel 1. Artikel 19
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta direktiv före den 1 oktober 1987. De skall genast underrätta kommissionen om detta.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 20
Om det vid tillämpningen av detta direktiv skulle uppstå allvarligare svårigheter för en medlemsstat inom vissa områden, skall kommissionen i samverkan med det landet undersöka dessa svårigheter och begära yttrande från den farmaceutiska nämnd som upprättats enligt beslut 75/320/EEG().
I mån av behov skall kommissionen föreslå rådet lämpliga åtgärder.
Artikel 21
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 20 december 1985 om samordning av lagar och andra författningar som avser företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag) (85/611/EEG)
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
med beaktande av följande:Medlemsstaternas författningsregler beträffande företag för kollektiva investeringar varierar avsevärt, särskilt i fråga om de skyldigheter och den övervakning som gäller för sådana företag. Dessa olikheter inverkar negativt på villkoren för konkurrens mellan företagen och ger inte likvärdigt skydd för andelsägarna.
Med hänsyn till dessa målsättningar bör gemensamma grundregler införas om auktorisation, tillsyn, organisation och verksamheter för medlemsstaternas företag för kollektiva investeringar hemmahörande i medlemsstaterna och för den information de skall offentliggöra.
Sådana gemensamma regler ger en tillräcklig garanti för att medlemsstaternas företag för kollektiva investeringar, med iakttagande av vad som skall gälla beträffande kapitalrörelser, skall kunna utbjuda sina andelar i andra medlemsstater utan att dessa skall ha möjlighet att för företagen eller deras andelar tillämpa några andra bestämmelser än sådana som faller utanför direktivets tillämpningsområde. Ett företag för kollektiva investeringar som utbjuder sina andelar i en annan medlemsstat än där företaget hör hemma, skall dock vidta alla åtgärder som krävs för att andelsägarna där skall kunna utöva sina finansiella rättigheter utan svårighet och få tillgång till nödvändig information.
Samordningen av medlemsstaternas lagstiftning skall till en början begränsas till att avse företag för kollektiva investeringar av icke sluten typ som utbjuder sina andelar till allmänheten inom gemenskapen och som har som enda syfte att investera i överlåtbara värdepapper (dvs. väsentligen överlåtbara värdepapper som är officiellt noterade vid fondbörser eller liknande reglerade marknadsplatser). Regleringen av företag för kollektiva investeringar som inte omfattas av direktivet erbjuder en mängd problem som måste lösas med hjälp av andra bestämmelser, och sådana företag kommer följaktligen att bli föremål för samordning i ett senare skede. I avvaktan på sådan samordning får varje enskild medlemsstat bl.a. från direktivets tillämpningsområde undanta kategorier av företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag) som har speciell placerings- och upplåningsinriktning och uppställa särskilda regler för dessa företags verksamhet inom den medlemsstaten.
Den fria marknadsföringen av andelar som utgivits av fondföretag som fått tillstånd att placera upp till 100% av sina tillgångar i överlåtbara värdepapper från samma emittent (stat, lokal myndighet, etc.) får varken direkt eller indirekt åstadkomma störningar i kapitalmarknadens funktion eller medlemsstaternas finansiering eller skapa ekonomiska situationer av det slag som artikel 68.3 i fördraget avser att förhindra.
Hänsyn bör tas till de särskilda omständigheter som råder beträffande de finansiella marknaderna i Grekland och Portugal genom att dessa länder medges en förlängd frist för att genomföra detta direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
AVSNITT I Allmänna bestämmelser och räckvidd
3. Sådana företag kan bildas med stöd av lag, antingen på kontraktsrättslig grund (som värdepappersfonder förvaltade av förvaltningsföretag) eller enligt trustlagstiftning (som "unit trusts") eller på bolagsrättslig grund (som investeringsbolag).
Vid tillämpningen av detta direktiv skall med värdepappersfonder avses även "unit trusts".
4. Detta direktiv skall emellertid inte tillämpas på investeringsbolag vars tillgångar via dotterbolag är placerade huvudsakligen i annat än överlåtbara värdepapper.
5. Medlemsstaterna skall förbjuda fondföretag för vilka detta direktiv gäller att ombilda sig till sådant företag för kollektiva investeringar som inte omfattas av direktivets bestämmelser.
6. Med förbehåll för bestämmelserna om kapitalrörelser och bestämmelserna i artiklarna 44, 45 och 52.2 får en medlemsstat, i de avseenden som regleras i detta direktiv, inte tillämpa andra bestämmelser för fondföretag hemmahörande i en annan medlemsstat, eller för andelar som utgivits av sådana företag, i de fall de utbjuder sina andelar inom medlemsstatens territorium.
7. Bestämmelserna i punkt 6 hindrar inte en medlemsstat att på fondföretag hemmahörande i den egna staten ställa krav som är strängare eller som går utöver vad som föreskrivs i artikel 4 och följande artiklar, förutsatt att kraven är generellt tillämpbara och inte står i strid med bestämmelserna i detta direktiv.
Artikel 2
- Fondföretag vars andelar enligt fondbestämmelserna eller bolagsordningen får säljas endast till allmänheten i icke-medlemsländer.
- Kategorier av fondföretag enligt vad som föreskrivs av medlemsstater där företagen hör hemma och för vilka bestämmelserna i avsnitt V och artikel 36 inte är ändamålsenliga med hänsyn till den placerings- och upplåningsinriktning som företagen har.
2. Senast fem år efter genomförandet av detta direktiv skall kommissionen överlämna en rapport till rådet över tillämpningen av bestämmelserna i punkt 1, särskilt dess fjärde strecksats. Om så erfordras skall kommissionen föreslå lämpliga åtgärder för att utöka bestämmelsernas tillämpningsområde.
Artikel 3
Vid tillämpningen av detta direktiv skall ett fondföretag anses hemmahörande i den medlemsstat där investeringsbolaget eller förvaltningsbolaget har sitt stadgeenliga säte; medlemsstaterna skall föreskriva att företagets huvudkontor skall vara beläget i samma medlemsstat som dess stadgeenliga säte.
AVSNITT II Auktorisation av fondföretag
Artikel 4
1. Inget fondföretag får bedriva verksamhet utan auktorisation av behöriga myndigheter i den medlemsstat där företaget hör hemma (i fortsättningen kallade "behöriga myndigheter").
Auktorisationen skall gälla i samtliga medlemsstater.
2. En värdepappersfond får auktoriseras endast om de behöriga myndigheterna godkänt förvaltningsbolaget, fondbestämmelserna och valet av förvaringsinstitut. Ett investeringsbolag får auktoriseras endast om de behöriga myndigheterna godkänt både dess bolagsordning och valet av förvaringsinstitut.
3. De behöriga myndigheterna får inte auktorisera ett fondföretag, om de som ingår i den verkställande ledningen för förvaltningsbolaget, investeringsbolaget eller förvaringsinstitutet inte har erforderlig vandel eller om de saknar tillräcklig erfarenhet för att kunna utföra sina uppgifter. För detta ändamål skall de behöriga myndigheterna utan dröjsmål underrättas om namnen på personer i sådan ledande ställning samt namnen på var och en som efterträder dem.
Med den verkställande ledningen avses de personer som, i enlighet med lag eller annan författning eller bolagsordning, företräder förvaltningsbolaget, investeringsbolaget eller förvaringsinstitutet eller som faktiskt bestämmer verksamhetsinriktningen för sådana företag.
4. Utan de behöriga myndigheternas godkännande får varken förvaltningsbolaget eller förvaringsinstitutet bytas ut, eller fondbestämmelserna eller investeringsbolagets bolagsordning ändras.
AVSNITT III Bestämmelser om värdepappersfonders organisation
Artikel 5
Ett förvaltningsbolag skall ha finansiella resurser som är tillräckliga för att bolaget skall kunna bedriva sin verksamhet på ett effektivt sätt och uppfylla sina förpliktelser.
Artikel 6
Ett förvaltningsbolag får inte ägna sig åt annan verksamhet än förvaltning av värdepappersfonder och investeringsbolag.
Artikel 7
1. Tillgångarna i en värdepappersfond skall förvaras hos ett förvaringsinstitut.
2. Ett förvaringsinstituts ansvarighet enligt artikel 9 skall gälla oberoende av om institutet anförtrott förvaringen av samtliga eller vissa tillgångar till någon annan.
d) tillse att ersättningar för transaktioner som berör en värdepappersfonds tillgångar inbetalas till institutet inom sedvanlig tid,
e) tillse att en värdepappersfonds intäkter används i enlighet med lag eller annan författning och med fondbestämmelserna.
Artikel 8
1. Ett förvaringsinstitut skall antingen ha sitt stadgeenliga säte i samma medlemsstat som förvaltningsbolaget eller vara etablerat där om det har sitt stadgeenliga säte i en annan medlemsstat.
2. Ett förvaringsinstitut skall stå under offentlig tillsyn. Det skall också kunna ställa erforderliga ekonomiska garantier samt besitta tillfredsställande sakkunskap och kompetens för att kunna effektivt bedriva verksamhet som förvaringsinstitut och uppfylla därmed förenade åtaganden.
3. Medlemsstaterna skall bestämma vilka av de kategorier av institut som avses i punkt 2 som skall kunna utses till förvaringsinstitut.
Artikel 9
Ett förvaringsinstitut skall i enlighet med den nationella lagstiftningen i den stat där förvaltningsbolaget har sitt stadgeenliga säte vara ansvarigt mot förvaltningsbolaget och andelsägarna för förluster som drabbar dem som följd av att institutet allvarligt försummat sina förpliktelser eller fullgjort dem på ett oriktigt sätt. Detta ansvar kan av andelsägarna åberopas antingen direkt eller indirekt genom förvaltningsbolaget, beroende på hur rättsförhållandet mellan förvaringsinstitutet, förvaltningsbolaget och andelsägarna är utformat.
Artikel 10
1. Ett företag får inte samtidigt vara förvaltningsbolag och förvaringsinstitut.
2. Förvaltningsbolaget och förvaringsinstitutet skall utföra sina respektive uppgifter självständigt och uteslutande i andelsägarnas intresse.
Artikel 11
Villkoren för utbyte av förvaltningsbolaget eller förvaringsinstitutet skall, liksom regler till skydd för andelsägare vid sådana utbyten, föreskrivas i lag eller annan författning eller anges i fondbestämmelserna.
AVSNITT IV Bestämmelser om investeringsbolags organisation och och om deras förvaringsinstitut
Artikel 12
Medlemsstaterna skall bestämma vilken rättslig form ett investeringsbolag skall ha. Ett investeringsbolag skall ha ett så stort inbetalt kapital att det kan bedriva verksamheten effektivt och uppfylla sina förpliktelser.
Artikel 13
Ett investeringsbolag får inte bedriva andra verksamheter än de som anges i artikel 1.2.
Artikel 14
1. Ett investeringsbolags tillgångar skall förvaras hos ett förvaringsinstitut.
2. Ett förvaringsinstituts ansvarighet enligt artikel 16 skall gälla oberoende av om institutet anförtrott förvaringen av samtliga eller vissa tillgångar till någon annan.
3. Ett förvaringsinstitut skall vidare
a) tillse att försäljning, utgivning, återköp, inlösen och makulering av andelar, som sker av eller på uppdrag av ett investeringsbolag, genomförs i enlighet med lag eller annan författning och med bolagsordningen,
c) tillse att ett bolags intäkter används i enlighet med lag eller annan författning och med bolagsordningen.
4. En medlemsstat får besluta att investeringsbolag som hör hemma i den staten och som utbjuder sina andelar uteslutande på en eller flera fondbörser där andelarna är officiellt noterade, inte skall vara skyldiga att anlita förvaringsinstitut som avses i detta direktiv.
Artiklarna 34, 37 och 38 skall inte gälla sådana bolag som nu sagts. Bestämmelserna om värdering av sådana bolags tillgångar måste emellertid vara angivna i lag eller annan författning eller i bolagsordningen.
5. En medlemsstat får bestämma att investeringsbolag som hör hemma i den staten och som utbjuder minst 80% av sina andelar på en eller flera fondbörser, vilka finns angivna i deras bolagsordningar, inte skall vara skyldiga att ha förvaringsinstitut som avses i detta direktiv, förutsatt att deras andelar noteras officiellt på fondbörserna i de medlemsstater där andelarna utbjuds, och att varje transaktion som ett sådant investeringsbolag kan komma att göra utanför fondbörserna sker uteslutande till börskurs. I ett investeringsbolags bolagsordning skall anges en fondbörs i varje land där andelar utbjuds och vars kursnotering skall vara bestämmande för de priser som skall gälla vid transaktioner som bolaget genomför utanför fondbörser i det landet.
En medlemsstat får utnyttja den möjlighet som ges i föregående stycke endast om den finner att andelsägarna har ett skydd som är likvärdigt med det som tillkommer andelsägare i fondföretag med förvaringsinstitut som avses i detta direktiv.
b) agera (intervenera) på marknaden för att hindra att marknadsvärdet för andelarna avviker mer än 5% från nettovärdet,
c) fastställa andelarnas nettovärde, lämna uppgift om nettovärdet till de behöriga myndigheterna minst två gånger per vecka och offentliggöra uppgifter om nettovärdet två gånger per månad.
Minst två gånger per månad skall en oberoende revisor kontrollera att andelarnas värde beräknas i enlighet med lag eller annan författning och med bolagsordningen. Vid sådana tillfällen skall revisorn kontrollera att bolagets tillgångar är placerade i enlighet med lag eller annan författning och med bolagsordningen.
6. Medlemsstaterna skall underrätta kommissionen om de investeringsbolag för vilka säregler, medgivna enligt punkterna 4 och 5, tillämpas.
Kommissionen skall senast inom fem år från det att detta direktiv genomförts underrätta kontaktkommittén om tillämpningen av bestämmelserna i punkterna 4 och 5. När kontaktkommitténs yttrande erhållits skall kommissionen, om det behövs, föreslå lämpliga åtgärder.
Artikel 15
1. Ett förvaringsinstitut skall antingen ha sitt stadgeenliga säte i samma medlemsstat som investeringsbolaget eller vara etablerat där om det har sitt stadgeenliga säte i en annan medlemsstat.
2. Ett förvaringsinstitut skall stå under offentlig tillsyn. Det skall också kunna ställa erforderliga ekonomiska garantier samt besitta tillfredsställande sakkunskap och kompetens för att kunna effektivt bedriva verksamhet som förvaringsinstitut och uppfylla därmed förenade åtaganden.
3. Medlemsstaterna skall bestämma vilka av de kategorier av institut som avses i punkt 2 som skall kunna utses till förvaringsinstitut.
Artikel 16
Ett förvaringsinstitut skall i enlighet med den nationella lagstiftningen i den stat där investeringsbolaget har sitt stadgeenliga säte vara ansvarigt mot investeringsbolaget och andelsägarna för förluster som drabbar dem som följd av att institutet allvarligt försummat sina förpliktelser eller fullgjort dem på ett oriktigt sätt.
Artikel 17
1. Ett företag får inte samtidigt vara investeringsbolag och förvaringsinstitut.
2. Ett förvaringsinstitut skall vid utförande av sina uppgifter handla uteslutande i andelsägarnas intresse.
Artikel 18
Villkoren för utbyte av förvaringsinstitut skall, liksom regler till skydd för andelsägarna vid sådana utbyten, föreskrivas i lag eller annan författning eller anges i investeringsbolagets bolagsordning.
AVSNITT V Placeringsbestämmelser för fondföretag
Artikel 19
b) överlåtbara värdepapper som är föremål för handel på någon annan reglerad marknad i en medlemsstat och vilken marknadsplats fungerar fortlöpande och är erkänd och öppen för allmänheten, och/eller
c) överlåtbara värdepapper som är officiellt noterade på en fondbörs i en icke-medlemsstat eller som är föremål för handel på någon annan reglerad marknadsplats i en icke-medlemsstat och vilken marknadsplats fungerar fortlöpande och är erkänd och öppen för allmänheten, förutsatt att valet av fondbörs eller annan marknadsplats godkänts av de behöriga myndigheterna eller är reglerat i lag eller annan författning eller i fondbestämmelserna eller i investeringsbolagets bolagsordning, och/eller
a) ett fondföretag får placera högst 10% av sina fondtillgångar i andra överlåtbara värdepapper än de som avses i punkt 1,
b) en medlemsstat får föreskriva att ett fondföretag får placera högst 10% av sina tillgångar i fordringsbevis som med hänsyn till sin natur kan jämställas med överlåtbara värdepapper och för vilka bland annat gäller att de är överlåtbara och likvida och vars värde kan nöjaktigt bestämmas när som helst eller i vart fall så ofta som sägs i artikel 34,
c) ett investeringsbolag får förvärva lös och fast egendom som det behöver för sin verksamhet,
d) ett fondföretag inte får förvärva ädla metaller eller värdepapper inlösbara i sådana metaller.
3. Summan av placeringar som nämns i punkt 2 a och b får aldrig motsvara mer än 10% av ett fondföretags tillgångar.
4. Värdepappersfonder och investeringsbolag får ha kompletterande likvida tillgångar.
Artikel 20
b) närmare upplysningar om alla ändringar de avser att göra i förteckningar enligt a eller om andra instrument som de avser att jämställa med överlåtbara värdepapper, med angivande av skälen.
1. Medlemsstaterna får ge fondföretag tillstånd att använda sig av sådan teknik och sådana instrument som hänför sig till överlåtbara värdepapper under de villkor och inom de ramar staterna föreskriver, förutsatt att sådan teknik och sådana instrument används i syfte att åstadkomma en effektiv förvaltning av värdepappersportföljen.
2. Medlemsstaterna får också ge fondföretag tillstånd att vid förvaltningen av sina tillgångar och skulder utnyttja sådan teknik och sådana instrument som syftar till att ge skydd mot valutarisker.
Artikel 22
1. Ett fondföretag får placera högst 5% av fondtillgångarna i överlåtbara värdepapper med samme utgivare.
2. Medlemsstaterna får höja den gräns som anges i punkt 1 till högst 10%. I den mån fondföretaget placerar mer än 5% av fondtillgångarna i överlåtbara värdepapper med samme utgivare, får det sammanlagda innehavet av sådana placeringar inte överstiga 40% av fondtillgångarna.
3. Medlemsstaterna får höja den gräns som anges i punkt 1 till högst 35% om de överlåtbara värdepapperen är utgivna eller garanterade av en medlemsstat, av dess lokala myndigheter, av en icke-medlemsstat eller av offentliga internationella organ i vilka en eller flera medlemsstater är medlemmar.
Artikel 23
1. Utan hinder av artikel 22, med förbehåll för artikel 68.3 i fördraget, får medlemsstaterna ge fondföretag tillstånd att med tillämpning av principen om riskspridning placera upp till 100% av fondtillgångarna i olika överlåtbara värdepapper utgivna eller garanterade av en medlemsstat, dess lokala myndigheter, en icke-medlemsstat eller offentliga internationella organ i vilka en eller flera medlemsstater är medlemmar.
De behöriga myndigheterna får medge sådana undantag endast om de finner att andelsägarna i fondföretaget har ett skydd likvärdigt med det som tillkommer andelsägarna i fondföretag som iakttar de gränsvärden som anges i artikel 22.
Ett sådant fondföretag skall inneha värdepapper från minst sex olika emissioner, varvid dock skall gälla att värdepapper från en och samma emission inte får motsvara mer än 30% av de samlade fondtillgångarna.
2. Fondbestämmelserna eller bolagsordningarna för de fondföretag som avses i punkt 1 skall innehålla uttrycklig uppgift om de stater, lokala myndigheter och offentliga internationella organ som utger eller garanterar sådana värdepapper i vilka fondföretaget avser att placera mer än 35% av fondtillgångarna; sådana fondbestämmelser och bolagsordningar måste godkännas av behöriga myndigheter.
3. De fondföretag som avses i punkt 1 skall vidare i sina prospekt och reklambroschyrer på framträdande plats omnämna tillståndet och ange de stater, lokala myndigheter och/eller offentliga internationella organ i vars värdepapper de har för avsikt att placera eller har placerat mer än 35% av fondtillgångarna.
Artikel 24
1. Ett fondföretag får inte förvärva fondandelar i andra företag för kollektiva investeringar av den öppna typen, såvida dessa inte är företag för kollektiva investeringar i den betydelse som avses i första och andra strecksatserna i artikel 1.2.
2. Ett fondföretag får placera högst 5% av sina tillgångar i andelar i sådana företag för kollektiva investeringar.
3. Placeringar i andelar i en värdepappersfond som förvaltas av samma förvaltningsbolag eller av ett annat företag med vilket förvaltningsbolaget är anknutet via gemensam företagsledning eller ägarkontroll eller genom ett betydande direkt eller indirekt ägande får tillåtas endast om det rör sig om en fond som, i enlighet med sina fondbestämmelser, har specialiserat sig på placeringar inom ett visst geografiskt område eller en viss ekonomisk sektor och förutsatt att sådana placeringar medges av de behöriga myndigheterna. Tillstånd skall ges endast om fonden har meddelat sin avsikt att utnyttja denna möjlighet och möjligheten uttryckligen angivits i dess fondbestämmelser.
Ett förvaltningsbolag får inte debitera några avgifter eller kostnader för transaktioner som hänför sig till en viss värdepappersfonds andelar i fall där några av en värdepappersfonds tillgångar är placerade i andelarna i en annan värdepappersfond som förvaltas av samma förvaltningsbolag eller av ett annat bolag med vilket förvaltningsbolaget är anknutet via gemensam företagsledning eller ägarkontroll eller genom ett betydande direkt eller indirekt ägande.
4. Punkt 3 skall även gälla i fall där ett investeringsbolag förvärvar fondandelar i ett annat investeringsbolag till vilket det är anknutet på det sätt som anges i punkt 3.
1. Ett investeringsbolag eller ett förvaltningsbolag får, såvitt gäller handhavandet av alla de värdepappersfonder som står under bolagets förvaltning och som omfattas av bestämmelserna i detta direktiv, inte förvärva aktier med sådan rösträtt som skulle göra det möjligt för bolaget att utöva ett väsentligt inflytande över ledningen hos en emittent.
I avvaktan på vidare samordning skall medlemsstaterna beakta gällande föreskrifter i andra medlemsstaters lagstiftning, som närmare uttrycker den i föregående stycke angivna principen.
- 10% av de skuldebrev som en enskild emittent givit ut,
- 10% av andelarna i ett sådant företag för kollektiva investeringar som avses i första och andra strecksatserna i artikel 1.2.
De gränsvärden som anges i andra och tredje strecksatserna behöver inte iakttas vid förvärvstillfället, om bruttomängden av skuldebreven eller nettomängden av de värdepapper som är under utgivning då inte kan uppskattas.
d) Ett fondföretags innehav av aktier i ett bolag beläget i en icke-medlemsstat och vars tillgångar placeras huvudsakligen i värdepapper utgivna av emittenter med sitt stadgeenliga säte i den staten, då den statens lagstiftning inte gör det möjligt för fondföretaget att på något annat sätt placera sina fondtillgångar i värdepapper med utgivare i staten. Detta undantag gäller dock endast om bolaget från icke-medlemsstaten vid sina placeringar följer de gränsvärden som anges i artiklarna 22, 24 och 25.1 och 25.2. Om gränsvärdena i artikel 22 och 24 har överskridits skall artikel 26 gälla i tillämpliga delar.
e) Ett investeringsbolags aktieinnehav i dotterbolag vars verksamhet består i förvaltning, rådgivning eller avsättning uteslutande för investeringsbolagets räkning.
Artikel 26
1. Fondföretag behöver inte iaktta de gränsvärden som anges i detta avsnitt när de utnyttjar teckningsrätter för överlåtbara värdepapper som ingår i fondtillgångarna.
Medlemsstaterna får, med beaktande av principen om riskspridning, tillåta nyligen auktoriserade fondföretag att under en tid av högst sex månader från auktorisationsdagen avvika från vad som föreskrivits i artiklarna 22 och 23.
2. Om gränsvärdena enligt punkt 1 överskrids av skäl som ligger utanför ett fondföretags rådighet eller som följd av att teckningsrätter utnyttjas, skall fondföretaget vid sina försäljningstransaktioner prioritera rättelse av detta förhållande under vederbörligt hänsynstagande till andelsägarnas intressen. AVSNITT VI
Bestämmelser om information till andelsägarna A. Offentliggörande av prospekt och periodiska rapporter
Artikel 27
1. Ett investeringsbolag och ett förvaltningsbolag, det senare för varje värdepappersfond det förvaltar, skall offentliggöra
- Två månader för halvårsrapporter.
Artikel 28
1. Ett prospekt skall innehålla den information som krävs för att investerare skall kunna göra en välgrundad bedömning av den erbjudna investeringen. Prospektet skall innehålla minst den information som anges i lista A i bilagan till detta direktiv, såvida inte informationen redan framgår av de handlingar som skall bifogas prospektet enligt artikel 29.1.
2. Årsrapporten skall innehålla en balansräkning eller en redovisning av tillgångar och skulder, en specificerad resultaträkning för räkenskapsåret, en verksamhetsberättelse för räkenskapsåret samt den information som anges i lista B i bilagan till detta direktiv, liksom all annan väsentlig information som möjliggör för investerare att göra en välgrundad bedömning av utvecklingen av fondföretagets verksamhet och av dess resultat.
3. Halvårsrapporten skall innehålla minst den information som anges i kapitel I-IV i lista B i bilagan till detta direktiv; om ett fondföretag har utbetalat eller föreslår utbetalning av interimsutdelning, skall i redovisningen anges resultatet efter skatt för halvårsperioden i fråga samt den interimsutdelning som utbetalats eller föreslås.
Artikel 29
1. Fondbestämmelserna eller investeringsbolagets bolagsordning skall utgöra en del av prospektet och skall bifogas till detta.
2. De handlingar som avses i punkt 1 behöver dock inte bifogas prospektet om andelsägarna informerats om att de på begäran kommer att tillställas dessa handlingar eller få upplysning om var i varje medlemsstat, där andelarna finns på marknaden, de kan ta del av handlingarna.
Artikel 30
All väsentlig information i ett prospekt måste hållas aktuell.
Artikel 31
De uppgifter om räkenskaperna som årsrapporten innehåller skall vara granskade av en eller flera personer som enligt lag eller annan författning bemyndigats att granska redovisningar i överensstämmelse med rådets direktiv 84/253/EEG av den 10 april 1984 grundat på artikel 54.3 g i Romfördraget, om godkännande av personer som har ansvar för lagstadgad revision av räkenskaper (4). Revisionsberättelsen, med eventuella anmärkningar, skall i sin helhet återges i årsrapporten.
Artikel 32
Ett fondföretag skall till de behöriga myndigheterna ge in sina prospekt och eventuella ändringar och tillägg i dessa, liksom årsrapporter och halvårsrapporter.
Artikel 33
1. Den som avser att teckna sig för förvärv av fondandelar skall innan avtalet ingås erbjudas att kostnadsfritt få prospektet, den senaste halvårsrapporten samt, i förekommande fall, den därpå följande halvårsrapporten.
2. Årsrapporterna och halvårsrapporterna skall finnas tillgängliga för allmänheten på i prospektet angivna platser.
3. Årsrapporterna och halvårsrapporterna skall på begäran kostnadsfritt tillställas andelsägarna.
B. Offentliggörande av annan information
Artikel 34
Ett fondföretag skall vid varje tillfälle då det emitterar, säljer, återköper eller löser in andelar, dock minst två gånger per månad, på lämpligt sätt offentliggöra emissions-, försäljnings-, återköps- och inlösenpriserna. De behöriga myndigheterna får dock medge ett fondföretag att offentliggöra sådana uppgifter endast en gång per månad, förutsatt att andelsägarnas intressen inte härigenom åsidosätts.
Artikel 35
Vid all marknadsföring av ett fondföretags andelar skall anges att ett prospekt finns och uppges var allmänheten kan få tillgång till prospektet. AVSNITT VII
Fondföretags allmänna förpliktelser
Artikel 36
2. Trots bestämmelserna i punkt 1 får en medlemsstat ge fondföretag tillstånd att låna
a) upp till 10% - av tillgångarna, i fråga om ett investeringsbolag eller,
- av fondens värde, i fråga om en värdepappersfond, förutsatt att upplåningen är av tillfällig art,
b) upp till 10% av tillgångarna, i fråga om ett investeringsbolag, förutsatt att upplåningen har till syfte att möjliggöra förvärv av fast egendom som det behöver för verksamheten; i detta fall får summan av denna upplåning och den som avses i a inte överstiga 15% av låntagarens tillgångar.
Artikel 37
1. Ett fondföretag skall återköpa eller inlösa andelar när andelsägare begär det.
b) Medlemsstaterna får tillåta de behöriga myndigheterna att kräva att återköp eller inlösen av andelar senareläggs med hänsyn till andelsägarnas eller allmänhetens intresse.
3. I de fall som avses i punkt 2 a, skall ett fondföretag utan dröjsmål underrätta de berörda myndigheterna och myndigheterna i samtliga medlemsstater där företaget utbjuder sina andelar om uppskovsbeslutet.
Artikel 38
Reglerna för värdering av tillgångar och för beräkning av försäljnings- eller emissionspris samt återköps- eller inlösenpris på ett fondföretags andelar skall vara föreskrivna i lag eller annan författning, i fondbestämmelserna eller i investeringsbolagets bolagsordning.
Artikel 39
Utdelningen eller återinvestering av en värdepappersfonds eller ett investeringsbolags intäkter skall ske i enlighet med lag eller annan författning och fondbestämmelserna eller investeringsbolagets bolagsordning.
Artikel 40
Ett fondföretags andelar får emitteras endast om fondtillgångarna inom sedvanlig tid tillförs betalning motsvarande emissionens nettopris. Denna bestämmelse skall inte utgöra hinder för tilldelning av bonusandelar.
Artikel 41
1. Med undantag för sådana fall som avses i artiklarna 19 och 21 gäller att varken
- ett förvaltningsbolag eller förvaringsinstitut som handlar för en värdepappersfonds räkning får bevilja lån eller ingå borgen för någon annans räkning.
2. Bestämmelserna i punkt 1 skall inte hindra sådana företag från att förvärva överlåtbara värdepapper som inte är till fullo betalda.
Artikel 42
Artikel 43
I lag eller annan författning eller i fondbestämmelserna skall det anges vilken ersättning och vilka kostnader ett förvaltningsbolag har rätt att debitera en värdepappersfond och vilken metod som skall tillämpas för beräkning av sådana vederlag.
I lag eller annan författning eller i ett investeringsbolags bolagsordning skall det anges vilka kostnader som skall bäras av bolaget.
AVSNITT VIII Särskilda bestämmelser för fondföretag som utbjuder sina andelar i andra medlemsstater än dem där företagen är hemmahörande
Artikel 44
1. Ett fondföretag som utbjuder sina andelar i en annan medlemsstat måste följa de lagar och andra författningar som gäller i den staten, och som inte faller inom tillämpningsområdet för detta direktiv.
2. Ett fondföretag får marknadsföra sina andelar i de medlemsstater där dessa utbjuds. Det måste därvid följa de bestämmelser om reklam som gäller i det landet.
3. Bestämmelserna i punkterna 1 och 2 får inte tillämpas på ett diskriminerande sätt.
Artikel 45
I det fall som avses i artikel 44 skall fondföretagen, i enlighet med de lagar och andra författningar som gäller i den medlemsstat där andelarna utbjuds, bl.a. vidta erforderliga åtgärder för att där kunna göra utbetalningar till andelsägarna, verkställa återköp och inlösen samt lämna ut den information som fondföretagen är skyldiga att tillhandahålla.
Artikel 46
- sina fondbestämmelser eller sin bolagsordning,
- sitt prospekt,
- där det anses lämpligt, sin senaste årsrapport och eventuell senare halvårsrapport, samt - upplysningar om de åtgärder som vidtagits för försäljning av dess andelar i den andra medlemsstaten.
Om ett fondföretag utbjuder sina andelar i en annan medlemsstat än den där företaget är beläget, skall det i den andra medlemsstaten, på minst ett av den andra medlemsstatens officiella språk, tillhandahålla de handlingar och den information som skall offentliggöras i den medlemsstat där det är hemmahörande, i den ordning som föreskrivs i den sistnämnda staten.
Artikel 48
Ett fondföretag skall i sin verksamhet ha rätt att använda samma företagsbeteckning (t.ex. investeringsbolag eller värdepappersfond) inom hela gemenskapen som det använder i den medlemsstat där det är hemmahörande. Om det finns risk för förväxling kan värdmedlemsstaten i förtydligande syfte begära att namnet skall åtföljas av något förklarande tillägg.
AVSNITT IX Bestämmelser om de myndigheter som svarar för auktorisation och tillsyn
Artikel 49
1. Medlemsstaterna skall utse de myndigheter som skall fullgöra de uppgifter som föreskrivs i detta direktiv. Medlemsstaterna skall underrätta kommissionen om detta och i förekommande fall ange hur uppgifterna fördelats mellan myndigheterna.
2. De myndigheter som avses i punkt 1 skall vara offentliga myndigheter eller institutioner utsedda av offentliga myndigheter.
3. Myndigheterna i den stat där ett fondföretag är hemmahörande skall vara behöriga att utöva tillsyn över företaget. Myndigheterna i den stat där ett fondföretag utbjuder sina andelar i enlighet med artikel 44 skall dock vara behöriga att kontrollera att bestämmelserna i avsnitt VIII följs.
4. De berörda myndigheterna skall ges alla de befogenheter som de behöver för att utföra sina uppgifter.
Artikel 50
1. De medlemsstaters myndigheter som avses i artikel 49 skall fullgöra sina uppgifter i nära samarbete och utbyta nödvändig information.
2. Medlemsstaterna skall föreskriva att alla som är eller har varit anställda hos de myndigheter som avses i artikel 49 skall vara bundna av tystnadsplikt. Detta innebär att ingen konfidentiell information som erhållits i tjänsten får röjas för någon person eller myndighet annat än med stöd av bestämmelser i lag eller annan författning.
3. Bestämmelserna i punkt 2 skall emellertid inte utesluta utbyte av information mellan de i artikel 49 angivna myndigheterna i olika medlemsstater i enlighet med bestämmelserna i detta direktiv. Beträffande sålunda utväxlad information skall anställda eller tidigare anställda hos myndigheter som erhåller information enligt ovan iaktta tystnadsplikt.
4. Utöver vad som följer av straffrättsliga föreskrifter får en myndighet som avses i artikel 49 och som erhåller ifrågavarande information använda denna endast för fullgörande av sina uppgifter samt vid överklaganden i administrativ ordning och vid rättsliga förfaranden som har samband med myndighetens verksamhet.
Artikel 51
1. Myndigheter som avses i artikel 49 skall uppge skälen för såväl beslut att vägra auktorisation som de övriga beslut med negativ innebörd som fattas i samband med införande av föreskrifter för tillämpning av detta direktiv, samt underrätta sökandena om skälen.
2. Medlemsstaterna skall sörja för att beslut som fattas med avseende på fondföretag med stöd av lag eller annan författning i enlighet med detta direktiv kan prövas av domstol. En möjlighet till domstolsprövning skall finnas också för fall då beslut inte fattats inom sex månader från det att ett fondföretag lämnat in auktorisationsansökan som innehåller all den information som krävs enligt gällande föreskrifter.
Artikel 52
1. Endast myndigheterna i den medlemsstat där ett fondföretag är beläget skall ha behörighet att vidta åtgärder mot företaget om det bryter mot lag eller annan författning eller fondbestämmelserna eller investeringsbolagets bolagsordning.
2. Myndigheterna i den medlemsstat där ett fondföretags andelar utbjuds får dock vidta åtgärder mot företaget, om det bryter mot de i avsnitt VIII nämnda bestämmelserna.
3. Myndigheterna i den medlemsstat där ett fondföretag är beläget skall utan dröjsmål underrätta myndigheterna i de medlemsstater där företaget utbjuder sina andelar om beslut som avser återkallelse av auktorisation, andra allvarliga åtgärder som riktar sig mot företaget samt uppskov med återköp eller inlösen.
AVSNITT X Kontaktkommitté
Artikel 53
1. En kontaktkommitté, i fortsättningen kallad kommittén, skall inrättas vid sidan av kommissionen. Dess funktion skall vara
a) att, så långt det inte strider mot artiklarna 169 och 170 i fördraget, underlätta ett samordnat genomförande av detta direktiv genom regelbundna samråd om praktiska problem som kan uppkomma vid dess tillämpning och beträffande vilka en diskussion bedöms ändamålsenlig,
b) att underlätta samråd mellan medlemsstater antingen beträffande skärpta eller kompletterande krav som de har rätt att uppställa i enlighet med artikel 1.7, eller beträffande föreskrifter som de får utfärda i enlighet med artiklarna 44 och 45,
c) att, om så erfordras, föreslå kommissionen tillägg till eller ändringar i detta direktiv.
2. Det skall inte ankomma på kommittén att pröva beslut som fattats i enskilda fall av de myndigheter som avses i artikel 49.
3. Kommittén skall vara sammansatt av personer utsedda av medlemsstaterna och av representanter för kommissionen. Ordföranden skall vara en representant för kommissionen. Sekretariatstjänster skall tillhandahållas av kommissionen.
4. Kommittén skall sammankallas av dess ordförande antingen på dennes eget initiativ eller på begäran av en medlemsstats delegation. Kommittén skall självständigt fastställa sin arbetsordning.
AVSNITT XI Övergångsbestämmelser, undantag och avslutande bestämmelser
Artikel 54
Uteslutande med avseende på danska fondföretag skall "pantebreve" utställda i Danmark jämställas med de överlåtbara värdepapper som avses i artikel 19.1 b.
Artikel 55
Trots bestämmelserna i artiklarna 7.1 och 14.1 får de behöriga myndigheterna tillåta sådana fondföretag som i enlighet med nationell lagstiftning hade två eller flera förvaringsinstitut vid tidpunkten för antagandet av detta direktiv att behålla dessa institut, om myndigheterna har garantier för att de uppgifter som föreskrivs i artiklarna 7.3. och 14.3 kommer att fullgöras i praktiken.
Artikel 56
1. Trots bestämmelserna i artikel 6 får medlemsstaterna tillåta förvaltningsbolag att emittera innehavarbevis avseende andra företags registrerade värdepapper.
2. Medlemsstaterna får bevilja förvaltningsbolag som, vid tidpunkten för antagande av detta direktiv bedriver andra verksamheter än sådana som tillåts enligt artikel 6, att fortsätta med dessa i fem år efter nämnda tidpunkt.
Artikel 57
1. Medlemsstaterna skall senast den 1 oktober 1989 sätta i kraft de beslut som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
2. Medlemsstaterna får bevilja fondföretag, som var verksamma vid tidpunkten för genomförandet av detta direktiv en frist om högst 12 månader från den tidpunkten att anpassa sig till den nya nationella lagstiftningen.
3. Grekland och Portugal tillåts att uppskjuta genomförandet av detta direktiv till senast den 1 april 1992.
Ett år före detta datum skall kommissionen rapportera till rådet om hur genomförandet av direktivet fortgår och om eventuella svårigheter som kan uppkomma för Grekland eller Portugal att genomföra direktivet per det datum som anges i föregående stycke.
Kommissionen skall, om så erfordras, föreslå att rådet förlänger uppskovet upp till fyra år.
Artikel 58
Medlemsstaterna skall se till att kommissionen erhåller uppgift om texterna till de viktigaste föreskrifterna som de antar inom det område som omfattas av detta direktiv.
Artikel 59
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 235 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
med beaktande av följande: En harmonisk utveckling av den ekonomiska verksamheten samt en varaktig och balanserad tillväxt inom gemenskapen som helhet är beroende av att det upprättas en gemensam marknad som fungerar tillfredsställande och erbjuder villkor som motsvarar dem som råder på den nationella marknaden. För att få till stånd denna gemensamma marknad och stärka dess enhet bör rättsliga grundvalar skapas som underlättar för fysiska personer, bolag och andra rättsliga enheter att anpassa sin verksamhet till gemenskapens ekonomiska villkor. Det är därför nödvändigt att dessa fysiska personer, bolag och andra rättsliga enheter kan samarbeta effektivt över gränserna.
Ett sådant samarbete kan möta svårigheter av rättslig, skattemässig eller psykologisk natur. Ett ändamålsenligt rättsligt instrument på gemenskapsnivå i form av en europeisk ekonomisk intressegruppering skulle bidra till att ovannämnda mål uppnås och behövs därför.
Fördraget innehåller inte tillräckliga bestämmelser för ett sådant rättsligt instrument.
En grupperings förmåga att anpassa sig till de ekonomiska villkoren bör garanteras genom en avsevärd handlingsfrihet för grupperingens medlemmar att reglera sina avtalsmässiga förbindelser och grupperingens interna organisation.
En gruppering skiljer sig från ett bolag främst i fråga om ändamålet, vilket endast är att underlätta eller utveckla medlemmarnas ekonomiska verksamhet för att göra det möjligt för dessa att förbättra sina egna resultat. På grund av denna stödjande karaktär måste grupperingens verksamhet ha samband med medlemmarnas ekonomiska verksamhet och får inte ersätta denna i sådan utsträckning att grupperingen t.ex. i förhållande till tredje man utövar en självständig yrkesmässig verksamhet, varvid begreppet ekonomisk verksamhet skall ges en vidsträckt tolkning.
Fysiska personer, bolag och andra rättsliga enheter bör enligt förordningens syfte i största möjliga utsträckning ha tillträde till denna företagsform. Förordningen hindrar dock inte att det på det nationella planet tillämpas rättsregler och/eller etiska regler som gäller utövningen av en verksamhet eller ett yrke.
Enbart denna förordning ger inte rätt att delta i en gruppering, även om villkoren som föreskrivs i förordningen är uppfyllda.
Förordningens bestämmelser om möjlighet att av hänsyn till allmänna intressen förbjuda eller begränsa rätten att delta i en gruppering inverkar inte på de rättsregler i medlemsstaterna som behandlar utövande av verksamhet och som kan föreskriva ytterligare förbud eller begränsningar eller annan kontroll eller tillsyn i fråga om rätten för fysiska personer, bolag eller andra rättsliga enheter eller kategorier därav att delta i en gruppering.
För att en gruppering skall kunna fylla sitt ändamål skall den ha rättskapacitet. Ett organ som är rättsligt skilt från grupperingens medlemmar skall representera grupperingen mot tredje man.
Skyddet för tredje man kräver en hög grad av offentlighet. Medlemmarna ansvarar obegränsat solidariskt för grupperingens skulder och andra förbindelser, inklusive skulder avseende skatter och sociala avgifter, dock utan att denna princip inverkar på rätten att genom ett särskilt avtal mellan grupperingen och en tredje man bestämma att ansvaret skall uteslutas eller begränsas i fråga om en eller flera medlemmar när det gäller en viss skuld eller någon annan förbindelse.
Frågor om fysiska personers rättsliga handlingsförmåga och rättskapacitet samt om juridiska personers rättskapacitet regleras av nationell lagstiftning.
Regler bör ges om särskilda grunder för upplösning av grupperingen, dock bör hänvisning ske till nationella rättsregler om likvidation och avslutning av denna.
En gruppering omfattas av bestämmelserna i nationell lagstiftning om obestånd och betalningsinställelse. Dessa bestämmelser kan ange ytterligare grunder för upplösning av grupperingen.
Denna förordning föreskriver att det endast är grupperingens medlemmar som skall beskattas för resultatet av grupperingens verksamhet. Därutöver tillämpas nationella skatteregler, bl.a. när det gäller fördelningen av vinst, taxeringsförfarandet och alla förpliktelser som medlemsstaternas skattelagstiftning innehåller.
I frågor som inte omfattas av denna förordning tillämpas medlemsstaternas rättsregler och gemenskapsrätten, t.ex. när det gäller
- social- och arbetsrätt,
- konkurrensrätt,
- immaterialrätt.
En gruppering är underkastad medlemsstaternas rättsregler om utövande av verksamheten och kontroll av denna. Om en gruppering eller dess medlemmar missbrukar eller kringgår en medlemsstats lagstiftning får medlemsstaten tillgripa lämpliga sanktioner.
Det står medlemsstaterna fritt att tillämpa eller anta lagar eller förordningar eller vidta administrativa åtgärder som inte strider mot tillämpningsområdet för eller syftet med denna förordning.
Denna förordning skall i sin helhet omedelbart träda i kraft. Tillämpningen av vissa bestämmelser skall dock senareläggas för att ge medlemsstaterna möjlighet att inrätta den administration inom sina respektive områden som behövs för registrering av grupperingarna och för att säkerställa att handlingar angående dessa blir offentliga. Från den dag förordningen tillämpas skall de grupperingar som bildas kunna verka utan territoriella inskränkningar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
De som avser att bilda en gruppering skall ingå ett avtal och låta registrera grupperingen enligt artikel 6.
1. Syftet med en grupperings verksamhet är att underlätta eller utveckla medlemmarnas ekonomiska verksamhet och att förbättra resultatet av denna verksamhet; en gruppering har inte till syfte att skapa vinst för egen del. En grupperings verksamhet skall knyta an till medlemmarnas ekonomiska verksamhet och får endast vara av understödjande karaktär i förhållande till den senare verksamheten.
2. En gruppering får därför inte
a) direkt eller indirekt utöva någon form av styrning eller kontroll över medlemmarnas egen verksamhet eller över något annat företags verksamhet, särskilt inte i personal-, finansierings- eller investeringsfrågor,
b) under några omständigheter, varken direkt eller indirekt, inneha andelar eller aktier av något slag i ett företag som är medlem i grupperingen; innehav av andelar eller aktier i andra företag tillåts endast i den mån det är nödvändigt för att syftet med grupperingen skall uppnås och om det sker för medlemmarnas räkning,
c) ha fler än 500 anställda,
d) utnyttjas av ett bolag för att lämna lån till ledningen i ett bolag eller till någon ledningen närstående person, om rätten att bevilja sådana lån är begränsad eller underkastad kontroll enligt medlemsstaternas bolagsrätt; en gruppering får inte heller utnyttjas för att föra över egendom mellan ett bolag och dess ledning eller någon ledningen närstående person utöver vad som är tillåtet enligt medlemsstaternas bolagsrätt; i denna bestämmelse avses med att lämna lån även att medverka i transaktioner med motsvarande verkan, och med egendom avses lös och fast egendom,
e) vara medlem av någon annan europeisk ekonomisk intressegruppering.
Artikel 4
1. Endast följande kan vara medlemmar i en gruppering:
a) Bolag som avses i artikel 58 andra stycket i fördraget och andra rättsliga enheter av offentligrättsligt eller privaträttsligt slag, som har bildats enligt en medlemsstats lagstiftning och som har sitt registrerade eller i lag bestämda säte samt sitt huvudkontor inom gemenskapen; om ett bolag eller en annan rättslig enhet enligt en medlemsstats lagstiftning inte behöver ha ett registrerat eller i lag bestämt säte, räcker det att bolaget eller den rättsliga enheten har sitt huvudkontor inom gemenskapen.
b) Fysiska personer som utövar industri-, handels-, hant- verks- eller jordbruksverksamhet eller ett fritt yrke eller annan verksamhet inom gemenskapen.
2. En gruppering skall omfatta minst
a) två bolag eller andra rättsliga enheter som avses i punkt 1 och som har sina huvudkontor i olika medlemsstater, eller
b) två fysiska personer som avses i punkt 1 och som bedriver sin huvudsakliga verksamhet i olika medlemsstater, eller
c) ett bolag eller någon annan rättslig enhet som avses i punkt 1 och en fysisk person, av vilka den förstnämnda har sitt huvudkontor i en medlemsstat och den senare utövar sin huvudsakliga verksamhet i någon annan medlemsstat.
3. En medlemsstat kan bestämma att grupperingar som enligt artikel 6 är intagna i den statens register inte får ha mer än 20 medlemmar. Med hänsyn därtill får en sådan medlemsstat även bestämma att enligt dess lagstiftning varje medlem i en rättslig enhet, som har bildats enligt den lagstiftningen och som inte är ett registrerat bolag, skall behandlas som en särskild medlem när det gäller medlemskap i en gruppering.
4. Varje medlemsstat kan med hänsyn till sina allmänna intressen förbjuda eller begränsa rätten för vissa kategorier av fysiska personer, bolag eller andra rättsliga enheter att delta i grupperingar.
Artikel 5
Ett avtal om att bilda en gruppering skall innehålla minst följande uppgifter:
a) Grupperingens namn, föregånget eller följt av antingen orden "europeisk ekonomisk intressegruppering" eller förkortningen "EEIG", om inte dessa ord eller denna förkortning redan ingår i namnet.
b) Grupperingens säte.
c) Föremålet för grupperingens verksamhet.
d) För varje medlem namn, firma, rättslig organisationsform, bostadsadress eller adress för säte samt i förekommande fall registreringsnummer och registreringsort.
e) Tiden för grupperingens bestånd, om inte denna tid är obestämd.
Artikel 6
I den stat där en gruppering har sitt säte skall den tas in i ett register enligt artikel 39.1.
Artikel 7
Avtalet om att bilda en gruppering skall ges in till det register som anges i artikel 6.
Följande handlingar och uppgifter skall också ges in till registret: a) Varje ändring i avtalet om att bilda grupperingen, däribland varje ändring i grupperingens sammansättning.
b) Uppgift om inrättande eller nedläggning av ett huvudkontor eller avdelningskontor för grupperingen.
c) Ett rättsligt avgörande som enligt artikel 15 fastställer eller tillkännager att grupperingen är ogiltig.
d) Uppgift om vem eller vilka som har utsetts till företagsledare för grupperingen, vederbörandes namn och övriga personuppgifter som krävs enligt lagstiftningen i den medlemsstat där registret förs, uppgift huruvida företagsledarna kan handla var för sig eller om de måste handla i förening samt uppgift om när uppdraget för en företagsledare har upphört.
e) Uppgift om när en medlem enligt artikel 22.1 har överlåtit sin andel eller en del av denna.
f) Ett beslut av medlemmarna varigenom grupperingen förklaras upplöst enligt artikel 31 eller ett rättsligt avgörande om upplösning enligt artikel 31 eller 32.
g) Uppgift om att enligt artikel 35 en eller flera likvidatorer har tillsatts för en gruppering, vederbörandes namn och övriga personuppgifter som krävs enligt lagstiftningen i den medlemsstat där registret förs samt uppgift om när uppdraget för en likvidator har upphört.
h) Uppgift om att likvidationen av en gruppering har avslutats enligt artikel 35.2.
i) Förslag till byte av säte enligt artikel 14.1.
j) Avtalsvillkor enligt artikel 26.2 som befriar en ny medlem från ansvar för skulder och andra förpliktelser som har uppkommit innan han antogs som medlem.
Artikel 8
Följande skall offentliggöras enligt artikel 39 i den tidning som där anges i punkt 1:
a) De obligatoriska uppgifter som enligt artikel 5 skall anges i avtalet om att bilda en gruppering och ändring i dessa uppgifter.
b) Registreringsnummer, datum och ort för registreringen samt uppgift om att denna har upphört.
c) I artikel 7 b-j avsedda handlingar och uppgifter.
De i a och b angivna uppgifterna skall offentliggöras i sin helhet. I c angivna handlingar och uppgifter skall offentliggöras antingen i sin helhet eller i form av ett utdrag eller ett meddelande om att de har givits in till registret enligt tillämplig nationell lagstiftning.
Artikel 9
1. De handlingar och uppgifter som skall offentliggöras på grund av denna förordning kan åberopas av en gruppering mot tredje man enligt vad som har bestämts i tillämplig nationell lagstiftning med stöd av artikel 3.5 och 3.7 i rådets direktiv 68/151/EEG av den 9 mars 1968 om samordning av de skyddsåtgärder som krävs i medlemsstaterna av de i artikel 58 andra stycket i Romfördraget avsedda bolagen i bolagsmännens och tredje mans intressen, i syfte att göra skyddsåtgärderna likvärdiga inom gemenskapen (4).
2. Har handlingar företagits i en grupperings namn innan grupperingen registrerats enligt artikel 6 och åtar sig inte grupperingen efter registreringen att svara för de förbindelser som följer med dessa handlingar, svarar de fysiska personer, bolag eller andra rättsliga enheter som har företagit handlingarna obegränsat solidariskt för dessa.
Artikel 10
Ett huvudkontor eller avdelningskontor i någon annan medlemsstat än den där grupperingen har sitt säte skall registreras i den stat där kontoret är beläget. För detta ändamål skall grupperingen till den sistnämnda statens register ge in kopior av de handlingar som måste ges in till registret i den medlemsstat där grupperingen har sitt säte och, om det behövs, en översättning som uppfyller kraven vid det register där kontoret skall registreras.
Artikel 11
Efter offentliggörandet i den i artikel 39.1 avsedda tidningen skall i Europeiska gemenskapernas officiella tidning föras in uppgifter om bildandet av en gruppering och om avslutandet av en grupperings likvidation med uppgift om grupperingens registreringsnummer, datum och plats för registreringen, datum och plats för offentliggörandet samt den förstnämnda tidningens namn.
Artikel 12
Det säte som anges i avtalet om att bilda en gruppering skall finnas inom gemenskapen.
Sätet skall vara beläget
a) i den ort där grupperingen har sitt huvudkontor, eller
b) i den ort där någon av grupperingens medlemmar har sitt huvudkontor eller, när det är fråga om en fysisk person, utövar sin huvudsakliga verksamhet, förutsatt att grupperingen är verksam där.
Artikel 13
En gruppering får byta säte inom gemenskapen.
Beslut om bytet skall fattas enligt vad som är bestämt i avtalet om att bilda grupperingen, om inte bytet medför att enligt artikel 2 någon annan lagstiftning blir tillämplig.
Artikel 14
1. Om byte av säte medför att enligt artikel 2 någon annan lagstiftning blir tillämplig, skall förslag till bytet upprättas samt ges in och offentliggöras enligt föreskrifterna i artiklarna 7 och 8.
Beslut om bytet får fattas först två månader efter det att förslaget har offentliggjorts. Beslutet fattas enhälligt av medlemmarna. Det får verkan från den dag då grupperingen enligt artikel 6 tas in i det nya registret. Innan registreringen äger rum måste det visas att förslaget till byte har offentliggjorts.
2. En gruppering får avföras ur det tidigare registret först sedan det visats att grupperingen har tagits in i det nya registret.
3. Sedan den nya registreringen har offentliggjorts kan det nya sätet åberopas mot tredje man enligt artikel 9.1; innan grupperingens avförande ur det tidigare registret har offentliggjorts får dock tredje man fortfarande åberopa det tidigare sätet, om grupperingen inte visar att tredje man kände till det nya.
4. En medlemsstat kan i fråga om grupperingar som enligt artikel 6 är registrerade i den staten föreskriva i sin lagstiftning att ett byte av säte, som skulle medföra att annan lagstiftning blev tillämplig, inte skall få verkan om en behörig myndighet i den nämnda staten motsätter sig bytet inom den i punkt 1 angivna tvåmånadersfristen. En sådan invändning får endast grunda sig på allmänna intressen. Den skall kunna prövas av domstol.
Artikel 15
1. Om en gruppering är ogiltig på grund av den lagstiftning som enligt artikel 2 är tillämplig, skall ogiltigheten fastställas eller tillkännages genom avgörande av en domstol. Den domstol som handlägger saken skall dock bestämma en frist inom vilken rättelse får ske, om grupperingens förhållanden kan bringas i överensstämmelse med gällande rätt.
2. En grupperings ogiltighet medför likvidation av grupperingen enligt artikel 35.
3. Ett avgörande varigenom ogiltigheten av en gruppering fastställs eller tillkännages kan göras gällande mot tredje man enligt artikel 9.1.
Ett sådant avgörande enbart inverkar inte på giltigheten av de förpliktelser som grupperingen har ådragit sig eller som gäller till förmån för denna, om förpliktelserna har uppkommit innan avgörandet enligt föregående stycke kan göras gällande mot tredje man.
Artikel 16
1. Medlemmarna gemensamt och en eller flera företagsledare utgör grupperingens organ.
Avtalet om att bilda grupperingen kan innehålla bestämmelser om andra organ; i så fall skall avtalet ange dessas befogenheter.
2. Grupperingens medlemmar kan i egenskap av organ för denna fatta alla beslut som syftar till att förverkliga ändamålet med grupperingen.
Artikel 17
1. Varje medlem har en röst. Avtalet om att bilda grupperingen kan dock tilldela vissa medlemmar flera röster förutsatt att ingen medlem får röstmajoritet.
2. Medlemmarna kan endast enhälligt besluta att
a) ändra föremålet för grupperingens verksamhet,
b) ändra det antal röster som varje medlem har tilldelats,
c) ändra förutsättningarna för att fatta beslut,
d) förlänga grupperingens varaktighet utöver den tid som har bestämts i avtalet om att bilda grupperingen,
e) ändra det belopp med vilket varje medlem eller vissa medlemmar skall bidra till grupperingens finansiering,
f) ändra någon annan förpliktelse som åligger en medlem, om inte annat är bestämt i avtalet om att bilda grupperingen,
g) vidta andra ändringar i avtalet om att bilda grupperingen än som anges i denna punkt, om inte annat är bestämt i avtalet.
Artikel 18
Varje medlem har rätt att få upplysningar av företagsledarna om grupperingens verksamhet samt att granska grupperingens böcker och affärshandlingar.
Artikel 19
1. En gruppering leds av en eller flera fysiska personer som utses i avtalet om att bilda grupperingen eller genom beslut av medlemmarna.
Till företagsledare i en gruppering kan inte utses någon som
- enligt den lagstiftning som gäller för honom, eller
- enligt den interna lagstiftningen i den stat där grupperingen har sitt säte, eller
- enligt ett avgörande av domstol eller annan myndighet som har beslutats eller erkänts inom en medlemsstat
inte får tillhöra styrelsen eller direktionen i ett bolag, inte får leda ett företag eller inte får vara företagsledare i en europeisk ekonomisk intressegruppering.
2. En medlemsstat kan för grupperingar som enligt artikel 6 är intagna i den statens register föreskriva att en juridisk person får vara företagsledare, under förutsättning att denne till sina representanter utser en eller flera fysiska personer för vilka bestämmelserna i artikel 7 d skall gälla.
En medlemsstat som begagnar sig av den nu angivna möjligheten skall föreskriva att representanterna skall ha samma ansvar som företagsledarna.
Förbuden enligt punkt 1 gäller också för representanterna.
3. Förutsättningarna för att utse och entlediga företagsledarna samt dessas befogenheter skall bestämmas i avtalet om att bilda grupperingen eller genom enhälligt beslut av medlemmarna.
Artikel 20
1. Endast företagsledaren eller, om de är flera, var och en av dem företräder grupperingen mot tredje man.
När en företagsledare handlar på grupperingens vägnar förpliktar han denna mot tredje man även om hans handlingar faller utanför föremålet för grupperingens verksamhet, såvida inte grupperingen visar att tredje man kände till eller med hänsyn till omständigheterna inte kunde vara obekant med att handlingen föll utanför föremålet för grupperingens verksamhet; enbart offentliggörandet av den i artikel 5 c angivna uppgiften skall därvid inte anses tillräckligt som bevis.
En begränsning i företagsledarnas rätt att företräda grupperingen i avtalet om att bilda denna eller genom beslut av medlemmarna får inte åberopas mot tredje man, även om begränsningen har offentliggjorts.
2. I avtalet om att bilda grupperingen kan bestämmas att endast två eller flera företagsledare i förening får företräda denna. En sådan bestämmelse kan göras gällande mot tredje man enligt artikel 9.1 endast om den har offentliggjorts enligt artikel 8.
Artikel 21
1. Vinsten av en grupperings verksamhet skall anses som medlemmarnas egen vinst och delas mellan dem enligt vad som är bestämt i avtalet om att bilda grupperingen eller, om sådana bestämmelser saknas, i lika delar.
2. Grupperingens medlemmar skall bidra till att betala belopp varmed utgifterna överstiger inkomsterna enligt vad som är bestämt i avtalet om att bilda grupperingen eller, om sådana bestämmelser saknas, med lika delar.
Artikel 22
1. Varje medlem i en gruppering kan överlåta sin andel i denna eller en del av andelen till någon annan medlem eller till tredje man; överlåtelsen får verkan endast om grupperingens övriga medlemmar enhälligt har tillåtit denna.
2. En medlem kan endast med de övriga medlemmarnas enhälliga medgivande använda sin andel i grupperingen som säkerhet, om inte något annat är bestämt i avtalet om att bilda grupperingen. Innehavaren av en sådan säkerhet kan inte bli medlem på grund av säkerheten.
Artikel 23
En gruppering får inte rikta placeringserbjudanden till allmänheten. Artikel 24
1. Medlemmarna svarar obegränsat solidariskt för alla grupperingens förbindelser. Följderna av detta ansvar bestäms av den nationella lagstiftningen.
2. Innan likvidationen av en gruppering är avslutad får grupperingens borgenärer inte väcka talan mot en medlem för att få betalt enligt punkt 1, om de inte först har anmodat grupperingen att betala och betalning inte har erlagts inom skälig tid.
Artikel 25
På brev, beställningssedlar och liknande handlingar skall följande tydligt anges:
a) Grupperingens namn föregånget eller följt av orden "europeisk ekonomisk intressegruppering" eller förkortningen "EEIG", om inte orden eller förkortningen redan ingår i namnet.
b) Orten för det register enligt artikel 6 i vilket grupperingen är införd och grupperingens registreringsnummer.
c) Adressen för grupperingens säte.
d) I förekommande fall att företagsledarna endast får handla i förening.
e) I förekommande fall att grupperingen har trätt i likvidation enligt artikel 15, 31, 32 eller 36.
Varje enligt artikel 10 registrerat kontor skall på de nu nämnda handlingarna som härrör från kontoret lämna de angivna uppgifterna och motsvarande uppgifter som gäller kontorets egen registrering.
Artikel 26
1. Ett beslut att anta en ny medlem skall fattas enhälligt av medlemmarna.
2. Varje ny medlem svarar enligt artikel 24 för grupperingens förbindelser, inräknat sådana som har uppkommit i verksamheten före medlemmens inträde.
En medlem kan dock genom en bestämmelse i avtalet om att bilda grupperingen eller i inträdeshandlingen fritas från ansvar för förbindelser som har uppkommit före inträdet. En sådan bestämmelse kan göras gällande enligt artikel 9.1 mot tredje man, om den har offentliggjorts enligt artikel 8.
Artikel 27
2. En medlem kan uteslutas på de grunder som anges i avtalet om att bilda grupperingen och under alla förhållanden, om medlemmen väsentligt åsidosätter sina skyldigheter eller vållar eller hotar att vålla allvarliga störningar i grupperingens verksamhet.
En sådan uteslutning får ske endast genom ett domstolsavgörande efter gemensam ansökan av en majoritet av de övriga medlemmarna, om inte något annat är bestämt i avtalet om att bilda grupperingen.
Artikel 28
1. Ett medlemskap upphör när medlemmen dör eller inte längre uppfyller de i artikel 4.1 angivna villkoren.
Dessutom kan en medlemsstat med hänsyn till sin lagstiftning om upplösning, likvidation, obestånd och betalningsinställelse bestämma att ett medlemskap skall upphöra vid tidpunkter som anges i den nämnda lagstiftningen.
2. Om en medlem dör, kan någon annan inträda i grupperingen i den avlidnes ställe endast på de villkor som är bestämda i avtalet om att bilda grupperingen eller efter samtycke av alla övriga medlemmar.
Artikel 29
Så snart någon upphör att vara medlem skall företagsledarna underrätta de övriga medlemmarna om det; företagsledarna skall dessutom vidta de åtgärder som krävs enligt artiklarna 7 och 8. De sistnämnda åtgärderna får även vidtas av var och en som saken angår.
Artikel 30
Utom då avtalet att bilda grupperingen föreskriver något annat och med förbehåll för den rätt som någon kan ha förvärvat enligt artiklarna 22.1 och 28.2, skall grupperingen efter det att ett medlemskap har upphört fortsätta att bestå med de kvarvarande medlemmarna och på de villkor som är bestämda i avtalet om att bilda grupperingen eller som de sistnämnda medlemmarna enhälligt beslutar.
Artikel 31
1. En gruppering får upplösas genom ett beslut av medlemmarna om detta. Ett sådant beslut skall fattas enhälligt om inte något annat är bestämt i avtalet om att bilda grupperingen. 2. En gruppering skall upplösas genom ett beslut av medlemmarna, om
a) tiden för grupperingens bestånd enligt avtalet om att bilda denna har löpt ut eller någon annan i avtalet angiven grund för upplösning föreligger, eller
b) ändamålet med grupperingen har uppnåtts eller inte längre kan uppnås.
Varje medlem får ansöka om att rätten skall bestämma att upplösning skall ske, om medlemmarna ännu tre månader efter det att en i a eller b angiven omständighet har inträffat inte har beslutat om upplösning.
3. En gruppering skall även upplösas genom ett beslut av medlemmarna eller den kvarvarande medlemmen om de i artikel 4.2 angivna villkoren inte längre är uppfyllda.
4. Efter upplösning av en gruppering genom beslut av medlemmarna skall företagsledarna vidta de åtgärder som krävs enligt artiklarna 7 och 8. Dessa åtgärder får även vidtas av var och en som saken angår.
Artikel 32
1. På ansökan av den som saken angår eller en behörig myndighet skall rätten förordna att en gruppering skall upplösas om bestämmelserna i artikel 3, 12 eller 31.3 har åsidosatts, såvida inte rättelse vidtas innan rätten har avgjort ärendet.
2. På ansökan av en medlem får rätten förordna att en gruppering skall upplösas, om det föreligger en riktig grund för det.
3. En medlemsstat kan bestämma att rätten på ansökan av en behörig myndighet inom den staten får förordna att en gruppering med säte inom staten skall upplösas om grupperingen åsidosätter allmänna intressen inom staten, allt under förutsättning att det enligt statens lagstiftning är möjligt att på sådan grund upplösa registrerade bolag eller andra rättsliga enheter.
Artikel 33
Om någon upphör att vara medlem i en gruppering på annan grund än överlåtelse av rättigheter enligt artikel 22.1, skall värdet av den avgående medlemmens rättigheter och skyldigheter bestämmas med hänsyn till grupperingens förmögenhetsförhållanden vid tidpunkten för medlemskapets upphörande.
Värdet av en avgående medlems rättigheter och skyldigheter får inte bestämmas i förväg.
Artikel 34
Med den begränsning som anges i artikel 37.1 svarar en avgången medlem enligt artikel 24 för de förbindelser som har uppkommit genom grupperingens verksamhet före avgången.
Artikel 35
1. Avvecklingen av en gruppering skall ske genom likvidation.
2. Likvidationen och avslutningen av denna skall ske enligt nationell rätt.
3. Grupperingen behåller sin rättskapacitet enligt artikel 1.2 till dess likvidationen är avslutad.
4. Likvidatorerna skall vidta de åtgärder som avses i artiklarna 7 och 8.
Artikel 36
En gruppering omfattas av nationell lagstiftning om obestånd och betalningsinställelse. Enbart det förhållandet att ett rättsligt förfarande inleds mot en gruppering på grund av dennas obestånd eller betalningsinställelse får inte medföra att ett sådant förfarande inleds mot medlemmarna.
Artikel 37
1. En preskriptionstid på fem år räknat från offentliggörandet enligt artikel 8 av en medlems avgång gäller i stället för längre preskriptionstider i nationell lagstiftning i fråga om åtgärder mot den avgångne medlemmen med anledning av förbindelser som har uppkommit genom grupperingens verksamhet före avgången.
2. En preskriptionstid på fem år räknat från offentliggörandet enligt artikel 8 av avslutandet av en grupperings likvidation gäller i stället för längre preskriptionstider i nationell lagstiftning i fråga om åtgärder mot en medlem med anledning av förbindelser som har uppkommit genom grupperingens verksamhet.
Artikel 38
En behörig myndighet i en medlemsstat får förbjuda en gruppering att utöva verksamhet varigenom grupperingen åsidosätter allmänna intressen i den staten. Förbudet skall kunna prövas av domstol. Artikel 39
1. Medlemsstaterna skall inrätta det eller de register som skall svara för registrering enligt artiklarna 6 och 10, samt meddela regler om registreringen. De skall bestämma hur handlingarna som avses i artiklarna 7 och 10 skall ges in. De skall se till att de handlingar och uppgifter som avses i artikel 8 offentliggörs i en lämplig officiell tidning inom den medlemsstat där grupperingen har sitt säte, samt får bestämma hur de handlingar och uppgifter som avses i artikel 8 c skall offentliggöras.
Medlemsstaterna skall vidare se till att var och en har möjlighet att vid det register som avses i artikel 6 respektive 10 ta del av de i artikel 7 angivna handlingarna och att, även med post, få fullständiga eller partiella kopior av dessa handlingar.
Medlemsstaterna får bestämma att avgifter skall erläggas för den verksamhet som avses i de två föregående styckena; avgifterna får dock inte överstiga de administrativa kostnaderna för verksamheten.
2. Medlemsstaterna skall se till att de upplysningar som enligt artikel 11 skall offentliggöras i Europeiska gemenskapernas officiella tidning sänds till kontoret för de Europeiska gemenskapernas officiella publikationer inom en månad efter offentliggörandet i den officiella tidning som avses i punkt 1.
3. Medlemsstaterna skall bestämma lämpliga påföljder för underlåtenhet att iaktta föreskrifterna om offentliggörande i artiklarna 7, 8 och 10 och föreskrifterna i artikel 25.
Artikel 40
Endast medlemmarna skall beskattas för resultatet av en grupperings verksamhet.
Artikel 41
1. Medlemsstaterna skall före den 1 juli 1989 vidta de åtgärder som krävs av dem enligt artikel 39. De skall underrätta kommissionen så snart åtgärderna har vidtagits.
2. För kännedom skall en medlemsstat underrätta kommissionen om vilka kategorier av fysiska personer, bolag och andra rättsliga enheter som medlemsstaten enligt artikel 4.4 har förbjudit att delta i en gruppering. Kommissionen skall underrätta de övriga medlemsstaterna om förbudet.
Artikel 42
1. När denna förordning har antagits skall en kontaktkommitté tillsättas under kommissionens överinseende. Kontaktkommitténs uppgift skall vara att
a) med förbehåll för artiklarna 169 och 170 i Romfördraget underlätta tillämpningen av förordningen genom regelbundet samråd, särskilt om praktiska problem i samband med tillämpningen,
b) vid behov ge kommissionen råd om tillägg till eller ändringar i förordningen.
2. Kontaktkommittén skall bestå av representanter för medlemsstaterna och kommissionen. En representant för kommissionen skall vara ordförande. Kommissionen skall tillhandahålla ett sekretariat.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1035/72/EEG(1) av den 18 maj 1972 om den gemensamma organisationen av marknaden för frukt och grönsaker, senast ändrad genom förordning (EEG) nr 1332/84(2),
med beaktande av rådets förordning (EEG) nr 449/69 av den 11 mars 1969 om återbetalning av stöd som medlemsstaterna har beviljat frukt- och grönsaksproducenters organisationer(3), särskilt artikel 7.3 i denna, och
med beaktande av följande: Genom rådets förordning (EEG) nr 3284/83(4) ändras bestämmelserna för beviljande av stöd till frukt- och grönsaksproducenters organisationer.
De blanketter som avses i rådets förordning (EEG) nr 850/80(5) bör därför anpassas till de nya bestämmelserna.
Det åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för Europeiska utvecklings- och garantifonden för jordbruket.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Enda artikel
Bilagorna 1 och 2 i rådets förordning (EEG) nr 2264/69(6) skall ersättas med bilagorna 1 och 2 till denna förordning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av Anslutningsakten för Spanien och Portugal, särskilt artiklarna 171 och 358 i denna,
med beaktande av rådets förordning (EEG) nr 3117/85 av den 4 november 1985 om allmänna bestämmelser för beviljande av ekonomisk kompensation avseende sardiner(), särskilt artikel 4 i denna, och
med beaktande av följande: I artikel 2 i förordning (EEG) nr 3117/85 fastställs vissa villkor för beviljande av ekonomisk kompensation för produkterna, att den kvantitativa begränsningen skall vara 2 000 ton, vilka mottagarna av stödet skall vara samt metoden för beräkning av detta.
Detta program måste tillämpas på de kategorier av sardiner som kan förutses vara lättast att avsätta på marknaden efter beredning.
De hygienföreskrifter och tekniska bestämmelser som fastställts av de nationella myndigheterna bör säkerställa att produkterna i fråga fullständigt och slutligt beretts i någon av de former som anges i artikel 3.1 i förordning (EEG) nr 3117/85. Det bör kontrolleras att de beredda produkterna överensstämmer med dessa bestämmelser.
De former av beredning som är tillåtna bör preciseras i syfte att klart ange omfattningen av den aktuella ordningen.
När det gäller de kvantiteter som berättigar till bidrag bör närmare bestämmelser införas för hur ansökningarna om utbetalning av bidraget skall lämnas in.
För att kunna möjliggöra en fortlöpande kontroll bör bidragsmottagarna hela tiden hålla tillsynsmyndigheten underrättad om sin beredningsverksamhet.
Enligt artikel 2.3 i anslutningsfördraget får gemenskapens institutioner före anslutningen vidta de åtgärder som anges i artiklarna 171 och 358 i akten.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fiskeriprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- fångats av medlemmarna,
- sålts till en beredare för fullständig och slutlig beredning i enlighet med de hygienföreskrifter och tekniska bestämmelser som gäller för livsmedelsprodukter i den medlemsstat där beredaren är etablerad.
2. De beredningsprocesser som avses i punkt 1 är
a) frysning,
b) framställning av konserver enligt nr 16.04 i gemensamma tulltaxan,
c) filetering eller styckning i förening med en av de beredningsformer som avses i a och b.
Artikel 3
För varje parti av samma kommersiella kategori som säljs skall bidragets storlek bestämmas i enlighet med artikel 2.4 i förordning (EEG) nr 3117/85.
Artikel 4
Om någon av de beredningsprocesser som anges i artikel 2.2 utförs i en annan medlemsstat än den som erkänt den producentorganisation som säljer produkten, skall bevis om att sådan beredning ägt rum företes i form av kontrollformulär T nr 5 i enlighet med bestämmelserna i kommissionens förordning (EEG) nr 223/77() och i denna förordning.
Av kontrollformuläret skall följande uppgifter framgå:
- I fält 41 en beskrivning av varorna i det tillstånd de befann sig vid tidpunkten för avsändandet.
- I fält 104 en av följande angivelser med versaler:
"VERARBEITUNG, FÜR DIE EINE AUSGLEICHS- ENTSCHÄDIGUNG GEWÄHRT WIRD
såvida det vid utbetalningstillfället inte finns uppgifter som tyder på att produkterna inte har beretts fullständigt och slutligt.
2. Beredaren skall skriftligt åta sig att bereda de produkter som ingår i avtalet i enlighet med bestämmelserna i artikel 2. Han måste därför i sin lagerförteckning kunna identifiera de kvantiteter som inköpts i samband därmed. Beredaren skall förplikta sig att upplåta sina lokaler för varje form av inspektion av de behöriga myndigheterna.
3. Producentorganisationen skall lämna in ansökan om utbetalning av bidraget till de behöriga myndigheterna i den berörda medlemsstaten före slutet av den första månaden efter det att försäljningsavtalet ingåtts.
Artikel 6
1. De berörda medlemsstaterna skall införa ett kontrollsystem för att säkerställa att de produkter för vilka ansökan om bidrag lämnats in berättigar till sådant och att bestämmelserna i denna förordning följts.
2. De närmare bestämmelserna för hur kontrollen skall gå till skall utarbetas av medlemsstaten och omfatta minst följande krav:
- Inspektioner av beredningsföretagen på plats.
- Mottagaren av bidraget skall lämna in de handlingar på vilka han grundar sina anspråk på rätt till bidraget.
- Närmare angivande av de uppgifter som skall ingå i den ansökan om bidrag som anges i artikel 5.
- Identifiering genom producentorganisationens försäljningsjournal av de kvantiteter som sålts enligt denna ordning.
Artikel 7
1. De berörda medlemsstaterna skall senast två månader efter ikraftträdandet av denna förordning anmäla till kommissionen vilka kontrollåtgärder som införts i enlighet med artikel 6.1.
2. Medlemsstaterna skall också varje månad till kommissionen anmäla de kvantiteter som sålts under den föregående månaden som berättigar till stöd, fördelade på handelskategorier och beredningsformer, samt kostnaderna för beviljandet av stödet i fråga.
3. På grundval av den information som framkommit vid kontrollen enligt artikel 6 skall i förekommande fall bidragets storlek korrigeras.
Artikel 8
Den omvandlingskurs som skall gälla för bidraget är den på försäljningsdagen gällande representativa kursen.
Artikel 9
Denna förordning träder i kraft den 1 mars 1986, förutsatt att Anslutningsfördraget för Spanien och Portugal då trätt i kraft. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), senast ändrad genom förordning (EEG) nr 1298/85(2), särskilt artikel 6.7 i denna, och
med beaktande av följande: I kommissionens förordning (EEG) nr 3143/85 av den 11 november 1985 om försäljning till sänkt pris av interventionssmör för användning till direkt konsumtion i form av koncentrerat smör(3), senast ändrad genom förordning (EEG) nr 3338/85(4), föreskrivs att förpackningar med koncentrerat smör skall vara försedda med vissa påskrifter som är skrivna med klart synliga och läsliga tryckbokstäver. På grund av ett fel motsvarar påskriften på italienska språket inte den påskrift som antagits i den text som förelagts Förvaltningskommittén för mjölk och mjölkprodukter för röstning. Följaktligen bör nämnda förordning rättas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 5.4 första stycket skall den näst sista strecksatsen ersättas med följande:
"- burro concentrato".
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS BESLUT av den 22 december 1986 om införande av en ordning för samråd och samarbete på turistområdet (86/664/EEG)
med beaktande av kommissionens förslag (),
med beaktande av Europaparlamentets yttrande (),
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
med beaktande av följande: Enligt artikel 2 i fördraget har gemenskapen särskilt till uppgift att främja en harmonisk utveckling av den ekonomiska verksamheten inom gemenskapen som helhet, en fortgående och balanserad tillväxt, en ökad stabilitet, samt närmare förbindelser mellan de stater som gemenskapen förenar. Turism kan bidra till att uppnå dessa mål.
Rådets resolution av den 10 april 1984 om gemenskapspolitik på turistområdet () understryker behovet av samråd mellan medlemsstaterna och kommissionen i fråga om turism.
Samråd är ett bra medel för att underlätta samarbetet mellan medlemsstaterna och kommissionen i avsikt att uppnå fördragets mål.
Varje medlemsstat bör låta de andra medlemsstaterna och kommissionen dra fördel av sin erfarenhet inom turistområdet.
I avsikt att ha samråd inom turistområdet bör informationsutbyte säkerställas mellan medlemsstaterna och kommissionen.
Sådant samråd bör inte upprepa det arbete som utförts inom andra gemenskapsorgan.
HÄRIGENOM FÖRESKRIVS FÖLJANDE
Artikel 1
En rådgivande turistkommitté, härefter kallad "kommittén", skall inrättas hos kommissionen. Den skall bestå av medlemmar utsedda av varje medlemsstat.
Artikel 2
Kommitténs uppgift skall vara att underlätta informationsutbyte, samråd och, när så är lämpligt, samarbete om turism och då i synnerhet tjänster för turister.
Artikel 3
För de ändamål som anges i artikel 2 skall varje medlemsstat översända en rapport till kommissionen en gång om året om de viktigaste åtgärderna som den har vidtagit och, så långt möjligt, om de åtgärder den avser att vidta i fråga om sådana tjänster för turister som skulle kunna få konsekvenser för resande från andra medlemsstater.
Kommissionen skall underrätta de andra medlemsstaterna om detta.
Artikel 4
3. Kommittén skall också råda kommissionen i de frågor där kommissionen har begärt ett yttrande.
4. Den information och det samråd som föreskrivs i detta beslut skall omfattas av tystnadsplikt.
Artikel 5
Kommissionen skall utöva ordförandeskapet i kommittén.
Kommissionen skall tillhandahålla sekreterartjänster åt kommittén.
med beaktande av Anslutningsakten för Spanien och Portugal, särskilt artikel 396 i denna, och
med beaktande av följande: Med anledning av Portugals anslutning är det nödvändigt att göra vissa ytterligare tekniska ändringar av direktiv 85/384/EEG() i dess lydelse enligt direktiv 85/614/EEG() för att säkerställa att det tillämpas på samma sätt av Portugal och de andra medlemsstaterna.
I enlighet med artikel 2.3 i Fördraget om Spaniens och Portugals anslutning får gemenskapens institutioner besluta om de åtgärder som åsyftas i artikel 396 i anslutningsakten, vilka åtgärder skall träda i kraft om och när fördraget träder i kraft.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Med verkan från den 1 januari 1986 skall artikel 11 k i direktiv 85/384/EEG kompletteras med följande:
med beaktande av rådets förordning (EEG) nr 426/86 av den 24 februari 1986 om den gemensamma organisationen av marknaden för bearbetade produkter av frukt och grönsaker (), särskilt artikel 6.4 i denna, och
med beaktande av följande: I artikel 2.1 i förordning (EEG) nr 426/86 föreskrivs ett system för produktionsstöd för vissa produkter. I artikel 6.1 b i samma förordning föreskrivs att stödet endast skall betalas ut för produkter som uppfyller vissa minimikvalitetskrav som skall fastställas.
Syftet med sådana minimikrav på kvalitet är att förhindra framställning av produkter som inte efterfrågas eller produkter som skulle leda till en snedvridning av marknaden. Kraven måste baseras på traditionella och sunda framställningsmetoder.
Med tanke på genomförandet av systemet med produktionsstöd måste denna förordning tillämpas tillsammans med kommissionens förordning (EEG) nr 1599/84 av den 5 juni 1984 om tillämpningsföreskrifter för produktionsstödet för bearbetade produkter av frukt och grönsaker (), senast ändrad genom förordning (EEG) nr 1155/86 (), särskilt vad gäller undersökning av de bearbetade produkterna.
De kvalitetskrav som fastställs i denna förordning ingår i åtgärderna för genomförandet av systemet med produktionsstöd. Gemenskapen har ännu inte fastställt kvalitetskraven i samband med saluföring av produkterna. Medlemsstaterna får för detta ändamål fortsätta att tillämpa nationella krav under förutsättning att de är förenliga med fördragets bestämmelser om fri rörlighet för varor.
Förvaltningskommittén för bearbetade produkter av frukt och grönsaker har inte lämnat något yttrande inom den tidsfrist som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Denna förordning fastställer de minimikvalitetskrav som produkter som framställs av tomater enligt definitionen i artikel 1.2 i förordning (EEG) nr 1599/84 skall uppfylla för att få del av det produktionsstöd som avses i artikel 2.1 i förordning (EEG) nr 426/86.
Artikel 2
Artikel 3
I denna avdelning betyder "skalade tomater"
P hela tomater eller tomater i bitar, skalade och konserverade enligt definitionen i artikel 1.2 h, ij, k och l i förordning (EEG) nr 1599/84.
Artikel 4
1. Skalade tomater får endast tillsättas
P vatten,
P tomatsaft,
P tomatkoncentrat,
P vanligt salt (natriumklorid),
P naturliga kryddor, kryddörter och extrakt av dessa samt naturliga aromämnen.
Som tillsatsämnen vid framställning av skalade tomater får endast citronsyra (E 330) och kalciumklorid (509) användas.
2. Den totala tillsatsen av vanligt salt får inte överstiga 3 % av nettovikten och vid tillsättning av kalciumklorid får det totala kalciuminnehållet inte överstiga 0,045 % i hela tomater och 0,080 % i tomater i bitar. Vid bestämningen av tillsatsen vanligt salt skall det naturliga kloridinnehållet anses vara lika med 2 % av torrsubstansen.
3. Tillsatt tomatsaft och tomatkoncentrat skall uppfylla de minimikrav som fastställs i avdelning II.
Artikel 5
1. Skalade tomater skall vara fria från främmande smaker och lukter och färgen skall vara karakteristisk för den sort som används och för korrekt bearbetade skalade tomater.
2. Skalade tomater skall vara praktiskt taget fria från skal. Hela skalade tomater skall dessutom vara praktiskt taget fria från skadade delar.
3. Mögeltalet för skalade tomater (tomaterna och den omgivande vätskan) skall inte överstiga 50 % positiva fält och pH-värdet får inte överstiga 4,5.
Artikel 6
1. Produkterna skall anses uppfylla kraven i artikel 5.2 om följande gränsvärden för skador inte överskrids:
P skador: 35 cm2 sammantagen yta,
P skal:
P hela tomater: 300 cm2 sammantagen yta,
P tomater i bitar: 1 250 cm2 sammantagen yta.
De fastställda gränsvärdena gäller per 10 kg nettovikt.
2. I punkt 1 avses med
a) skador: områden där skador på ytan har trängt igenom och som därigenom skiljer sig starkt i färg eller konsistens från den normala tomatvävnaden och som normalt borde ha avlägsnats under bearbetningen,
b) skal: både skal som sitter fast på tomatköttet och skal som påträffas löst i behållaren.
Artikel 7
1. Vad avser skalade konserverade tomater skall tomaterna och den omgivande vätskan uppta minst 90 % av behållarens volym.
2. Den avrunna nettovikten för hela skalade tomater skall i genomsnitt vara lika med minst 56 % av behållarens volym uttryckt i gram.
3. Om skalade konserverade tomater förpackas i glasburkar skall volymen minskas med 20 ml innan de procenttal som avses i punkterna 1 och 2 beräknas.
Artikel 8
I denna avdelning skall "tomatsaft" och "tomatkoncentrat" avse de produkter som definieras i artikel 1.2 n och o i förordning (EEG) nr 1599/84.
Artikel 9
1. Tomatsaft och tomatkoncentrat får endast tillsättas följande:
P vanligt salt (natriumklorid),
P naturliga kryddor, kryddörter och extrakt av dessa samt naturliga aromämnen.
2. Som tillsatsämne vid framställning av tomatsaft och tomatkoncentrat får citronsyra (E 330) användas. Vidare, vid framställning av
P tomatsaft med ett torrsubstansinnehåll på mindre än 7 %, får askorbinsyra (E 300) användas. Innehållet av askorbinsyra skall dock inte överstiga 0,03 % av den färdiga produktens vikt,
P tomatkoncentrat i pulverform, får kiseldioxid (551) användas. Innehållet av kiseldioxid skall dock inte överstiga 1 % av den färdiga produktens vikt.
3. Kvantiteten tillsatt vanligt salt får inte överstiga
a) 15 viktprocent av torrsubstansinnehållet i tomatkoncentrat med ett torrrsubstansinnehåll som överstiger 20 %, och
b) 3 viktprocent av nettovikten för andra tomatkoncentrat och för tomatsaft.
Vid bestämning av kvantiteten tillsatt vanligt salt skall det naturliga innehållet av klorider anses vara lika med 2 % av torrsubstansinnehållet.
Artikel 10
1. Tomatsaft och tomatkoncentrat skall ha
a) en karakteristisk röd färg, och
b) en god smak som är karakteristisk för en korrekt bearbetad produkt.
Produkterna skall vara fria från främmande smaker, särskilt smaken av bränd eller karamelliserad produkt. 2. Tomatsaft och tomatkoncentrat skall vara
a) fria från synligt främmande beståndsdelar av vegetabiliskt ursprung, däribland skal, frön och andra hårda delar av tomater,
b) praktiskt taget fria från oorganiska orenheter.
3. De krav som fastställs i punkt 2 skall anses vara uppfyllda om
a) eventuella främmande beståndsdelar av vegetabiliskt ursprung endast kan urskiljas genom en noggrann undersökning med blotta ögat, och
b) halten av oorganiska orenheter inte överstiger 0,1 % av torrsubstansinnehållet, reducerat med eventuell tillsats av vanligt salt och vad avser tomatkoncentrat i pulverform, eventuell tillsats av kiseldioxid.
4. Tomatsaft och tomatkoncentrat skall ha
a) en jämnt fördelad konsistens och beskaffenhet som visar att en korrekt bearbetningsmetod har använts,
b) en sockerhalt uttryckt som invertsocker på minst 42 viktprocent av torrsubstansinnehållet minskat med eventuell tillsats av vanligt salt,
c) en total titrerbar surhet, uttryckt som kristalliserad citronsyremonohydrat, på högst 10 viktprocent av torrsubstansinnehållet minskat med eventuell tillsats av vanligt salt,
d) en flyktig surhet, uttryckt som ättiksyra på högst 0,4 viktprocent av torrsubstansen, minskat med eventuell tillsats av vanligt salt,
e) ett pH-värde på högst 4,5.
5. Mögeltalet för tomatsaft och tomatkoncentrat skall, vid spädning med så mycket vatten att torrsubstanshalten uppgår till 8 %, inte överstiga 70 % positiva fält. För tomatsaft med en torrsubstanshalt på mindre än 8 %, skall procenttalet för positiva fält minskas i proportion till torrsubstanshalten.
Artikel 11
I denna avdelning skall "tomatflingor" avse den produkt som definieras i artikel 1.2 m i förordning (EEG) nr 1599/84.
Artikel 12
1. Tomatflingor skall
a) ha en karakteristisk röd färg, och
b) ha en god smak som är karakteristisk för en korrekt bearbetad produkt, och
c) vara fria från främmande smaker och lukter.
2. Tomatflingors torrsubstanshalt skall vara minst 93 %.
3. Det sammanlagda innehållet av oorganiska och vegetabiliska orenheter får inte överstiga 1 % av produktens vikt. Med "vegetabiliska orenheter" avses här ett material av vegetabiliskt ursprung som kan urskiljas med blotta ögat och som inte är en del av själva tomaten eller som har suttit fast vid den färska tomaten men skulle ha avlägsnats vid bearbetningen, särskilt blad, stjälkar och foderblad från tomatplantan.
4. Som tillsatsämne vid framställning av tomatflingor får endast kiseldioxid (551) användas. Kiseldioxidinnehållet får dock inte överstiga 1 viktprocent.
Artikel 13
1. Behållare med konserverade skalade tomater, hela eller i bitar, och tomatsaft skall märkas med en referens som anger tillverkningsdatum och -år samt bearbetningsföretag. Om tomatsaft som har producerats på olika dagar har lagrats tillsammans innan den förpackas skall märkningen göra det möjligt att fastställa alla tillverkningsdagarna.
2. Bestämmelserna i punkt 1 skall även gälla andra tomatbaserade produkter om sådana produkter vid bearbetningstillfället förpackas i behållare i vilka de skall lämna bearbetningsanläggningen. Om de förvaras i tankar eller liknande behållare ämnade för senare förpackning eller vidare bearbetning, skall datumet eller datumen för framställningen anges på behållarna. När sådana produkter förpackas i de slutliga behållarna skall det på dessa finnas en referens som gör det möjligt att fastställa datumet eller datumen för framställningen samt bearbetningsföretaget.
3. Märkningen som avses i denna artikel kan vara i form av en kod och skall godkännas av de behöriga myndigheterna i den medlemsstat där framställningen sker. Dessa myndigheter får fastställa ytterligare föreskrifter angående själva märkningen.
Artikel 14
Bearbetningsföretaget skall dagligen och med jämna mellanrum under bearbetningen kontrollera att produkterna uppfyller kraven för beviljande av stöd. Resultatet av kontrollen skall registreras. Artikel 15
1. I bilagan fastställs analysmetoderna för att bestämma
a) torrsubstansinnehållet,
b) naturliga lösliga substanser,
c) saltinnehållet,
d) sockerinnehållet,
e) den totala surheten,
f) innehållet av flyktiga syror,
g) innehållet av oorganiska orenheter,
h) pH-värde,
i) innehållet av kalciumjoner, och
3. De metoder som avses i punkterna 1 och 2 skall användas för att slutgiltigt fastställa om produktionsstöd skall beviljas. Andra metoder får användas för rutinmässiga analyser.
Artikel 16
Denna förordning träder i kraft den 1 juli 1986.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av följande: Artikel 30 och följande i fördraget, om avskaffande av kvantitativa restriktioner och alla åtgärder med motsvarande verkan, gäller utan åtskillnad för de varor som har sitt ursprung i gemenskapen och sådana som har övergått till fri omsättning i någon av medlemsstaterna oberoende av ursprung.
Enligt dessa regler är krav på importlicens eller liknande förfarande, även om de är rent formella, förbjudna i handeln mellan medlemsstaterna.
Dessutom utesluter artikel 9.2 i fördraget varje administrativt förfarande som är avsett att skapa olika regler för rörelse av varor, beroende på om varorna har sitt ursprung i gemenskapen eller i tredje land och har övergått till fri omsättning i någon av medlemsstaterna.
En fullständig tillämpning av dessa principer förutsätter emellertid en fungerande gemensam handelspolitik.
Genomförandet av en gemensam handelspolitik är ännu inte slutfört. Åtgärder från medlemsstaters sida för vissa varor från tredje land har ännu inte ersatts av enhetliga, gemensamma regler.
Att en gemensam handelspolitik ännu inte helt genomförts innebär att det fortfarande kommer att finnas skillnader mellan medlemsstaterna i fråga om handelspolitiken, vilket kan vålla störning i handeln, något som artikel 115 i fördraget är avsedd att hindra.
För detta ändamål har kommissionen befogenhet att til låta medlemsstater att, utan hinder av principen om fri rörlighet inom gemenskapen, besluta om övervakningsåtgärder eller skyddsåtgärder inom gemenskapen gentemot varor som har sitt ursprung i tredje land och som övergått till fri omsättning i någon av medlemsstaterna. I artikel 115 föreskrivs emellertid att sådana åtgärder enbart kan tillåtas om de är nödvändiga och att kommissionen skall ge företräde åt åtgärder som vållar de minsta störningarna när det gäller den gemensamma marknadens funktion. Följden är att på det nuvarande stadiet av genomförandet av den gemensamma marknaden åtgärder enligt artikel 115 i fördraget bör tillåtas endast i fall där en störning i handeln leder till ekonomiska svårigheter eller äventyrar effektiviteten av handelspolitiska åtgärder som medlemsstater har vidtagit i överensstämmelse med gemenskapens internationella åtaganden.
Enligt Europeiska enhetsakten kommer den 1 januari 1993 ett område utan inre gränser att upprättas inom vilket varor, tjänster och kapital fritt kan röra sig. Detta innebär å ena sidan att de kvarstående skillnaderna i medlemsstaternas handelspolitik gradvis kommer att försvinna eller minska, och å andra sidan att kommissionen måste vara fullt medveten om dessa mål när den bedömer behovet av att tillåta åtgärder enligt artikel 115 i fördraget. Genom kommissionens beslut 80/47/EEG av den 20 december 1979 om övervaknings- och skyddsåtgärder som medlemsstater kan tillåtas vidta för import av vissa varor med ursprung i tredje land och som har övergått till fri omsättning i någon medlemsstat(1) fastställdes vissa kriterier och förfaranden vid tillämpning av artikel 115 i fördraget.
Med hänsyn till erfarenheterna och det åtgärdsprogram gemenskapen har fastställt för genomförandet av den enhetliga marknaden bör beslut 80/47/EEG ändras. I synnerhet bör dess räckvidd utsträckas till alla de fall där det kvarstår skillnader inom de handelspolitiska åtgärder som har vidtagits av medlemsstater i enlighet med fördraget, däribland fall där skillnader inom tulltaxebestämmelser fortfarande tillåts, och vissa av de i beslutet angivna kriterierna och förfarandena bör specificeras. För att inarbeta dessa ändringar bör beslutet omarbetas till en enda rättsakt.
I de fall då en övervakningsåtgärd tillåts måste en importhandling utfärdas automatiskt och utan avgift, inom en given frist och för varje begärd mängd. Om övervakningsåtgärder begärs på grund av att import kan leda till ekonomiska svårigheter för en medlemsstat, bör en sådan risk bedömas mot bakgrund av de störningar i handeln som dittills iakttagits och av storleken av de importmöjligheter gemenskapen har beviljat tredje land i fråga.
Om en medlemsstat begär att få tillämpa skyddsåtgärder, måste fristen för utfärdande av importhandlingar förlängas om den volym som omfattas av ansökningar under prövning når en viss nivå.
De uppgifter och de grunder som medlemsstaterna åberopar till stöd för en begäran om tillstånd för åtgärderna i fråga måste vara av sådan beskaffenhet att kommissionen fullt ut kan bedöma behovet av ett sådant tillstånd.
Om så är nödvändigt bör kommissionen få företa en undersökning för att kontrollera giltigheten av de uppgifter som den har fått till sitt förfogande.
Eftersom de skyddsåtgärder som har beslutats enligt artikel 115 i fördraget, inte bara utgör undantag från bestämmelserna i artiklarna 9 och 30 i fördraget, utan också hindrar upprättandet av en gemensam handelspolitik i enlighet med artikel 113 i fördraget, måste de tolkas och tillämpas strikt. Med hänsyn till detta och till de mål som har fastställts i som har fastställts i Europeiska enhetsakten bör sådana åtgärder bara tillämpas under en begränsad tid och när lägets allvar så kräver.
För att handeln mellan medlemsstaterna inte skall hindras, bör det föreskrivas att medlemsstaterna som regel bara skall begära vissa uppgifter från importören som ett led i uppfyllandet av formaliteterna vid import av en vara från en annan medlemsstat. Vad beträffar kontroll av ursprung skall medlemsstaterna i regel bara begära en enkel ursprungsdeklaration för varan, eftersom importören rimligen kan antas känna till ursprunget.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Räckvidd
Detta beslut gäller för import till en medlemsstat av varor med ursprung i tredje land, som har övergått till fri omsättning inom gemenskapen och inte är underkastade enhetliga importvillkor i medlemsstaterna.
Artikel 2
Övervakning inom gemenskapen
1. När det kan befaras att import till en medlemsstat av en sådan vara som avses i artikel 1 kan leda till ekonomiska svårigheter, får som villkor för import med tidsbegränsat tillstånd från kommissionen, krävas att en importhandling utfärdas.
2. I regel skall kommissionen inte ge sådant tillstånd som avses i punkt 1 om
a) det inte har skett betydande import av den ifrågavarande varan från andra medlemsstater under kalenderåret före det år då ansökan görs,
b) importmöjligheter som gemenskapen har öppnat för varan gentemot det tredje land som är ursprungsland inte överstiger 1 % av de sammanlagda importmöjligheterna som gemenskapen har öppnat gentemot alla tredje länder för vilka liknande regler gäller.
3. Utan att det påverkar tillämpningen av artikel 3, skall importhandlingen utfärdas av medlemsstaten i fråga, för varje begärd kvantitet och utan avgift, inom högst fem arbetsdagar från dagen för importörens ansökan, oberoende av var hans företag är beläget inom gemenskapen.
4. För att erhålla det tillstånd som avses i punkt 1 skall medlemsstaten lämna följande uppgifter i sin ansökan till kommissionen:
a) En beskrivning av varan med närmare uppgifter om dess handelsbeteckning, dess nummer i Gemensamma tulltaxan, dess NIMEXE-nummer och dess ursprungsland.
b) De regler som gäller för direkt import gentemot ursprungslandet och andra tredje länder, däribland i förekommande fall tullregler, importmöjligheternas storlek eller volym samt de ekonomiska överväganden på vilka reglerna är grundade.
c) Den volym eller den mängd av varan som har sitt ursprung
- i tredje landet i fråga, med fördelning på direkt import och varor i fri omsättning,
- i alla tredje länder,
- inom gemenskapen.
d) Risken för ekonomiska svårigheter som åberopas och huruvida de framgår av sådana faktorer som förbrukningen av varan och de marknadsandelar som gäller för inhemsk produktion, för tredje landet i fråga och för alla tredje länder.
De uppgifter som krävs enligt punkterna c och d skall omfatta de två närmast föregående åren och det aktuella året. Om dessa uppgifter inte kan tillhandahållas i tid eller med den noggrannhet som krävs, skall medlemsstatens ansökan innehålla de uppgifter som finns tillgängliga.
5. En medlemsstat som har fått det tillstånd som avses i punkt 1 får av den som ansöker om importhandling bara begära följande uppgifter:
a) Uppgifter som identifierar importören samt avsändaren i den exporterande medlemsstaten.
b) Uppgift om ursprungslandet och den exporterande medlemsstaten.
c) En beskrivning av varan med uppgift om
- dess handelsbeteckning,
- dess nummer i Gemensamma tulltaxan samt dess NIMEXE-nummer.
d) Varans värde och kvantitet i de enheter som vanligen används i handeln.
e) Planerad dag eller planerade dagar för leverans.
f) Uppgifter som styrker att varorna är i fri omsättning. Om varorna ännu inte är i fri omsättning den dag då ansökan om import görs eller om det vid den tidpunkten inte går att styrka att de är i fri omsättning, skall en importhandling utfärdas, men giltigheten begränsas till en månad efter den tidpunkt då den sökande tar emot handlingen.
Artikel 3
Skyddsåtgärder
1. I de fall då import till en medlemsstat av en vara som avses i artikel 1 medför ekonomiska svårigheter får medlemsstaten i fråga vidta skyddsåtgärder efter att ha fått tillstånd från kommissionen, som skall bestämma villkor och närmare regler för sådana åtgärder.
2. Kommissionen skall bevilja tillståndet bara för en begränsad period och bara när lägets allvar så kräver.
3. För att få tillstånd skall medlemsstaten i sin ansökan till kommissionen lämna följande uppgifter utöver de uppgifter som avses i artikel 2.4 a och 2.4 b:
a) Den exporterande medlemsstaten.
b) Den dag då ansökan om importhandling lämnades in.
c) Den faktiska eller tillåtna importvolymen eller importmängden för varan i fråga
- när den har sitt ursprung i tredje landet i fråga, med fördelning på direkt import och import av varor i fri omsättning,
- när den har sitt ursprung i andra tredje länder gentemot vilka den ansökande medlemsstaten til lämpar liknande importregler eller regler med motsvarande verkan,
- med ursprung i alla tredje länder,
- med ursprung i gemenskapen.
d) Där så är möjligt, den volym eller den mängd av varan med ursprung i tredje landet i fråga som återexporteras till andra medlemsstater och till tredje land.
e) De åberopade ekonomiska svårigheterna, vilka framgår av sådana faktorer som produktion, kapacitetsutnyttjande, förbrukning, försäljning, marknadsandelarna för det tredje landet i fråga, för alla tredje länder och för inhemsk produktion, samt priser (dvs. pressade priser eller uteblivna normala prisstegringar), vinster eller förluster, sysselsättning.
f) Om kommissionen begär det, de åtgärder som har vidtagits eller föreslagits för att avhjälpa situationen för den berörda sektorn.
De uppgifter som begärs enligt punkterna c-e skall omfatta de två närmast föregående åren och det aktuella året.
5. I de fall då medlemsstaten finner att den volym eller den sammanlagda mängd som omfattas av ansökningar under prövning avseende import av varan i fråga med ursprung i tredje landet överstiger antingen 5 % av eventuell direkt import från det tredje landet eller 1 % av den sammanlagda importen från länder utanför EEG under den senaste tolvmånadsperiod för vilken statistiska uppgifter finns tillgängliga, skall dock följande gälla:
- Fristen för utfärdande av importhandlingar skall ökas till tio arbetsdagar från den dag då importören lämnade in sin ansökan.
- Medlemsstaten får avslå ansökan om en importhandling om kommissionens beslut tillåter detta.
6. Medlemsstaten skall sända in sin ansökan om tillstånd till skyddsåtgärder med telex eller telefax. En kopia skall samtidigt och på samma sätt sändas till de behöriga myndigheter som för detta syfte har utsetts av de andra medlemsstaterna. Medlemsstaten skall vidare underrätta dem som har ansökt om importhandlingar om att en ansökan om skyddsåtgärder har lämnats in.
7. Kommissionen skall ta ställning till medlemsstatens begäran inom fem arbetsdagar efter mottagandet.
Artikel 4
Ursprungsbevis
1. Som ett led i uppfyllandet av formaliteterna i samband med import av varor som är föremål för övervaknings- eller skyddsåtgärder inom gemenskapen får medlemsstatens behöriga myndigheter anmoda importören att ange ursprunget av de varor som är upptagna i tulldeklarationen eller i ansökan om en importhandling.
Artikel 5
Slutbestämmelser De förfaranden som fastställs genom detta beslut skall gälla när verkan av de handelspolitiska åtgärder som en medlemsstat tillämpar i överensstämmelse med gemenskapens internationella åtaganden äventyras av en störning i handeln med undantag för vad som avses i artiklarna 2.4 d och 3.3 e.
Artikel 6
1. Detta beslut skall tillämpas från och med den 1 oktober 1987.
2. Kommissionens beslut 80/47/EEG skall upphöra att gälla från och med samma dag. Hänvisningar till det upphävda beslutet skall betraktas som hänvisningar till detta beslut.
Artikel 7
Detta beslut riktar sig till medlemsstaterna.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2), och
med beaktande av följande: Direktiv 70/156/EEG(3), senast ändrat genom Anslutningsakten för Spanien och Portugal, fastställde gemenskapens förfarande för typgodkännande av fordon som tillverkas i enlighet med de tekniska krav som specificerats i särdirektiv, och även förteckningen över fordonsdelar och egenskaper som ingår i dessa direktiv.
För att undanröja risken för missförstånd på grund av ordalydelsen i vissa artiklar i nämnda direktiv, är det nödvändigt att införa mindre rättelser.
För att förfarandet för typgodkännande skall kunna tillämpas fullständigt är det nödvändigt att det omfattar såväl komponenter som särskilda tekniska enheter och att varje begrepp definieras noggrant.
För att tillämpa förfarandet för typgodkännande på ett riktigt sätt bör kontroller av produktionens överensstämmelse även avse åtgärder som vidtagits av tillverkaren i syfte att säkerställa att fordon, särskilda tekniska enheter eller komponenter i serietillverkning överensstämmer med den godkända typen.
För att minska antalet dokument som nu cirkulerar mellan medlemsstaterna bör ett typgodkännandeintyg, antingen i enlighet med det tillämpliga särdirektivet eller med förebilden i direktiv 70/156/EEG, anses uppfylla medlemsstaternas normala informationskrav. Medlemsstaterna har dock rätt att begära utförligare tekniska upplysningar.
Ett förtydligande behövs för de administrativa förfaranden som styr förhållandet mellan medlemsstaterna, i det fall en medlemsstat påvisar att ett antal fordon inte överensstämmer med den godkända typen för den medlemsstat som har utfärdat typgodkännandet och att det därför finns skäl att anta att produktionens överensstämmelse inte har kontrollerats i tillräcklig grad.
I de fall där det i särdirektiven föreskrivs att en särskild teknisk enhet måste förses med typgodkännandenummer behöver varje enhet inte nödvändigtvis åtföljas av ett intyg om överensstämmelse. Tillverkaren av en särskild teknisk enhet måste i varje enskilt fall tillhandahålla upplysningar om begränsningar i användningen av enheten och villkoren för dess montering.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 70/156/EEG ändras på följande sätt:
I detta direktiv avses med:
- fordon: dels varje motordrivet fordon avsett att användas på väg, med eller utan karosseri, som har minst fyra hjul och som är konstruerad för en högsta hastighet som överstiger 25 km/tim, dels släpvagnar till dessa fordon, spårbundna fordon, jordbrukstraktorer och lantbruksmaskiner är undantagna,
- särskild teknisk enhet: en anordning för vilken det fastställs krav i ett särdirektiv, som är avsedd att vara en del av ett fordon och som kan vara typgodkänt särskilt men endast i samband med en eller flera, specificerade fordonstyper,
- komponent: en anordning för vilken det fastställs krav i ett särdirektiv, som är avsedd att vara en del av ett fordon och som kan vara typgodkänd oberoende av ett fordon.
Artikel 2
I detta direktiv avses med:
a) nationellt typgodkännande ett administrativt förfarande som benämns:
-"agrément par type"/"typegoedkeuring" i belgisk lagstiftning,
- "standardtypegodkendelse" i dansk lagstiftning,
- "allgemeine Betriebserlaubnis" i tysk lagstiftning,
- "Ýãêñéóç ôýðïõ" i grekisk lagstiftning,
- "homologacion de tipo" i spansk lagstiftning,
- "réception par type" i fransk lagstiftning,
- "type approval" i irländsk lagstiftning,
- "omologazione" eller "approvazione del tipo" i italiensk lagstiftning,
- "agrément" i luxemburgsk lagstiftning,
- "typegoedkeuring" i nederländsk lagstiftning,
- "aprovaço de marca e modelo" i portugisisk lagstiftning,
- "type approval" i brittisk lagstiftning.
b) EEG-typgodkännande avser det förfarande genom vilket en medlemsstat fastställer att en fordonstyp, en särskild teknisk enhet eller komponent, uppfyller de tekniska kraven i särdirektiven och de kontroller som anges i EEG-typgodkännandeintyget. En förebild för detta visas i bilaga 2 och skall, i tillämpliga fall, kompletteras enligt bilagan till typgodkännandeintyget i det berörda direktivet."
2. Artiklarna 4 och 5 skall ersättas med följande:
"Artikel 4
1. Varje medlemsstat skall godkänna alla fordonstyper som uppfyller följande villkor:
a) Fordonstypen måste överensstämma med specifikationerna i det tekniska underlaget.
b) Fordonstypen måste uppfylla de kontrollkrav som anges i den förebild för typgodkännandeintyg som avses i artikel 2 b.
2. En medlemsstat som har beviljat ett typgodkännande skall vidta nödvändiga åtgärder för att, i nödvändig utsträckning och vid behov i samarbete med behöriga myndigheter i andra medlemsstater, kontrollera att tillräckliga åtgärder har gjorts som säkerställer att serietillverkade fordon överensstämmer med den godkända typen.
3. En medlemsstat som har beviljat typgodkännande skall i nödvändig utsträckning och vid behov i samarbete med behöriga myndigheter i andra medlemsstater, vidta nödvändiga åtgärder för att kontrollera att de åtgärder som avses i punkt 2 även fortsättningsvis är tillräckliga och att serietillverkade fordon överensstämmer med den godkända typen. Kontroll av att serietillverkade fordon överensstämmer med den godkända typen skall begränsas till stickprovskontroller, såvida inte annat anges i särdirektiven.
4. Varje medlemsstat skall fylla i alla avsnitt av ett typgodkännandeintyg för varje fordonstyp som den godkänner.
Artikel 5
1. De behöriga myndigheterna i varje medlemsstat skall inom en månad sända en kopia av typgodkännandeintyget för varje fordonstyp som har godkänts eller vägrats godkännande till de behöriga myndigheterna i de andra medlemsstaterna.
2. Medlemsstater har dock rätt att från en medlemsstat som har utfärdat typgodkännandet, eller från tillverkaren eller dennes representant, begära ytterligare sådana upplysningar som anges i de tekniska dokumenten i typgodkännandeintyget.
3. Tillverkaren eller dennes representant i registreringslandet skall för varje fordon som tillverkas i enlighet med den godkända typen utfärda ett intyg om överensstämmelse, för vilket en förebild visas i bilaga 3.
4. Artikel 7.2 skall ersättas med följande:
"2. Ett sådant intyg får dock inte hindra en medlemsstat från att vidta sådana åtgärder mot fordon som inte överensstämmer med den godkända typen.
Ett fordon anses inte överensstämma med den godkända typen om det avviker från uppgifterna i typgodkännandeintyget och/eller det tekniska underlaget förutsatt att dessa avvikelser inte har godkänts under artikel 6.2 eller 6.3 av den medlemsstat som har beviljat typgodkännandet. Ett fordon skall inte anses avvika från den godkända typen om toleranser som anges i särdirektiv inte överskrids."
5. Artikel 8 skall ersättas med följande:
"Artikel 8
1. Om en medlemsstat som har utfärdat EEG-typgodkännandet finner att ett antal fordon med intyg om överensstämmelse inte överensstämmer med den godkända typen, skall den vidta nödvändiga åtgärder för att säkerställa att serietillverkade exemplar överensstämmer med den godkända typen. De behöriga myndigheterna i denna stat skall upplysa motsvarande myndigheter i de andra medlemsstaterna om vidtagna åtgärder vilket, om så är påkallat, kan leda till att EEG-typgodkännandet återkallas. 2. Om en medlemsstat påvisar att ett antal fordon med intyg om överensstämmelse inte överensstämmer med den godkända typen kan denna stat begära att medlemsstaten som har utfärdat EEG-typgodkännandet visar att serietillverkade fordon överensstämmer med den godkända typen. Medlemsstaten som utfärdade EEG-typgodkännandet skall, inom sex månader räknat från dagen för en begäran, kontrollera att produktionen är i överensstämmelse med den godkända typen. Kontrollen kan, om så bedöms nödvändigt, utföras i samarbete med den medlemsstat som begärde att en sådan kontroll skulle utföras.
Om bristande överensstämmelse konstateras skall de behöriga myndigheterna i den medlemsstat som utfärdade typgodkännandet vidta de åtgärder som beskrivs under punkt 1.
3. De behöriga myndigheterna i medlemsstaterna skall inom en månad upplysa varandra om varje återkallat EEG-typgodkännande, och orsakerna till en sådan åtgärd.
4. Om medlemsstaten som beviljade EEG-typgodkännandet ifrågasätter den påpekade avvikelsen, skall de berörda medlemsstaterna bemöda sig att bilägga tvisten.
Kommissionen skall hållas informerad och, den skall vid behov, hålla erforderliga överläggningar i syfte att nå en överenskommelse."
6. Artikel 9a skall ändras enligt följande:
"Artikel 9a
1. EEG-typgodkännande kan, när detta uttryckligen föreskrivs i särdirektiven, även utfärdas för typer av system eller fordonsdelar som utgör en särskild teknisk enhet och för komponenter i överensstämmelse med artiklarna 3 till 9 och 14.
2. När den särskilda tekniska enheten eller komponenten som skall godkännas fyller sin funktion eller erbjuder en särskild egenskap endast tillsammans med andra fordonskomponenter och dess överensstämmelse med ett eller flera krav av denna anledning endast kan visas när den tekniska enheten eller komponenten som skall godkännas används tillsammans med andra fordonskomponenter, antingen på verkliga eller simulerade, måste omfattningen av EEG-typgodkännandet för den tekniska enheten eller komponenten begränsas i motsvarande grad. EEG-typgodkännandeintyget för en särskild teknisk enhet eller komponent skall i detta fall innehålla uppgifter om begränsning av dess användning och skall utvisa varje villkor för dess montering. Efterlevnaden av dessa begränsningar och villkor skall kontrolleras då fordonet EEG-typgodkänns.
3. Emellertid skall innehavaren av EEG-typgodkännande för en särskild teknisk enhet eller en komponent, vilka beviljats i enlighet med denna artikel, utfärda intyget som beskrivs i artikel 5.3 och märka varje enhet eller komponent som tillverkats i enlighet med den godkända typen med handelsbeteckning eller varumärke, typen och, om så anges i särdirektivet, typgodkännandets nummer. I det senare fallet medför detta ingen skyldighet att utfärda intyget som föreskrivs i artikel 5.3.
4. Innehavaren av ett EEG-typgodkännandeintyg, vilket, i enlighet med bestämmelserna i punkt 2, innehåller uppgifter om begränsningar i fråga om användning, skall för varje tillverkad enhet eller komponent tillhandahålla detaljerade upplysningar om dessa begränsningar och varje villkor för montering."
7. Det tredje indraget i artikel 10.1 skall ersättas med följande:
"- vid ansökan från en tillverkare eller dennes representant och inlämnandet av de upplysningar som krävs enligt särdirektivet, skall den berörda medlemsstaten färdigställa intyget om typgodkännande i enlighet med det tillgängliga särdirektivet. En kopia av intyget skall sändas till sökanden. Andra medlemsstater skall, för fordon av samma typ, acceptera denna kopia som bevis på att nödvändiga provningar har utförts."
Artikel 2
De dokument som anges i bilagan till detta direktiv skall anses likvärdiga med de typgodkännandeintyg, vilka nämns i det tredje indraget i artikel 10.1 i direktiv 70/156/EEG.
Artikel 3
1. Medlemsstaterna skall till den 1 oktober 1988 sätta i kraft de författningar som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
2. Medlemsstaterna skall se till att kommissionen tillställs texten till de viktigaste bestämmelser i den nationella lagstiftningen som de antar inom det område som omfattas av detta direktiv.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av rådets direktiv 79/117/EEG av den 21 december 1978 om förbud mot att växtskyddsprodukter som innehåller vissa verksamma ämnen släpps ut på marknaden och används(), särskilt artikel 6 i detta, senast ändrat genom direktiv 87/181/EEG(), och
med beaktande av följande: Vetenskapliga och tekniska framsteg medför att vissa ändringar måste göras i bilagan till direktiv 79/117/EEG.
Det finns skäl att upphäva vissa av de tillfälliga undantagen från förbuden i direktivet, eftersom mindre farliga behandlingsmetoder nu finns att tillgå.
Samtliga medlemsstater har meddelat kommissionen att de inte kommer att eller inte längre avser att utnyttja dessa undantag.
De åtgärder som föreskrivs genom detta direktiv är förenliga med yttrandet från Ständiga kommittén för växtskydd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
b) under 5, "Alkoxyalkyl- och arylkvicksilverföreningar", skall texten i andra kolumnen ersättas med: "Behandling av utsäde till spannmål och betor".
2. I del B, "Svårnedbrytbara organiska klorföreningar", under 1, "Aldrin", skall texten till b i andra kolumnen ändras genom att orden "Irland och" utgår.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(1), senast ändrad genom förordning nr (EEG) 1454/86(2), särskilt artikel 5.4 i denna,
med beaktande av kommissionens förslag, och
med beaktande av följande: I artikel 13 i förordning (EEG) nr 2261/84(3), senast ändrad genom förordning (EEG) nr 3788/85(4), föreskrivs att tillfälligt godkännande får beviljas för fabriker som lämnar in en ansökan om godkännande under regleringssåren 1984/85 och 1985/86. Erfarenheten har visat att de berörda medlemsstaterna inte är i stånd att genomföra de kontroller som behövs inom den fastställda tiden. Dessa tider bör därför förlängas.
Innan medlemsstaterna har möjlighet att definitivt godkänna en fabrik skall de utföra vissa kontroller. För att göra det möjligt för fabrikerna att börja sin verksamhet bör bestämmelser införas för beviljande av ett tillfälligt tillstånd under en begränsad tid, så snart som ansökan har lämnats in.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Första stycket i artikel 13.3 i förordning (EEG) nr 2261/84 skall ersättas med följande:
"Tillfälligt tillstånd får beviljas för en fabrik som börjar sin verksamhet enligt det program för produktionsstöd som fastställs i denna förordning. Tillståndet skall beviljas så snart en ansökan om godkännande har lämnats in enligt de i punkt 1 angivna villkoren. Giltighetstiden för det tillfälliga tillståndet får inte vara längre än till slutet av det regleringsår då det beviljades. Giltighetstiden för tillfälliga tillstånd som beviljades under regleringsåren 1984/85, 1985/86 och 1986/87 skall upphöra vid utgången av regleringsåret 1986/87."
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
RÅDETS FÖRORDNING (EEG) nr 678/87 av den 26 januari 1987 om tillämpningen av systemet med ursprungscertifikat som föreskrivs enligt Internationella kaffeavtalet 1983 när kvoterna är tillfälligt upphävda
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 113 i detta,
med beaktande av rådets förordning (EEG) nr 288/82 av den 5 februari 1982 om gemenskapsregler för import(1), senast ändrad genom förordning (EEG) nr 899/83(2), särskilt artikel 16.1 b i denna,
med beaktande av kommissionens förslag, och
med beaktande av följande: Enligt beslut 83/539/EEG(3) har gemenskapen provisoriskt tillämpat Internationella kaffeavtalet 1983 sedan denna provisoriskt trädde i kraft den 1 oktober 1983.
Förordning (EEG) nr 3761/83(4) införde det system med ursprungsintyg som föreskrivs i Internationella kaffeavtalet 1983 när kvoterna tillämpas.
Lämpliga åtgärder skall vidtas för att genomföra det nya systemet med intyg inom gemenskapen och för att se till att det tillämpas utan att några importörer i gemenskapen missgynnas.
För att säkerställa en effektiv förvaltning av systemet och för att klargöra frågan under vilken tid denna förordning faktiskt kommer att gälla, och för att uppfylla regel 11 i bilagan till denna förordning och till regel 47 i bilagan till förordning (EEG) nr 3761/83, bör åtgärder vidtas för kommissionen, enligt de beslut som fattats av de behöriga organen i Internationella kaffeorganisationen och vid den tid då kvoterna är tillfälligt upphävda eller återinförs, för att ange den dag då åtgärderna i fråga skall bli tillämpliga eller upphöra att vara tillämpliga.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Export från gemenskapen av kaffe och extrakt, essenser eller koncentrat av kaffe enligt undernummer 09.01 A och 21.02 A i Gemensamma tulltaxan skall inte vara beroende av inlämnande av de intyg som föreskrivs i avtalet.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av rådets förordning (EEG) nr 170/83 av den 25 januari 1983 om ett gemenskapssystem för bevarande och förvaltning av fiskeresurserna(),
med beaktande av rådets förordning (EEG) nr 3094/86 av den 7 oktober 1986 om vissa tekniska åtgärder för bevarande av fiskeresurserna(), ändrad genom förordning (EEG) nr 4026/86(), särskilt artikel 15 i denna, och med beaktande av följande:
I artikel 6.3 i kommissionens förordning (EEG) nr 3440/84() fastställs att det är tillåtet att sätta fast en förstärkande nätkasse på trålar, danska snurrevadar och liknande nätredskap under förutsättning att dess maskstorlek är minst 80 millimeter.
Om en förstärkande nätkasse med denna maskstorlek används på nätredskap med en maskstorlek som är mindre än 40 millimeter har det visat sig att det bildas nätfickor, som leder till skador på fångsten beroende på tekniska problem med att få ut denna ur lyftet, vilket leder till att lyftet slits ut och rivs sönder.
Om en förstärkande nätkasse med mindre maskstorlek användes skulle dessa problem kunna undvikas utan negativ inverkan på fiskebeståndet.
Definitionerna på nätkategorierna i artiklarna 5 och 6 i förordning (EEG) nr 3440/84 behöver därför ändras.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fiskeresurser.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 3440/84 ändras på följande sätt:
1. Artikel 5.5 skall ersättas med följande:
"5. Det är förbjudet att använda ett övre slitskydd tillsammans med förstärkande nätkassar, med undantag för trålar med en maskstorlek på 60 mm eller mindre."
2. Artikel 6 skall ändras enligt följande:
- Punkt 2 skall ersättas med följande:
"2. Det är bara tillåtet att använda en förstärkande nätkasse åt gången, med undantag för trålar med en maskstorlek på högst 60 mm, för vilka två förstärkande nätkassar får användas."
- Punkt 3 skall ersättas med följande:
"3. Maskstorleken skall vara minst dubbelt så stor som lyftets. Om en andra förstärkande nätkasse används skall den ha en maskstorlek på minst 120 mm."
- Punkt 6 skall ersättas med följande:
"6. En förstärkande nätkasse som är fastsatt på en trål med en maskstorlek på över 60 mm får sträcka sig högst två meter framför den bakre lyftstoppen."
- Punkt 7 skall ersättas med följande:
"7. Trots punkt 1 får en förstärkande nätkasse som är mindre än lyftet sättas fast på redskap med en maskstorlek på högst 60 mm."
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EEG) nr 4155/87 av den 22 december 1987 om ändring av vissa förordningar om tillämpningen av den gemensamma organisationen av marknaden för ägg till följd av införandet av Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (), ändrad genom förordning (EEG) nr 3985/87 (), särskilt artikel 15.1 andra stycket i denna, och med beaktande av följande: I enlighet med artikel 15.1 andra stycket i förordning (EEG) nr 2658/87 skall kommissionen göra anpassningar av teknisk art av gemenskapens rättsakter som hänvisar till tulltaxe- eller statistiknomenklaturen. Rådets förordning (EEG) nr 2771/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för ägg () har ändrats genom kommissionens förordning (EEG) nr 4000/87 (), varvid varubeskrivningarna och de tulltaxenummer som anges i dessa anpassades i enlighet med Kombinerade nomenklaturen. Många andra förordningar om äggsektorn måste bli föremål för en teknisk anpassning varvid hänsyn skall tas till nya Kombinerade nomenklaturen som är baserad på systemet för harmoniserad varubeskrivning- och kodifiering som skall ersätta konventionen av den 15 december 1950 om nomenklaturen för klassificering av handelsvaror i tulltaxor. På grund av antalet och innehållet i de texter där en anpassning är nödvändig, bör alla förordningar som skall anpassas samlas i en ändringsförordning. I samband med denna anpassning av kommissionens förordning 164/67/EEG () bör vissa faktorer som används vid beräkningen av slusspriserna och som i nämnda förordning fortfarande anges i beräkningsenheter, uttryckas i ecu med användning av den koefficient på 1,208 953 som avses i artikel 13 i rådets förordning (EEG) nr 1676/85 (), senast ändrad genom förordning (EEG) nr 1636/87 (). HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 1 i kommissionens förordning nr 54/65/EEG () av den 7 april 1965 om icke-fastställande av en tilläggsavgift för polska ägg skall ersättas med följande: "Artikel 1 I enlighet med artikel 8.2 i förordning (EEG) nr 2771/75 skall de importavgifter som skall betalas vid import av fjäderfäägg med skal (undernummer 0407 00 i Kombinerade nomenklaturen) som har sitt ursprung i och kommer från Polen, inte höjas med en tilläggsavgift."
Artikel 2
Artikel 1 i kommissionens förordning nr 183/66/EEG av den 18 november 1966 om icke-fastställande av en tilläggsavgift för sydafrikanska ägg () skall ersättas med följande: "Artikel 1 I enlighet med artikel 8.2 i förordning (EEG) nr 2771/75 skall de importavgifter som fastställts i enlighet med artikel 3 i samma förordning inte höjas med en tilläggsavgift i samband med import av ägg med skal (undernummer 0407 00 i Kombinerade nomenklaturen) som har sitt ursprung i och kommer från Sydafrika."
Artikel 3
Bilagan till kommissionens förordning nr 164/67/EEG av den 26 juni 1967 om fastställande av faktorerna för beräkning av importavgifter och slusspriser för härledda äggprodukter, senast ändrad genom förordning (EEG) nr 1775/74 (), skall ersättas med bilaga 1 till den här förordningen.
Artikel 4
Artikel 1 i kommissionens förordning nr 765/67/EEG av den 26 oktober 1967 om icke-fastställande av en tilläggsavgift för australiska ägg () skall ersättas med följande: "Artikel 1 Importavgifter som fastställts i enlighet med artikel 3 i förordning (EEG) nr 2771/75 skall inte höjas med en tilläggsavgift när det gäller import av färska, konserverade, kokta eller på annat sätt värmebehandlade fjäderfäägg med skal, undantaget kläckägg som omfattas av undernummer 0407 00 30 i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Australien."
Artikel 5
1. Artikel 1 skall ersättas med följande: "Artikel 1 Importavgifter som fastställs i enlighet med artikel 3 i förordning (EEG) nr 2771/75 skall inte höjas med en tilläggsavgift i samband med import av produkter som omfattas av följande nummer i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Österrike: >Plats för tabell>
2. Artikel 2 skall ersättas med följande: "Artikel 2 Importförändringar som fastställts i enlighet med artikel 2 i förordning (EEG) nr 2783/75 avseende produkter som omfattas av följande undernummer i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Österrike, skall inte höjas med en tilläggsavgift: () EGT nr L 186, 1.7.1974, s. 14. () EGT nr 260, 27.10.1967, s. 24. () EGT nr L 130, 31.5.1969, s. 4. >Plats för tabell>
Artikel 6
Artikel 1 i kommissionens förordning (EEG) nr 59/70 av den 14 januari 1970 om ickefastställande av tilläggsavgifter för ägg med skal som importeras från Rumänien () skall ersättas med följande: "Artikel 1 Importavgifter som fastställts i enlighet med artikel 3 i förordning (EEG) nr 2771/75 skall inte höjas med en tilläggsavgift i samband med import av fjäderfäägg med skal, färska eller konserverade, undantaget kläckägg, som omfattas av undernummer 0407 00 30 i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Rumänien."
Artikel 7
Bilagorna 1 och 2 till rådets förordning (EEG) nr 2773/75 av den 29 oktober 1975 om fastställande av bestämmelser för beräkning av importavgiften och slusspriset för ägg (), senast ändrad genom förordning (EEG) nr 3232/86 (), skall ersättas med bilaga 2 och 3 till denna förordning.
Artikel 8
Denna förordning träder i kraft den 1 januari 1988.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater. ()()()
KOMMISSIONENS BESLUT av den 28 oktober 1988 om upprättande av en förteckning över produkter som avses i artikel 3.1 andra stycket i rådets förordning (EEG) nr 1898/87 (88/566/EEG)
med beaktande av rådets förordning (EEG) nr 1898/87 av den 2 juli 1987 om skydd för beteckningar som används vid saluförande av mjölk och mjölkprodukter(1), senast ändrad genom förordning (EEG) nr 222/88(2), särskilt artikel 4.2 b i denna, och
med beaktande av följande: Genom förordning (EEG) nr 1898/87 fastställs principen att beteckningarna mjölk och mjölkprodukter inte får användas för andra produkter än de som upptas i förordningens artikel 2. Ett undantag från denna princip är beteckningen på produkter vars beskaffenhet är känd genom traditionellt bruk eller beteckningar som uppenbarligen används för att beskriva en karakteristisk egenskap hos produkten.
Artikel 1 De produkter inom gemenskapens territorium som motsvarar de produkter som avses i artikel 3.1 andra stycket i förordning (EEG) nr 1898/87 upptas i förteckningen i bilagan.
Artikel 2 Detta beslut riktar sig till medlemsstaterna.
med beaktande av rådets direktiv 71/127/EEG av den 1 mars 1971 om tillnärmning av medlemsstaternas lagstiftning om backspeglar för motorfordon(1), i dess lydelse enligt kommissionens direktiv 86/562/EEG(2), särskilt artikel 9 i detta, och
med beaktande av följande: Med hänsyn till vunna erfarenheter och teknikens nuvarande utvecklingsnivå är det nu möjligt att skärpa vissa krav i direktiv 71/127/EEG i syfte att förbättra trafiksäkerheten.
För fordon i kategori N2 med en massa över 7,5 ton och andra fordon än dragfordon för påhängsvagn i kategori N3 har nuvarande krav visat sig otillräckliga vad avser det yttre siktfältet längs fordonets sida och bakåt. För att råda bot på denna brist är det nödvändigt att möjliggöra montering av en extra backspegel av s.k. vidvinkeltyp.
För fordon i kategori N2 med en massa över 7,5 ton har nuvarande krav även visat sig otillräckliga vad avser siktfältet längs den sida av förarhytten som är längst bort från föraren. För att råda bot på denna brist är det nödvändigt att möjliggöra montering av en närzonsbackpegel.
De i detta direktiv fastställda åtgärderna har tillstyrkts av Kommittén för anpassning till teknisk utveckling av direktiv om avskaffande av tekniska handelshinder inom motorfordonssektorn.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagorna 2 och 3 till direktiv 71/127/EEG ändras härigenom i enlighet med bilagan till detta direktiv.
Artikel 2
1. Från och med den 1 januari 1989 får medlemsstaterna inte, av skäl som hänför sig till backspeglar
- vare sig vägra att bevilja EEG-typgodkännande eller att utfärda dokumentet enligt artikel 10.1. tredje strecksatsen i rådets direktiv 70/156/EEG(3), eller att bevilja nationellt typgodkännande,
- eller förbjuda att fordon tas i bruk,
om backspeglarna på denna fordonstyp eller dessa fordonstyper överensstämmer med bestämmelserna i detta direktiv.
2. Från och med den 1 oktober 1990 gäller följande:
- Medlemsstaterna får inte längre utfärda dokumentet enligt artikel 10.1 tredje strecksatsen i direktiv 70/156/EEG för en typ av fordon, vars backspeglar inte överensstämmer med bestämmelserna i det här direktivet.
- Medlemsstaterna får vägra nationellt typgodkännande för en fordonstyp, vars backspeglar inte överensstämmer med bestämmelserna i detta direktiv.
- De får förbjuda att fordon, vars backspeglar inte överensstämmer med bestämmelserna i detta direktiv tas i bruk.
Artikel 3
Medlemsstaterna skall senast den 1 januari 1989 sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(),
Direktiv 83/181/EEG bestämmer inte bara räckvidden av artikel 14.1 d i direktiv 77/388/EEG(), senast ändrat genom direktiv 84/386/EEG(), utan syftar även till upprättandet av gemenskapsregler för momsbefrielse vid slutlig införsel av varor som går utöver räckvidden av den nämnda artikeln. Dessa regler bör ändras eller kompletteras på ett sådant sätt att de åstadkommer en mer enhetlig tillämpning av detta på gemenskapsnivå.
För den juridiska klarhetens skull bör ordalydelsen av artikel 11.2 i direktiv 83/181/EEG preciseras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 83/181/EEG ändras på följande sätt:
1. Artikel 11.2 skall ersättas med följande:
"2. Befrielse skall också beviljas när det gäller sedvanliga bröllopsgåvor som ges till en person som uppfyller de villkor som fastställs i punkt 1 av personer som har sin normala bosättningsort i ett land utanför gemenskapen. Befrielsen skall tillämpas på gåvor med ett värde av högst 200 ecu per styck. Medlemsstater får dock bevilja befrielse för mer än 200 ecu, om värdet av varje skattebefriad gåva inte överstiger 1 000 ecu."
2. Artikel 22 skall ersättas med följande:
"Artikel 22
3. I artikel 35.1 b andra strecksatsen skall orden "artikel 60.1 b" ersättas med "artikel 60".
4. Följande kapitel införs efter artikel 38:
"Kapitel IIa
Referenssubstanser för kvalitetskontroll av läkemedel
Artikel 38 a
Sändningar som innehåller varuprov av referenssubstanser som godkänts av Världshälsoorganisationen för kvalitetskontroll av material som används vid tillverkning av läkemedel och som är adresserade till mottagare som är bemyndigade av medlemsstaternas behöriga myndigheter att ta emot sådana försändelser utan att erlägga skatt skall vara skattebefriade vid införsel."
5. Följande tillfogas till artikel 56:
"d) Priser, troféer och souvenirer av symbolisk natur och med begränsat värde, avsedda för gratisutdelning till personer som normalt är bosatta i ett annat land än införsellandet vid affärskonferenser eller liknande internationella evenemang, och vars beskaffenhet, värde per styck eller övriga kännetecken inte är sådana att de skulle kunna vara avsedda för kommersiella ändamål."
6. Artiklarna 62 och 63 skall ersättas med följande:
"Artikel 62
Med förbehåll för vad som föreskrivs i artikel 63 skall tryckt reklammaterial såsom kataloger, prislistor, bruksanvisningar eller broschyrer vara skattebefriade vid införsel, om de hänför sig till:
a) varor som är till salu eller uthyrning av en person som är etablerad utanför införselmedlemsstaten, eller
b) tjänster som erbjuds av en person som är etablerad i en annan medlemsstat, eller
c) transport-, handels-, försäkrings- eller banktjänster som erbjuds av en person som är etablerad i ett tredje land.
Artikel 63
Den befrielse som avses i artikel 62 skall begränsas till reklamtrycksaker som uppfyller följande villkor:
a) Trycksakerna måste tydligt utvisa namnet på det företag som producerar, säljer eller hyr ut de varor eller som erbjuder de tjänster till vilka de hänför sig.
b) Varje försändelse får innehålla högst ett dokument eller ett enda exemplar av varje dokument om det består av flera dokument. Försändelser innefattande flera exemplar av samma dokument får emellertid beviljas befrielse, om deras sammanlagda bruttovikt inte överstiger ett kilogram.
c) Trycksakerna får inte vara skickade som gruppförsändelser från samma avsändare till samma mottagare.
Villkoren i punkterna b och c skall dock inte tillämpas på trycksaker som avser antingen varor till salu eller uthyrning eller tjänster som erbjuds av en person som är etablerad i en annan medlemsstat, om trycksakerna har införts och kommer att distribueras gratis."
7. Följande tillfogas till artikel 79:
"s) Införsel av officiella publikationer som utgör språkrör för utförsellandet, internationella institutioner, regionala eller lokala myndigheter eller offentligrättsliga organ, som är etablerade i utförsellandet liksom av trycksaker som distribueras inför val till Europaparlamentet eller nationella val i det land från vilket trycksakerna härrör av utländska politiska organisationer som är officiellt erkända i medlemsstaterna, försåvitt publikationerna och trycksakerna har beskattats i utförsellandet och inte åtnjutit restitution av skatt vid utförsel."
8. Titeln på kapitel VI skall ersättas med följande:
"Bränslen och smörjmedel som finns i motorfordon och specialcontainrar"
1. Om inte annat sägs i artikel 83 85 skall följande varor vara skattebefriade vid införsel:
- specialcontainrar,
b) bränsle som finns i reservdunkar som fraktas av privata motorfordon och motorcyklar, dock högst 10 liter per fordon, med förbehåll för nationella bestämmelser om innehav och transport av bränsle.
2. I punkt 1 används nedan angivna beteckningar med de betydelser som här anges:
a) kommersiella motorfordon: motordrivna vägfordon (även traktor med släpvagn) som genom sin konstruktionstyp och utrustning är utformade för och ägnade att transportera, mot eller utan betalning: - mer än nio personer inräknat föraren,
- varor,
eller vägfordon för annat särskilt ändamål än transport.
b) privata motorfordon: motorfordon som inte omfattas av definitionen i punkt a.
- tankar som av tillverkaren är fast monterade i alla containrar av samma typ som containern i fråga och vars fasta installation gör det möjligt att använda bränslet direkt för att under transporten driva kylsystem och övriga system som specialcontainrar är utrustade med.
d) specialcontainer: container som är försedd med en särskilt utformad anordning för kylsystem, syrsättningssystem, system för termisk isolering eller andra system."
10. Första punkten i artikel 83 ändras på följande sätt:
- I inledningen införs orden "och specialcontainrar" efter orden "kommersiella motorfordon".
- Efter punkt b tillfogas följande:
"c) till 200 liter per specialcontainer och resa."
12. Följande tillfogas till artikel 91:
"c) skattebefrielser i samband med överenskommelser som med hänsyn till principen om reciprocitet ingås med icke-medlemsländer som är avtalsslutande parter till konventionen om internationell civil luftfart (Chicago 1944) i syfte att genomföra rekommenderade praxis enligt 4.42 och 4.44 i bilaga 9 till konventionen (åttonde upplagan, juli 1980)."
Artikel 2
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta direktiv senast den 1 januari 1989. De skall genast underrätta kommissionen om detta.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av rådets förordning (EEG) nr 3878/87 av den 18 december 1987 om produktionsstöd för vissa rissorter(1), senast ändrad genom förordning (EEG) nr 1424/88(2), särskilt artikel 2.3 i denna, och med beaktande av följande:
I artikel 2.1 i förordning (EEG) nr 3878/87 fastställs vilka morfologiska kännetecken rissorterna skall ha för att berättiga till produktionsstöd. I punkt 2 i samma artikel föreskrivs att från och med regleringsåret 1988/89 skall ingen sort berättiga till produktionsstöd som inte också har vissa kvalitativa kännetecken med avseende på klibbighet, konsistens och amylosinnehåll.
Dessa kvalitativa kännetecken bör motsvara de egenskaper som konstateras för sorter som importeras från områden där indicaris traditionellt odlas.
De analysmetoder som skall användas när dessa morfologiska och kvalitativa kännetecknen fastställs, bör närmare anges.
Förfarandet vid ändring av den sortlista som anges i bilaga B till förordning (EEG) nr 3878/87 bör inbegripa årliga kontroller som omfattar provtagning som gör det möjligt att genomföra de nödvändiga sortanalyserna.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Från och med regleringsåret 1988/89 skall endast de rissorter förtecknas i bilaga B till förordning (EEG) nr 3878/87 som har de morfologiska kännetecken som anges i artikel 2.1 i förordningen och följande kvalitativa kännetecken:
- En klibbighet på högst 2,50 gcm.
- En konsistens på minst 0,85 kg/cm².
- Ett amylosinnehåll på minst 21 %.
1. De medlemsstater som vill få en rissort som berättigar till stöd införd i bilaga B till förordning (EEG) nr 3878/87, skall senast den 31 juli varje år till kommissionen överlämna en ansökan där sortens namn anges samt dess inskrivningsreferenser i den nationella sortlistan över jordbruksgrödor.
Artikel 3
1. Det laboratorium som ansvarar för bearbetningen av riset, skall efter att ha genomfört grobarhetsprov och bearbetat riset, översända prover märkta med en kod till samtliga laboratorier som förtecknas i bilaga 2 samt översända ett förseglat meddelande som möjliggör avkodning av proverna till kommissionens tjänstemän.
2. Varje prov som sänds in till laboratorierna för analys skall bestå av minst 100 g råris och minst 750 g helt slipat ris. Proven skall endast bestå av hela riskorn, dock skall hela men kritaktiga korn avlägsnas från prov av helt slipat ris.
Artikel 4
1. Kommissionens personal skall bestämma de aktuella sorternas kännetecken på grundval av det aritmetiska medelvärdet av analysresultaten, sedan det högsta och det lägsta värdet uteslutits.
2. Om en och samma sort är föremål för två eller flera ansökningar, skall dess kännetecken bestämmas som medelvärdet av provresultaten enligt punkt 1.
3. Kommissionens tjänstemän skall före den 31 mars varje år meddela medlemsstaterna om analysresultaten.
Artikel 5
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av rådets förordning (EEG) nr 2658/87(1) av den 23 juli 1978, om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan, senast ändrad genom förordning (EEG) nr 1315/88(2), särskilt artikel 9, och
med beaktande av följande: För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser angående klassificering av de varor som anges i bilagan till den här förordningen.
Förordning (EEG) nr 2658/87 fastställer de allmänna bestämmelserna för tolkningen av Kombinerade nomenklaturen och dessa bestämmelser gäller också varje annan nomenklatur som helt eller delvis grundar sig på denna eller som lägger ytterligare underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser med tanke på tillämpningen av tulltaxebestämmelser eller andra bestämmelser som rör varuhandeln.
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt de tillämpliga KN-nummer som anges i kolumn 2 av de skäl som anges i kolumn 3.
Nomenklaturkommittén har inte yttrat sig över förslaget inom den tid som ordföranden bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i tabellen i bilagan klassificeras nu inom Kombinerade nomenklaturen enligt de tillämpliga KN-nummer som anges i kolumn 2 i denna tabell.
Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2), och
med beaktande av följande: Enligt artikel 1.1 i förordning (EEG) nr 2262/84(3), senast ändrad genom förordning (EEG) nr 3462/87(4), skall de producerande medlemsstaterna upprätta organ som skall utföra vissa kontroller och uppgifter i samband med programmet för produktionsstöd för olivolja. Enligt artikel 1.5 i den förordningen skall rådet före den 1 januari 1989 fastställa metoden för finansiering av organens utgifter från och med regleringsåret 1989/90.
Med hänsyn till den viktiga roll som dessa organ kan spela för att säkerställa att avtalen om produktionsstöd tillämpas på ett korrekt och enhetligt sätt, bör en metod föreskrivas för finansiering av deras faktiska utgifter som gör det möjligt för dem att ha en smidig och effektiv verksamhet inom ramen för en självständig administration som föreskrivs i dessa bestämmelser. Det syftet kan uppnås genom en metod som förenar gemenskapsfinansiering med finansiering av medlemsstaten.
Organen i de fyra producerande medlemsstaterna befinner sig inte i samma läge. På grund av administrativa och juridiska svårigheter har upprättandet av organen och organens verksamhet försenats i vissa medlemsstater. Dessa medlemsstater utnyttjade inte i tillräcklig grad de högsta belopp som var reserverade för dem under inledningsfasen, när utgifterna helt kunde debiteras gemenskapen. Den tid som denna fas omfattar bör därför förlängas med ett år utan höjning av de högsta belopp som redan är tilldelade enligt nuvarande bestämmelser.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 1.5 i förordning (EEG) nr 2262/84 skall ersättas med följande:
"5. Under en tid av fem år från och med den 1 november 1984 skall följande procentsatser av organets faktiska utgifter debiteras de europeiska gemenskapernas allmänna budget:
- För Italien 100 % för de första tre åren upp till högst 14 miljoner ecu och 50 % för det fjärde och femte året,
- För Grekland 100 % upp till högst 7 miljoner ecu.
Under en tid av tre år från och med den 1 november 1989 skall 50 % av de faktiska utgifterna för organen i Italien och Grekland belasta de europeiska gemenskapernas allmänna budget.
För Spanien och Portugal skall 100 % av organets faktiska utgifter under tiden från den 1 mars 1986 till den 31 oktober 1990 täckas av de europeiska gemenskapernas allmänna budget upp till högst 9 300 000 ecu för Spanien och 4 700 000 ecu för Portugal. Under tiden från den 1:a november 1990 till den 31 oktober 1992 skall 50 % av de ifrågavarande utgifterna täckas av denna budget.
Medlemsstaterna får, enligt villkor som skall bestämmas i enlighet med det förfarande som anges i artikel 38 i förordning nr 136/66/EEG, täcka en del av de utgifter som de själva skall bära genom avdrag från det beviljade gemenskapsstödet för olivolja.
Rådet skall med kvalificerad majoritet på förslag från kommissionen senast den 1 januari 1992 fastställa metoden för finansiering av utgifterna i fråga från och med regleringsåret 1992/93."
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
RÅDETS DIREKTIV av den 12 juni 1989 om åtgärder för att främja förbättringar av arbetstagarnas säkerhet och hälsa i arbetet (89/391/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 118a i detta,
med beaktande av kommissionens förslag(1), utarbetat efter samråd med Rådgivande kommittén för arbetarskyddsfrågor,
i samarbete med Europaparlamentet(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Enligt artikel 118a i fördraget skall rådet genom direktiv fastställa minimikrav i syfte att främja förbättringar, framför allt på arbetsmiljöområdet, för att trygga en högre skyddsnivå för arbetstagarnas säkerhet och hälsa.
Direktiv enligt artikel 118a i fördraget får inte medföra sådana administrativa, ekonomiska och rättsliga hinder, som skulle kunna hämma bildandet och utvecklingen av små och medelstora företag.
Kommissionens meddelande om dess program arbetarskyddsfrågor(4) förutsätter att direktiv antas i syfte att säkerställa arbetstagarnas säkerhet och hälsa.
Rådet uppmärksammade i sin resolution av den 21 december 1987 om arbetarskyddsfrågor(5) att kommissionen avsåg att inom en snar framtid föreslå rådet ett direktiv om organisationen av verksamheten för arbetstagarnas säkerhet och hälsa på arbetsplatsen.
Europaparlamentet antog i februari 1988 fyra resolutioner i anslutning till debatten om den inre marknaden och arbetarskydd; i dessa resolutioner anmodas kommissionen uttryckligen att utarbeta ett ramdirektiv, som skall ligga till grund för särdirektiv, vilka skall omfatta alla risker förknippade med säkerhet och hälsa på arbetsplatsen.
Det åligger medlemsstaterna att inom sina territorier verka för förbättringar av arbetstagarnas säkerhet och hälsa; åtgärder, som vidtas för att skydda arbetstagarnas säkerhet och hälsa i arbetet bidrar även, i vissa fall, till att bibehålla hälsan och möjligen säkerheten hos personer i arbetstagarens hushåll.
Medlemsstaternas arbetarskyddslagstiftning varierar avsevärt och behöver förbättras; nationella bestämmelser, som ofta innehåller tekniska föreskrifter och/eller vägledande normer, kan leda till skilda skyddsnivåer och möjliggöra konkurrens på bekostnad av säkerhet och hälsa.
Antalet arbetsolycksfall och arbetssjukdomar är alltjämt för högt; förebyggande åtgärder måste införas eller förbättras utan dröjsmål för att trygga arbetstagarnas säkerhet och hälsa och säkra en högre skyddsnivå.
För att säkerställa en förbättrad skyddsnivå måste arbetstagarna och/eller deras representanter informeras om de risker som föreligger för deras säkerhet och hälsa och om de åtgärder, som krävs för att minska eller eliminera dessa risker; de måste ha förutsättningar att medverka till att tillräckliga skyddsåtgärder vidtas genom avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis.
Information, dialog och avvägd medverkan i frågor som rör säkerhet och hälsa i arbetet måste utvecklas mellan arbetsgivare och arbetstagare och/eller deras representanter med hjälp av ändamålsenliga metoder och medel i överensstämmelse med nationell lagstiftning och/eller praxis.
Förbättring av arbetarskyddet för arbetstagarna är ett mål som inte skall underordnas rent ekonomiska hänsyn.
Arbetsgivare skall vara skyldiga att hålla sig à jour med de senaste tekniska och vetenskapliga framstegen vad gäller arbetsplatsens utformning med beaktande av de risker som är förbundna med deras verksamhet och att informera de arbetstagarrepresentanter, som enligt detta direktiv har rätt att ta del av sådan information, på ett sådant sätt att en högre skyddsnivå kan säkerställas.
Utan att det inskränker strängare existerande eller framtida gemenskapsbestämmelser skall detta direktiv tillämpas på alla risker och i synnerhet på dem som härrör från hanteringen av de kemiska, fysiologiska och biologiska agenser, som omfattas av direktiv 80/1107/EEG(6), senast ändrat genom direktiv 88/642/EEG(7).
En kommitté bestående av ledamöter nominerade av medlemsstaterna behöver tillsättas för att bistå kommissionen med de tekniska bearbetningarna för de särdirektiv, som föreskrivs i detta direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. För det ändamålet innehåller direktivet dels allmänna principer för att förebygga yrkesbetingade risker, för arbetarskydd, för att eliminera riskfaktorer och faktorer, som kan förorsaka olycksfall, för information, samråd, avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis samt utbildning av arbetstagarna och deras representanter, dels allmänna riktlinjer för genomförandet av dessa principer.
3. Detta direktiv skall inte hindra tillämpningen av sådana gällande eller framtida bestämmelser i medlemsstaterna och i gemenskapen som är gynnsammare vad gäller skyddet för arbetstagarnas säkerhet och hälsa.
Artikel 2
Räckvidd
1. Detta direktiv skall tillämpas på all verksamhet, såväl privat som offentlig ( industri, jordbruk, handel, förvaltning, tjänster, undervisning, kultur- och fritidsverksamhet etc.).
2. Detta direktiv skall inte tillämpas på sådana offentliga verksamheter, där det inte kan undvikas att förhållanden som är speciella för dessa verksamheter kommer i konflikt med direktivet, exempelvis försvaret eller polisen eller viss specifik verksamhet inom civilförsvaret.
I dessa fall skall arbetstagarnas säkerhet och hälsa tryggas så långt möjligt mot bakgrund av direktivets syften.
Artikel 3
Definitioner
I detta direktiv avses med
a) arbetstagare, varje person anställd av en arbetsgivare, inklusive praktikanter och lärlingar men inte arbetstagare i arbetsgivarens hushåll,
b) arbetsgivare, varje fysisk eller juridisk person som står i ett arbetsgivarförhållande till arbetstagare och har ansvar för företaget och/eller verksamheten,
c) arbetstagarrepresentanter med särskilt ansvar för arbetstagarnas säkerhet och hälsa, varje person, som i enlighet med nationell lagstiftning och/eller praxis har utsetts, valts eller utnämnts att representera arbetstagarna i arbetarskyddsfrågor,
d) förebyggande, alla mått och steg som vidtas eller planeras i något skede av verksamheten för att förebygga eller minska risker i arbetet.
Artikel 4
1. Medlemsstaterna skall vidta tillräckliga åtgärder för att säkerställa att arbetsgivare, arbetstagare och arbetstagarrepresentanter omfattas av sådana lagar och andra författningar som behövs för att bestämmelserna i detta direktiv skall kunna genomföras i praktiken.
2. Medlemsstaterna skall i synnerhet se till att en ändamålsenlig kontroll och tillsyn säkerställs.
AVSNITT II ARBETSGIVARNAS SKYLDIGHETER
Artikel 5
Allmänna bestämmelser
1. Arbetsgivaren är skyldig att svara för att arbetstagarens säkerhet och hälsa tryggas i alla avseenden som är förbundna med arbetet.
2. I de fall en arbetsgivare i överensstämmelse med artikel 7.3 anlitar tjänster eller personer utifrån skall han inte fritas från sitt ansvar på detta område.
3. Arbetstagarnas skyldigheter på arbetarskyddsområdet skall inte inverka på arbetsgivarens ansvar.
Artikel 6
Arbetsgivarens allmänna skyldigheter
1. Inom ramen för sina skyldigheter skall arbetsgivaren vidta tillräckliga åtgärder till skydd för arbetstagarnas säkerhet och hälsa, inbegripet förebyggande av risker i arbetet och tillhandahållande av information och utbildning samt iordningställande av erforderlig organisation och nödvändiga resurser.
Arbetsgivaren skall vara uppmärksam på behovet av att avpassa dessa åtgärder med hänsyn till ändrade omständigheter och sträva efter att förbättra de rådande förhållandena.
2. Arbetsgivaren skall verkställa de åtgärder som avses i punkt 1 första stycket med utgångspunkt från följande allmänna principer för förebyggande arbete:
3. Utan att det inskränker de övriga bestämmelserna i detta direktiv skall arbetsgivaren göra följande med beaktande av verksamhetens art:
a) Arbetsgivaren skall utvärdera riskerna för arbetstagarnas säkerhet och hälsa, bland annat vid val av arbetsutrustning, de kemiska ämnen och preparat som används samt arbetsplatsernas utformning.
Som en följd av denna utvärdering, skall vid behov de förebyggande åtgärder samt de arbets- och produktionsmetoder, som tillämpas av arbetsgivaren
- garantera en förbättring av skyddsnivån för arbetstagarna med avseende på säkerhet och hälsa,
- integreras i all verksamhet och på alla nivåer inom företaget och/eller verksamheten.
b) Då arbetsgivaren uppdrar åt arbetstagaren att utföra vissa arbetsuppgifter skall han ta hänsyn till dennes kunskaper på arbetarskyddsområdet.
c) Arbetsgivaren skall se till att planläggning och införande av ny teknik blir föremål för överläggningar med arbetstagarna och/eller deras representanter i fråga om följdverkningarna för arbetstagarnas säkerhet och hälsa i samband med val av utrustning och förändringar i arbetsbetingelser och arbetsmiljön.
d) Arbetsgivaren skall vidta lämpliga åtgärder för att säkerställa att endast de arbetstagare, som fått tillräckliga instruktioner, får tillträde till särskilt riskfyllda och farliga områden.
4. Utan att det inskränker övriga bestämmelser i detta direktiv skall arbetsgivare, där flera företag samtidigt driver verksamhet på ett arbetsställe, samverka vid tillämpningen av reglerna om säkerhet, hälsa och arbetshygien samt, med beaktande av verksamhetens art, samordna sina åtgärder i skyddshänseende och i frågor som rör förebyggande av risker i arbetet samt underrätta varandra och sina respektive arbetstagare och/eller arbetstagarrepresentanter om dessa risker.
5. Åtgärder som rör säkerhet, hygien och hälsa i arbetet får under inga förhållanden medföra några kostnader för arbetstagarna.
Artikel 7
Skydds- och förebyggande åtgärder
1. Utan att det inskränker skyldigheterna enligt artiklarna 5 och 6 skall arbetsgivaren ge en eller flera arbetstagare i uppgift att verka för skydd mot och förebyggande av risker i arbetet inom företaget och/eller verksamheten.
2. De utsedda arbetstagarna skall inte på något sätt missgynnas på grund av sin verksamhet med avseende på skyddsfrågor och förebyggande arbete.
De utsedda arbetstagarna skall ges skälig tid för att kunna fullgöra sina skyldigheter enligt detta direktiv.
4. I de fall då arbetsgivaren anlitar sakkunnig hjälp utifrån skall han informera de personer som anlitas om de faktorer som påverkar eller misstänks påverka arbetstagarnas säkerhet och hälsa och personerna skall ha tillgång till sådan information som avses i artikel 10.2.
5. Under alla omständigheter skall
- de utsedda arbetstagarna ha tillräckliga kunskaper och resurser,
- utifrån anlitade företag eller personer ha tillräckliga kunskaper och tillräckliga personella och professionella resurser, och
6. Ansvaret för åtgärder till skydd mot och förebyggande av de risker för säkerhet och hälsa, som avses i denna artikel, skall åligga en eller flera arbetstagare eller en eller flera enheter inom eller utanför företaget och/eller verksamheten.
Arbetstagaren/arbetstagarna och/eller enheten/enheterna skall vid behov samarbeta.
7. Med hänsyn tagen till verksamheternas art och företagens storlek skall medlemsstaterna ange de verksamhetsgrenar, där arbetsgivaren, under förutsättning att han har kompetens, själv kan ta ansvaret för de åtgärder som avses i punkt 1.
8. Medlemsstaterna skall definiera de erforderliga färdigheter och kvalifikationer som avses i punkt 5.
De kan fastställa det erforderliga antal, som åsyftas i punkt 5.
Artikel 8
Första hjälpen, brandbekämpning, utrymning, allvarlig och överhängande fara
1. Arbetsgivaren skall
- upprätta alla behövliga kontakter med utomstående serviceorgan, framför allt i fråga om första hjälpen, akutvård, räddningsarbete och brandbekämpning.
2. I överensstämmelse med punkt 1 skall arbetsgivaren framför allt ifråga om första hjälpen och utrymning avdela de arbetstagare som behövs för att genomföra sådana åtgärder.
Dessa arbetstagare skall vara tillräckligt många, de skall erhålla fullgod utbildning och ha tillgång till ändamålsenlig utrustning med beaktande av företagets och/eller verksamhetens storlek och särskilda risker.
3. Arbetsgivaren skall
a) så snart som möjligt informera alla arbetstagare, som utsätts eller kan utsättas för allvarlig och överhängande fara, om risken i fråga och om vidtagna eller planerade skyddsåtgärder,
b) vidta åtgärder och ge anvisningar så att alla arbetstagare i händelse av allvarlig, överhängande och oundviklig fara kan avbryta arbetet och/eller omedelbart avlägsna sig från sin arbetsplats och sätta sig i säkerhet,
c) utom i sådana undantagsfall då det finns väl underbyggda skäl för det, avhålla sig från att anmoda arbetstagarna att återgå till arbetet i ett läge, där en allvarlig och överhängande fara fortfarande föreligger.
4. Arbetstagare som vid en allvarlig, överhängande och oundviklig fara lämnar sin arbetsplats och/eller ett farligt område skall inte på något sätt missgynnas på grund av detta utan skall skyddas mot alla skadliga och orättfärdiga följdverkningar i enlighet med nationell lagstiftning och/eller praxis.
5. Arbetsgivaren skall säkerställa att alla arbetstagare, i fall då en allvarlig och överhängande fara för arbetstagarnas och/eller andras säkerhet föreligger, och då den närmast ansvariga arbetsledningen inte kan kontaktas, kan vidta lämpliga åtgärder med hänsyn till sin kunskap och de tekniska resurser, som står till deras förfogande, för att avvärja en sådan fara.
Arbetstagarnas åtgärder får inte leda till att de på något sätt missgynnas, såvida de inte handlat vårdslöst eller visat grov försumlighet.
Artikel 9
Arbetsgivarens skyldigheter i övrigt
1. Arbetsgivaren skall
a) se till att det finns en riskvärdering av miljöfaktorer på arbetsplatsen, inbegripet faktorer för sådana grupper som är utsatta för speciella risker,
b) besluta om de skyddsåtgärder som skall vidtas och den eventuella personliga skyddsutrustning som skall användas,
c) föra ett register över arbetsolycksfall, som resulterat i att arbetstagaren varit arbetsoförmögen under mer än tre dagar,
d) i enlighet med nationell lagstiftning och/eller praxis upprätta rapporter över arbetsolycksfall, som drabbat arbetstagarna.
2. Medlemsstaterna skall fastställa, med hänsyn till verksamhetens art och företagens storlek, de skyldigheter som åvilar skilda grupper av företag i fråga om upprättande av de handlingar som avses i punkt 1 a och b och vid utarbetande av handlingar enligt punkt 1 c och d.
Artikel 10
Information till arbetstagarna
1. I enlighet med nationell lagstiftning och/eller praxis som kan ta hänsyn till bland annat företagets/verksamhetens storlek skall arbetsgivaren vidta lämpliga åtgärder så att arbetstagare och /eller deras representanter i företaget och/eller verksamheten får all den information som behövs om
a) arbetsmiljörisker och skydds- och förebyggande åtgärder och verksamhet med avseende såväl på företaget och/eller verksamheten i stort som varje enskild arbetsplats och/eller varje enskilt arbete,
b) de åtgärder som vidtas i enlighet med artikel 8.2.
2. Arbetsgivaren skall vidta lämpliga åtgärder så att arbetsgivare för anställda i utomstående företag och/eller verksamheter, vilka utför arbete i den förstnämndes företag och/eller verksamhet, i enlighet med nationell lagstiftning och/eller praxis, får den information om förhållandena enligt punkterna 1 a och b som skall lämnas arbetstagarna ifråga.
3. Arbetsgivaren skall vidta lämpliga åtgärder, så att arbetstagare med särskilda uppgifter i skyddsfrågor eller arbetstagarrepresentanter med särskilt ansvar för skyddsfrågor, för de skall kunna utföra sina uppgifter och i enlighet med nationell lagstiftning och praxis, får tillgång till
a) den riskvärdering samt information om de skyddsåtgärder som avses i artikel 9.1 a och b,
b) det register och de rapporter som åsyftas i artikel 9.1 c och d,
c) den kunskap som skydds- och förebyggande åtgärder, tillsynsmyndigheter och arbetsmiljöansvariga organ avkastar.
Artikel 11
Samråd med och medverkan av arbetstagare
1. Arbetsgivarna skall inhämta synpunkter från arbetstagarna och/eller deras representanter och låta dem delta i diskussioner om alla frågor som gäller säkerhet och hälsa på arbetsplatsen.
Detta förutsätter
- överläggningar med arbetstagarna,
- rätt för arbetstagarna och/eller deras representanter att lägga fram förslag,
- avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis.
2. Arbetstagare eller arbetstagarrepresentanter med särskilt ansvar för skyddsfrågor skall ges rätt till avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis, eller rådfrågas i förväg och i god tid beträffande
a) varje åtgärd som på ett väsentligt sätt kan påverka arbetsmiljön,
b) utseende av arbetstagare enligt artikel 7.1 eller 8.2 och den verksamhet som avses i artikel 7.1,
c) den information som åsyftas i artiklarna 9.1 och 10,
d) i förekommande fall, anlitande av tjänster eller personer utifrån enligt artikel 7.3,
e) den planering och uppläggning av utbildningen som avses i artikel 12.
3. Arbetstagarrepresentanter med särskilt ansvar för skyddsfrågor skall ha rätt att anmoda arbetsgivaren att vidta lämpliga åtgärder och lägga fram förslag i syfte att minska riskerna för arbetstagarna och/eller undanröja källan till faran.
4. De arbetstagare, som avses i punkt 2, och de arbetstagarrepresentanter, som avses i punkterna 2 och 3, får inte missgynnas på något sätt på grund av sin verksamhet enligt punkterna 2 och 3.
6. I överensstämmelse med nationell lagstiftning och/eller praxis har arbetstagare och/eller arbetstagarrepresentanter rätt att vända sig till den arbetsmiljöansvariga myndigheten med klagomål, om de anser att de åtgärder som arbetsgivaren vidtagit inte är tillräckliga för att uppnå säkerhet och hälsa på arbetsplatsen.
Arbetstagarrepresentanter skall ges tillfälle att lägga fram sina iakttagelser i samband med inspektionsbesök av den behöriga myndigheten.
Artikel 12
Utbildning av arbetstagare
1. Arbetsgivaren skall säkerställa att varje arbetstagare får tillräcklig utbildning i arbetsmiljöfrågor, framför allt i form av information och instruktioner, som har direkt anknytning till platsen där han arbetar eller hans arbetsuppgifter i samband med
- anställning,
- förflyttning eller byte av arbete,
- införande av ny arbetsutrustning eller ändring av arbetsutrustning,
- införande av ny teknik.
Utbildningen skall
- anpassas till nya eller ändrade risksituationer, och
- vid behov upprepas regelbundet.
2. Arbetsgivaren skall säkerställa att anställda i utomstående företag och/eller verksamheter som utför arbete för arbetsgivarens räkning har fått tillräckliga instruktioner ifråga om arbetsmiljörisker som gäller deras arbete i arbetsgivarens företag och/eller verksamhet.
3. Arbetstagarrepresentanter med särskilda uppgifter i skyddsfrågor skall ha rätt till tillräcklig utbildning.
4. Den utbildning som avses i punkterna 1 och 3 får inte bekostas av arbetstagarna eller arbetstagarrepresentanterna.
Den utbildning som åsyftas i punkt 1 skall förläggas till arbetstid.
Den utbildning som avses i punkt 3 skall förläggas till arbetstid och i enlighet med nationell praxis äga rum inom eller utanför företaget och/eller verksamheten.
AVSNITT III ARBETSTAGARNAS SKYLDIGHETER
Artikel 13
1. Det åligger varje arbetstagare att så långt möjligt sörja för sin egen och andra personers säkerhet och hälsa, i den mån de påverkas av hans handlingar eller förtroendeuppdrag i arbetet, i enlighet med hans utbildning och arbetsgivarens instruktioner.
Artikel 14
Hälsokontroll
1. Åtgärder skall vidtas i enlighet med nationell lagstiftning och/eller praxis i syfte att tillförsäkra arbetstagarna hälsokontroller anpassade till de arbetsmiljörisker, som de utsätts för i arbetet.
2. De åtgärder som avses i punkt 1 skall vara av sådan karaktär att varje arbetstagare, som så önskar, kan genomgå regelbundna hälsokontroller.
3. Hälsokontrollen kan ingå som en del av den allmänna sjukvården.
Artikel 15
Riskgrupper
Särskilt utsatta riskgrupper skall skyddas mot de faror som speciellt berör dem.
Artikel 16
1. Efter förslag från kommissionen med stöd av artikel 118a i fördraget skall rådet anta särdirektiv, bland annat på de områden som uppräknas i bilagan.
2. Utan att det inskränker det förfarande som avses i artikel 17 i fråga om tekniska justeringar får detta direktiv och särdirektiven ändras i enlighet med artikel 118a i fördraget.
3. Bestämmelserna i detta direktiv skall fullt ut tillämpas på alla områden, som omfattas av särdirektiven utan att hindra tillämpningen av de strängare eller mer specifika bestämmelser som finns i särdirektiven.
Artikel 17
Kommitté
1. När rent tekniska justeringar av de särdirektiv som föreskrivs i artikel 16.1 görs för att ta hänsyn till
- antagandet av direktiv om teknisk harmonisering och standardisering, och/eller
- den tekniska utvecklingen, ändringar i internationella regler eller specifikationer och nya rön,
skall kommissionen biträdas av en kommitté bestående av företrädare för medlemsstaterna och med en företrädare för kommissionen som ordförande.
2. Kommissionens företrädare skall till kommittén lämna ett förslag till åtgärder som skall vidtas.
Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande ärendet är.
Beslut om yttrandet skall fattas med tillämpning av de omröstningsregler som enligt fördragets artikel 148.2 gäller för beslut som rådet skall fatta på förslag av kommissionen.
Vid omröstningen i kommittén skall de röster som avges av representanterna för medlemsstaterna vägas enligt artikeln i fördraget. Ordföranden får inte delta i omröstningen.
3. Kommissionen skall anta förslaget, om det har tillstyrkts av kommittén.
Om förslaget inte har tillstyrkts av kommittén eller om den inte avger något yttrande, skall kommissionen utan dröjsmål föreslå rådet åtgärder. Rådet skall besluta med kvalificerad majoritet.
Om rådet inte fattar beslut inom tre månader från det att förslaget har mottagits, skall kommissionen besluta att de föreslagna åtgärderna skall vidtas.
Artikel 18
Slutbestämmelser
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de redan har antagit eller som de antar på det område som omfattas av detta direktiv.
3. Medlemsstaterna skall vart femte år rapportera till kommissionen om den praktiska tillämpningen av bestämmelserna i detta direktiv, och om arbetsgivarnas och arbetstagarnas synpunkter.
Kommissionen skall informera Europaparlamentet, rådet, Ekonomiska och sociala kommittén och Rådgivande kommittén för arbetarskyddsfrågor.
4. Kommissionen skall regelbundet överlämna en rapport till Europaparlamentet, rådet och Ekonomiska och sociala kommittén om tillämpningen av detta direktiv med beaktande av punkterna 1, 2 och 3.
Artikel 19
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av kommissionens förslag(),
med beaktande av Europaparlamentets yttrande(),
med beaktande av Ekonomiska och sociala kommitténs yttrande(),
och med beaktande av följande: När rådet antog direktiv 83/183/EEG(), förband sig rådet att enhälligt på kommissionens förslag införa bestämmelser som tillåter en avsevärd lättnad i eller rent av avlägsnande av formaliteterna för beviljande av skattebefrielser vid permanent införsel från en medlemsstat av enskildas personliga egendom. Särskilda kommittén för ett Medborgarnas Europa inbjöd i sin första rapport, som bekräftades av Europeiska rådet i Bryssel av den 29 och 30 mars 1985, kommissionen att presentera ett sådant förslag.
Det är nödvändigt att i möjligaste mån underlätta den fria rörligheten för personer inom gemenskapen.
I avvaktan på att skattegränserna upphävs såsom behövs för att uppnå en verklig inre marknad, är det nödvändigt att harmonisera och lätta på vissa formaliteter som krävs för beviljandet av den införselbefrielse som föreskrivs i direktiv 83/183/EEG, särskilt vad beträffar upprättandet av en förteckning över egendomen och bevisning om den normala hemvisten. Det är nödvändigt att lätta på gällande regler om användningstiden för importerad egendom och de kvantitativa begränsningarna för vissa artiklar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 83/183/EEG ändras på följande sätt:
1. Artikel 2.2 b skall ersättas med följande:
"b) som personen i fråga faktiskt har haft i bruk innan bytet av hemvist genomfördes eller andrabostaden inrättades. I fråga om motorfordon (inklusive tillhörande släpvagnar), husvagnar och husbilar, nöjesbåtar och privatflygplan, får medlemsstaterna kräva att den flyttande har haft dem i bruk minst sex månader före bytet av hemvist.
För de varor som avses i punkt a andra meningen får medlemsstaterna kräva att den flyttande skall ha haft dem i bruk före flyttningen minst
- tolv månader då det gäller motorfordon (inklusive tillhörande släpvagnar), husvagnar och husbilar, nöjesbåtar och privatflygplan,
3. Artikel 5.1 skall ersättas med följande:
4. I artikel 7 görs följande ändringar:
a) Punkt 1 blir punkt 1 a,
b) I punkt 1 skall följande stycke tillfogas:
5. I artikel 8.2 görs följande ändringar:
a) Orden "under en tid av minst tolv månader" i slutet av första stycket skall ersättas med "före inrättandet av andrabostaden".
b) Tredje stycket skall utgå.
6. I artikel 9 görs följande ändringar:
a) Början av punkt 1 skall ersättas med följande:
"1. Utan att det påverkar tillämpningen av artiklarna 2 5, skall var och en vid giftermål vara berättigad till befrielse från de skatter som avses i artikel 1 när han till den medlemsstat dit han avser att flytta inför personlig egendom som han förvärvat eller har haft i bruk, förutsatt att".
b) Punkt 2 skall ersättas med följande:
"2. Skattebefrielse skall också beviljas för sedvanliga bröllopsgåvor till någon som uppfyller de villkor som fastställs i punkt 1 från personer som har sin normala hemvist i en annan medlemsstat än den dit införsel sker. Befrielsen skall gälla för gåvor med ett enhetsvärde av högst 350 ecu. Medlemsstaterna får dock bevilja skattebefrielse då gränsen 350 ecu överskrids förutsatt att värdet av varje skattebefriad gåva inte överstiger 1 400 ecu".
7. I artikel 11 görs följande ändringar:
a) I punkt 1 skall orden "Fram till ikraftträdandet av de gemenskapsskatteregler som införs i överensstämmelse med artikel 14.2 i direktiv 77/388/EEG skall medlemsstaterna" utgå och punkten inleds därefter med "Medlemsstaterna skall".
b) I punkt 2 skall hänvisningen till "artikel 2.2" ersättas med hänvisning till "artikel 2.2a".
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 11 december 1989 om veterinära kontroller vid handeln inom gemenskapen i syfte att fullborda den inre marknaden (89/662/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Gemenskapen kommer att vidta åtgärder för att stegvis upprätta den inre marknaden under tiden fram till den 31 december 1992.
För att samordningen av marknaden med kreatursprodukter och produkter av animaliskt ursprung skall fungera utan störningar krävs att veterinära hinder mot utvecklingen av handeln inom gemenskapen med dessa produkter undanröjs. Den fria rörligheten av jordbruksprodukter är ett grundläggande inslag i samordningen av marknaderna och bör kunna underlätta en rationell utveckling av jordbruksproduktionen och ett optimalt utnyttjande av produktionsmedlen.
På det veterinära området utnyttjas för närvarande gränserna för att utföra kontroller som syftar till att värna om hälsan hos människor och djur.
Det slutliga målet är att de veterinära kontrollerna skall utföras enbart vid avsändningsstället. För att uppnå detta krävs en harmonisering av de grundläggande krav som rör hälsoskyddet för människor och djur.
Målet är att förverkliga den inre marknaden och i avvaktan på att detta uppnås bör huvudvikten läggas på de kontroller som skall utföras hos avsändaren och på att organisera de kontroller som skulle kunna utföras på destinationsorten. En sådan lösning skulle innebära ett slopande av de veterinära kontrollerna vid gränserna mellan medlemsstaterna.
Denna lösning förutsätter ett ökat förtroende för de veterinära kontroller som utförs av den avsändande staten. Den senare måste säkerställa att dessa veterinära kontroller utförs på ett lämpligt sätt.
I destinationslandet skulle veterinära stickprovskontroller kunna utföras hos mottagarna. Vid allvarlig misstanke om felaktigheter skulle dock den veterinära kontrollen kunna utföras medan varorna är på väg.
Det är en uppgift för medlemsstaterna att lägga fram en plan över hur de avser att utföra kontrollerna. Dessa planer bör underställas gemenskapen för godkännande.
Ett förfarande bör fastställas för att bilägga eventuella tvister i fråga om sändningar från någon anläggning, något produktionsställe eller något företag.
Behovet av skyddsåtgärder måste uppmärksammas. Inom detta område, måste, inte minst med hänsyn till effektiviteten, ansvaret i första hand falla på den avsändande medlemsstaten. Kommissionen måste kunna vidta snabba åtgärder, särskilt genom att göra besök på platsen och vidta de åtgärder som läget kräver.
För att vara effektiva måste de regler som fastställs i detta direktiv täcka alla varor som är underkastade veterinära krav i samband med handel inom gemenskapen.
Dock föreligger alltjämt med avseende på vissa epizootiska sjukdomar olika hälsosituationer inom medlemsstaterna och i avvaktan på ett ställningstagande från gemenskapens sida vad gäller sätten att bekämpa dessa sjukdomar bör frågan om kontroll av handeln med husdjur inom gemenskapen tills vidare lämnas utanför och en kontroll av handlingar bör vara tillåten under transporten. Med hänsyn till det rådandet läget vad gäller frågan om harmonisering och i avvaktan på gemenskapsregler bör varor som inte är underkastade harmoniserade regler uppfylla de krav som gäller inom destinationslandet, förutsatt att de senare står i överensstämmelse med artikel 36 i fördraget.
Bestämmelserna i gällande direktiv bör anpassas till de nya regler som fastställs i detta direktiv.
Dessa regler bör ses över på nytt före utgången av år 1993.
Kommissionen bör bemyndigas att vidta åtgärder för tillämpningen av detta direktiv. I detta syfte bör det utarbetas rutiner för att upprätta ett nära och effektivt samarbete mellan kommissionen och medlemsstaterna inom Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Medlemsstaterna skall se till att de veterinära kontroller som skall utföras på produkter av animaliskt ursprung, som omfattas av de direktiv som räknas upp i bilaga A eller i artikel 14 och som är avsedda för handel, inte längre sker vid gränserna utan verkställs i enlighet med detta direktiv, utan att det påverkar tillämpningen av artikel 6.
Artikel 2
I detta direktiv avses med
1. veterinär kontroll: varje fysisk undersökning eller administrativt förfarande som gäller de varor som avses i artikel 1 och som syftar till att direkt eller på annat sätt värna om människors eller djurs hälsa,
2. handel: handel mellan medlemsstater med varor som avses i artikel 9.2 i fördraget,
3. anläggning: varje företag som producerar, lagrar eller bearbetar produkter som avses i artikel 1,
4. behörig myndighet: den centrala myndighet i en medlemsstat som det åligger att utföra veterinära kontroller eller varje myndighet till vilken denna uppgift har överförts,
5. officiell veterinär: den veterinär som förordnats av den behöriga centrala myndigheten i medlemsstaten.
Artikel 3
1. Medlemsstaterna skall se till att inga andra produkter görs till föremål för handel än sådana som avses i artikel 1 och som har anskaffats, kontrollerats, stämplats och märkts i enlighet med gemenskapens regler för den angivna destinationen och som fram till den slutlige mottagare som uppgivits åtföljs av ett hälsointyg, djurhälsocertifikat eller något annat dokument som fastställts genom gemenskapens veterinära bestämmelser.
De anläggningar som produkterna härrör ifrån skall genom kontinuerlig egenkontroll säkerställa att produkterna uppfyller de krav som uppställts i föregående stycke.
Utan att påverka de tillsynsskyldigheter som åligger den officiella veterinären i enlighet med gemenskapens lagstiftning skall den behöriga myndigheten utföra regelbunden kontroll vid anläggningarna för att försäkra sig om att de för handel avsedda produkterna uppfyller gemenskapens krav eller, i de fall som avses under punkt 3 i denna artikel och i artikel 14, de krav som gäller i den mottagande medlemsstaten.
När det finns anledning att misstänka att kraven inte uppfylls skall den behöriga myndigheten utföra nödvändiga kontroller och, i de fall misstanken bekräftas, vidta lämpliga åtgärder, vilket kan innefatta indragning av godkännandet.
2. När transporten innefattar flera destinationer skall produkterna sammanföras till ett antal partier som svarar mot antalet destinationer. Varje parti skall åtföljas av det ovannämnda certifikatet eller dokumentet.
När de produkter som åsyftas i artikel 1 är avsedda för export till ett tredje land skall transportproceduren stå under tullövervakning fram till den ort där sändningen lämnar gemenskapens territorium.
3. Medlemsstater som valt att föra in produkter från vissa länder utanför gemenskapen skall meddela kommissionen och övriga medlemsstater om förekomsten av sådan import.
När produkterna förs in till gemenskapens territorium via en annan medlemsstat än någon av dem som avses ovan skall denna medlemsstat verkställa en kontroll i handlingarna av ursprunget och varornas destination i enlighet med artikel 6.1.
De medlemsstater till vilka varorna är destinerade skall förbjuda att de berörda produkterna sänds vidare från deras territorium såvida de inte är avsedda för någon annan medlemsstat som begagnar sig av samma införselmöjlighet.
Artikel 4
1. Medlemsstater från vilka varorna avsänds skall vidta de åtgärder som krävs för att säkerställa att de berörda parterna uppfyller de veterinära kraven i samtliga led av produktion, lagring, saluföring och transport av de produkter som avses i artikel 1. De skall särskilt säkerställa att
- de produkter som anskaffats i enlighet med de direktiv som avses i bilaga A kontrolleras på samma sätt ur veterinär synpunkt, oavsett om de är avsedda för handel inom gemenskapen eller för den inhemska marknaden.
- de produkter som omfattas av bilaga B inte förs ut till någon annan medlemsstats territorium, om de inte kan försäljas inom medlemsstatens eget territorium av skäl som har stöd i artikel 36 i fördraget.
Artikel 5
1. Mottagande medlemsstater skall vidta följande åtgärder:
a) Den behöriga myndigheten får på destinationsorten för varorna genom icke-diskriminerande veterinära stickprov kontrollera att de krav som uppställs i artikel 3 har uppfyllts. Provtagning får ske samtidigt.
När den behöriga myndigheten i den medlemsstat genom vilken varorna transiteras eller den medlemsstat till vilken varorna avsänts har fått uppgifter som ger anledning till misstanke om att gällande bestämmelser överträtts, får kontroller som innefattar kontroll av transportsättet också utföras under transporten av varor till medlemsstatens territorium.
b) När de produkter som avses i artikel 1 och som härrör från en annan medlemsstat är avsedda
- för en anläggning som står under tillsyn av en officiell veterinär, skall denne se till att endast sådana produkter släpps in i denna anläggning som uppfyller kraven i artikel 3.1 med avseende på märkning och medföljande dokument eller, vad gäller de produkter som avses i bilaga B, åtföljs av de dokument som fastställs i destinationslandets bestämmelser,
- för en godkänd distributör som delar upp partierna eller för ett handelsföretag med många filialer, eller någon verksamhet som inte är underkastad ständig tillsyn skall den senare, innan partiet delas upp eller saluföras, kontrollera att varorna märkts och att de intyg eller dokument som avses i den första strecksatsen finns tillgängliga samt anmäla varje felaktighet eller avvikelse till den behöriga myndigheten.
- för andra mottagare, särskilt när partiet till en del har lossats under transporten, skall förpackningen i enlighet med artikel 3.1 åtföljas av originalet till det intyg som avses i den första strecksatsen.
De garantier som skall företes av de mottagare som avses i andra och tredje strecksatserna skall specificeras i ett avtal med den behöriga myndigheten att undertecknas vid tiden för den registrering som föreskrivits i punkt 3. Den behöriga myndigheten skall utföra stickprovskontroller för att förvissa sig om att dessa garantier uppfylls.
2. Om gemensamma varustandarder inte fastställts genom gemenskapsregler och i det fall som avses i artikel 14 kan den mottagande medlemsstaten, utan att det påverkar tillämpningen av artikel 4 och med vederbörlig hänsyn till de allmänna bestämmelserna i fördraget, kräva att ursprungsanläggningen skall följa de regler som gäller enligt den ifrågavarande medlemsstatens nationella lagstiftning. Den medlemsstat från vilken produkterna härrör skall se till att den ifrågavarande produkten uppfyller dessa normer.
3. För importörer som får produkter levererade till sig från en annan medlemsstat eller som helt delar upp ett parti av sådana produkter gäller att
a) de dessförinnan skall bli föremål för registrering, om den behöriga myndigheten kräver detta,
b) de skall föra ett register i vilket sådana leveranser noteras,
c) de skall, om den behöriga myndigheten kräver detta, anmäla ankomsten av sådana produkter från en annan medlemsstat i den mån detta är nödvändigt för att utföra de kontroller som avses under punkt 1,
d) de skall under den tid som fastställts av den behöriga myndigheten, dock under minst sex månader, arkivera de hälsointyg och dokument som avses i artikel 3 för att vid anfordran företes för den behöriga myndigheten.
4. Närmare bestämmelser för tillämpning av denna artikel skall utformas i enlighet med det förfarande som fastställs i artikel 18.
5. Rådet skall med ledning av en rapport från kommissionen som åtföljs av eventuella ändringsförslag på nytt se över denna artikel inom tre år från det att detta direktiv börjar tillämpas.
Artikel 6
1. I samband med den kontroll som företas på de platser där produkter kan införas till gemenskapens territorium från tredje land, däribland hamnar, flygplatser och gränsstationer mot tredje land, skall medlemsstaterna se till att följande åtgärder vidtas:
a) Kontroller av handlingar skall göras rörande produkternas ursprung.
b) Vid införsel av produkter från länder utanför gemenskapen, skall de sändas under tullövervakning till inspektionsställen där veterinär besiktning kan utföras.
De produkter som avses i bilaga A får inte godkännas vid tullklarering annat än om dessa kontroller har visat att de uppfyller gemenskapens bestämmelser.
De produkter som avses i bilaga B och de varor som medlemsstaterna har valt att importera i enlighet med artikel 3.3 och som efter att ha införts till gemenskapens territorium skall vidarebefordras till en annan medlemsstats territorium skall
- antingen underkastas veterinär besiktning som visar att de uppfyller de bestämmelser som utfärdats i den medlemsstat till vilken de destinerats, eller
- efter enbart visuell besiktning för att fastställa att dokument och produkter stämmer överens, vidarebefordras under tullövervakning till destinationsorten, där veterinär besiktning skall utföras.
c) Produkter som härrör från gemenskapen skall inspekteras i enlighet med de besiktningsbestämmelser som fastställs i artikel 5.
2. Dock skall från den 1 januari 1993 och utan hinder av punkt 1 alla produkter som transporteras genom reguljära och direkta transportmedel som förbinder två geografiska punkter inom gemenskapen vara underkastade de bestämmelser om inspektion som fastställs i artikel 5.
Artikel 7
1. Om den behöriga myndigheten i en medlemsstat i samband med den inspektion som utförs på destinationsorten eller under transporten konstaterar
a) förekomst av smittämnen som orsakar någon av de sjukdomar som nämns i direktiv 82/894/EEG(4), senast ändrat genom kommissionens beslut 89/162/EEG(5), någon zoonos eller sjukdom eller något annat som kan tänkas orsaka allvarlig fara för djur och människor eller om produkterna kommer från ett område som är smittat med en epizootisk sjukdom, skall de utom vad gäller djurhälsoaspekter, i fråga om produkter som är föremål för någon av de behandlingar som avses i artikel 4 i direktiv 80/215/EEG(6), senast ändrat genom direktiv 88/660/EEG(7), beordra att transportförpackningen i fråga förstörs eller används på något annat sätt som fastställts genom gemenskapsregler.
Kostnader i samband med förstöring av partiet skall betalas av avsändaren eller dennes ombud.
De behöriga myndigheterna i den mottagande medlemsstaten skall omedelbart genom telex delge de övriga medlemsstaternas behöriga myndigheter och kommissionen vad som framkommit vid inspektionen, vilka beslut som fattats och på vilka grunder de fattats.
De skyddsåtgärder som anges i artikel 9 får tillämpas.
Utöver detta får kommissionen på begäran av en medlemsstat och i enlighet med det förfarande som fastställs i artikel 17, när det uppkommer situationer som inte förutsetts av gemenskapens lagstiftning, vidta varje åtgärd som är nödvändig för att uppnå samstämmighet i medlemsstaternas handlande.
b) att varorna inte uppfyller de villkor som fastställts genom gemenskapens direktiv, eller nationella normer när ett beslut om de gemenskapsnormer som föreskrivits genom direktiven inte fattats, och förutsatt att hänsynen till människors och djurs hälsa tillåter det, låta avsändaren eller hans ombud välja mellan att
- förstöra varorna eller
- använda dem för något annat ändamål, däribland att sända tillbaka dem efter att att ha inhämtat medgivande från den behöriga myndigheten i ursprungslandet.
Om intyget eller dokumenten befinns innehålla felaktigheter skall dock avsändaren medges en tidsfrist innan den sistnämnda möjligheten tillgrips.
2. I enlighet med det förfarande som fastställs i artikel 18 skall kommissionen upprätta en förteckning över de smittämnen och sjukdomar som avses i punkt 1 och fastställa detaljerade regler för hur denna artikel skall tillämpas.
Artikel 8
1. I de fall som avses i artikel 7 skall den behöriga myndigheten i den mottagande medlemsstaten utan dröjsmål ta kontakt med de behöriga myndigheterna i den medlemsstat från vilken varorna avsänts. De sistnämnda myndigheterna skall vidta alla nödvändiga åtgärder och meddela den behöriga myndigheten i den förstnämnda medlemsstaten vilka kontroller som utförts, vilka beslut som fattats och motiveringen för dessa.
Om myndigheten i den första medlemsstaten befarar att dessa åtgärder är otillräckliga, skall de behöriga myndigheterna i de två medlemsstaterna gemensamt söka finna en lösning. Om det är lämpligt kan detta innefatta inspektion på platsen.
Om de kontroller som avses i artikel 7 visar upprepade oegentligheter, skall den behöriga myndigheten i den mottagande medlemsstaten underrätta kommissionen och de veterinära myndigheterna i de övriga medlemsstaterna.
Kommissionen får på begäran av den behöriga myndigheten i den mottagande medlemsstaten eller på eget initiativ och under hänsynstagande till arten av överträdelsen
- sända en inspektionsgrupp till den berörda anläggningen, eller
- uppdra åt en officiell veterinär, vars namn skall finnas med på en av kommissionen på förslag av medlemsstaterna upprättad förteckning och som kan godkännas av de olika berörda parterna, för att kontrollera fakta vid den berörda anläggningen,
- uppmana den behöriga myndigheten att intensifiera provtagningen av den berörda anläggningens produkter.
Den skall underrätta medlemsstaterna om vad som framkommit.
När dessa åtgärder vidtagits för att komma tillrätta med upprepade oegentligheter vid någon anläggning skall kommissionen debitera den berörda anläggningen alla utgifter som uppkommit genom tillämpning av strecksatserna i föregående stycke.
I avvaktan på vad kommissionen kommit fram till skall den medlemsstat från vilken sändningen härrör, på begäran av den mottagande medlemsstaten, utöka kontrollen av de produkter som kommer från den ifrågavarande anläggningen och tillfälligt dra in tillståndet om det föreligger starka skäl för detta med hänsyn till djurs och människors hälsa.
Den mottagande medlemsstaten får å sin sida utöka kontrollerna av produkter som kommer från samma anläggning.
På begäran av någon av de två berörda medlemsstaterna - om oegentligheterna har bekräftats av experternas utlåtanden - skall kommissionen i enlighet med det förfarande som fastställs i artikel 17, vidta lämpliga åtgärder som får utsträckas till att bemyndiga medlemsstaterna att införa ett tillfälligt förbud mot införsel till sina territorier av produkter som härrör från den berörda anläggningen. Dessa åtgärder skall bekräftas eller omprövas snarast möjligt i enlighet med det förfarande som fastställs i artikel 17.
De allmänna reglerna för tillämpningen av denna artikel skall fastställas i enlighet med förfarandet i artikel 18.
2. Rätten enligt medlemsstatens gällande lagstiftning att begära prövning av beslut som fattats av de behöriga myndigheterna skall inte påverkas av detta direktiv.
Beslut som fattats av den behöriga myndigheten i den mottagande staten skall tillsammans med en motivering delges avsändaren eller hans ombud och den behöriga myndigheten i den medlemsstat från vilken partiet avsänts.
Om avsändaren eller hans ombud begär detta, skall de ifrågavarande besluten tillsammans med motivering vidarebefordras till honom i skriftlig form med uppgifter om den rätt till prövning som står till buds i enlighet med gällande lagstiftning i den mottagande medlemsstaten, tillsammans med uppgift om hur och inom vilken tid detta skall ske.
Om tvist skulle uppkomma, och utan att det påverkar tillämpningen av den nyssnämnda rätten till prövning, får dock de två berörda parterna, om överenskommelse träffas om detta inom en period av högst två månader, hänskjuta tvisten för avgörande till någon expert vars namn finns med på en av kommissionen upprättad förteckning över gemenskapens experter. Kostnaden för att anlita denna expert skall betalas av gemenskapen.
Dessa experter skall yttra sig inom högst 72 timmar. Parterna skall avvakta expertens yttrande med vederbörlig hänsyn tagen till gemenskapens veterinära lagstiftning.
3. Kostnaderna för att sända tillbaka varorna, lagra dem, överföra dem till annan användning eller förstöra dem skall betalas av mottagaren.
Artikel 9
Den medlemsstat från vilken sändningen utgått skall omedelbart vidta de kontroll- och försiktighetsåtgärder som fastställs i gemenskapsreglerna, däribland särskilt fastställande av buffertzoner som avses i dessa regler eller vidta varje annan åtgärd som den finner lämplig.
Den mottagande medlemsstaten eller den genom vilken sändningen skall transiteras, som i samband med någon av de kontroller som avses i artikel 5 har konstaterat förekomst av någon av de sjukdomar eller orsaker som avses i första stycket, får om så krävs vidta de försiktighetsmått som fastställs i gemenskapens regler.
I avvaktan på att åtgärder vidtas i enlighet med punkt 4 får den mottagande medlemsstaten, när särskilt allvarliga folk- eller djurhälsoskäl föreligger, vidta tillfälliga skyddsåtgärder gentemot de berörda anläggningarna eller, i fråga om en epizootisk sjukdom, vad gäller det skyddsområde som fastställs i gemenskapens regler.
De åtgärder som vidtagits av medlemsstaterna skall utan dröjsmål anmälas till kommissionen och till de övriga medlemsstaterna.
2. På begäran av den medlemsstat som avses i första stycket i punkt 1, eller på initiativ av kommissionen, får en eller flera kommissionsledamöter omedelbart bege sig till den berörda platsen för att i samarbete med de behöriga myndigheterna undersöka vilka åtgärder som vidtagits. De skall avge ett yttrande om dessa åtgärder.
3. Om kommissionen inte har informerats om vilka åtgärder som vidtagits, eller om den anser de vidtagna åtgärderna otillräckliga, får den, i samarbete med den berörda medlemsstaten och i avvaktan på att den Ständiga veterinärkommittén sammanträder, vidta tillfälliga skyddsåtgärder gentemot produkter från den region som berörs av den epizootiska sjukdomen eller produkter från en viss anläggning. Dessa åtgärder skall underställas Ständiga veterinärkommittén snarast möjligt för att fastställas, ändras eller upphävas i enlighet med förfarandet i artikel 17.
4. Kommissionen skall i samtliga fall vid första lämpliga tillfälle ta ställning till situationen på nytt i Ständiga veterinärmedicinska kommittén. Den skall besluta om vilka åtgärder som behöver tillgripas för de produkter som avses i artikel 1 och, om situationen så kräver, för de ursprungliga produkterna eller de produkter som härletts från dessa produkter i enlighet med förfarandet i artikel 17. Kommissionen skall följa läget och i enlighet med samma förfarande ändra eller upphäva de beslut som fattats alltefter vad situationen kräver.
5. Utförliga regler för hur denna artikel skall tillämpas och särskilt förteckningen över de zoonoser eller orsaker som kan tänkas utgöra ett allvarlig hot mot människors hälsa skall utarbetas i enlighet med förfarandet i artikel 18.
Artikel 10
Varje medlemsstat och kommissionen skall utse den eller de veterinärmyndigheter som skall svara för de veterinära kontrollerna och samarbetet med de andra medlemsstaternas inspektionsmyndigheter.
Artikel 11
Medlemsstaterna skall se till att tjänstemännen inom deras veterinärmyndigheter, om så är lämpligt i samarbete med tjänstemännen inom andra myndigheter som anförtrotts denna uppgift särskilt ges fullmakt och möjlighet att
- verkställa inspektioner av lokaler, kontor, laboratorier, installationer, transportmedel, anläggningar och utrustning, rengörings- och underhållsmedel och de rutiner som används vid framställning, bearbetning, kontrollmärkning, märkning och presentation av dessa produkter,
- kontrollera att personalen uppfyller de krav som fastställs i de texter som avses i bilaga A,
- ta prover på produkter som finns i lager för att förvaras, släppas ut på marknaden eller transporteras,
- granska skriftligt eller datoriserat material som är av betydelse för de kontroller som verkställs utöver de åtgärder som vidtagits med stöd av artikel 3.1.
För detta ändamål skall de inspekterade anläggningarna vara beredda att samarbeta med kontrollanterna i den utsträckning som krävs för att de skall kunna fullgöra sina åligganden.
Artikel 12
1. Artikel 8.3 och artiklarna 10 och 11 i direktiv 64/433/EEG(8), senast ändrat genom direktiv 88/657/EEG(9), utgår.
2. Artikel 5.3 och 5.4 och artiklarna 9, 10 och 11 i direktiv 71/118/EEG(10), senast ändrat genom direktiv 88/657/EEG, utgår.
3. I direktiv 74/461/EEG(11), senast ändrat genom direktiv 87/489/EEG(12),
i) skall artiklarna 5.2, 5.3, 5.4 och 5.5 och artiklarna 6 och 8, utgå, och
ii) i artikel 8a skall hänvisningen till artikel 8 ersättas med en hänvisning till artikel 9 i direktiv 89/662/EEG.
4. Artikel 7.3 och artiklarna 12 och 16 i direktiv 77/99/EEG(13), senast ändrat genom direktiv 89/227/EEG(14), utgår.
5. I direktiv 80/215/EEG
i) skall artikel 5.2, 5.3, 5.4 och 5.5 och artiklarna 6 och 7 utgå, och
ii) i artikel 7a skall hänvisningarna till artikel 7 ersättas med en hänvisning till artikel 9 i direktiv 89/662/EEG.
6. Artikel 5.3 och 5.4 och artiklarna 7, 8 och 12 i direktiv 85/397/EEG(15), ändrat genom förordning (EEG) nr 3768/85(16), utgår.
7. Artikel 10.1 och 10.3 i direktiv 88/657/EEG utgår.
8. Artiklarna 8 och 9 i direktiv 89/437/EEG(17) utgår.
9. I bilaga B till direktiv 72/462/EEG(18) skall följande läggas till i intyget: "Första mottagarens namn och adress".
Artikel 13
1. Följande artikel skall läggas till direktiven 64/433/EEG och 71/118/EEG:
"Artikel 19
2. Följande artikel skall läggas till direktiven 72/461/EEG och 80/215/EEG:
"Artikel 15
3. Följande artikel läggs till direktiv 77/99/EEG:
"Artikel 24
4. Följande artikel skall läggas till direktiven 85/397/EEG och 88/657/EEG:
"Artikel 18
5. Följande artikel läggs till direktiv 88/437/EEG:
"Artikel 17
Artikel 14
Fram till och med den 31 december 1992 skall, i avvaktan på beslut om att gemenskapsregler skall antas, handeln med de produkter som räknas upp i bilaga B vara underkastade de regler om kontroll som fastställs i detta direktiv, särskilt de som fastställs i artikel 5.2.
Medlemsstaterna skall före det datum som fastställs i artikel 19 meddela vilka villkor och förfaranden som för närvarande tillämpas vid handeln med de produkter som avses i första stycket.
Rådet skall, efter förslag från kommissionen, före den 31 december 1991 fastställa de slutliga reglerna vad gäller handel med de produkter som räknas upp i bilaga B.
Artikel 15
I artikel 9 i direktiv 64/432/EEG(19)skall följande punkt införas:
"2 a En eller flera kommissionsledamöter får, på begäran av en medlemsstat eller på initiativ av kommissionen själv, genast bege sig till den berörda platsen för att, i samarbete med de behöriga myndigheterna, granska de åtgärder som vidtagits och avge ett yttrande om dessa åtgärder."
Artikel 16
1. Medlemsstaterna skall senast tre månader före det datum som fastställs i artikel 19.1 tillställa kommissionen ett program som redovisar de nationella åtgärder som kommer att vidtas för att förverkliga de angivna målen med detta direktiv, särskilt hur ofta kontrollerna kommer att utföras.
2. Kommissionen skall granska de program som överlämnats av medlemsstaterna i enlighet med punkt 1.
3. Varje år från och med 1991 skall kommissionen till medlemsstaterna överlämna en rekommendation till program för kontroller att genomföras påföljande år. Den ständiga veterinärkommittén skall i förväg ha avgivit sitt yttrande om rekommendationen som får bli föremål för senare anpassningar.
Artikel 17
3. Kommissionen skall själv anta förslaget om det är förenligt med yttrandet från kommittén.
4. Om förslaget inte är förenligt med yttrandet från kommittén eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas.
Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte har fattat något beslut inom 15 dagar från det att förslaget kommit det till handa, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas, såvida inte rådet med enkel majoritet har avvisat förslaget.
Artikel 18
1. När det förfarande som fastställs i denna artikel skall tillämpas, skall ordföranden utan dröjsmål hänskjuta ärendet till den ständiga veterinärmedicinska kommittén (i det följande kallad "kommittén") som inrättats genom beslut 68/361/EEG.
2. Företrädaren för kommissionen skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. De röster som avgivits av företrädarna för medlemsstaterna skall vägas enligt samma artikel i fördraget. Ordföranden får inte rösta.
3. Kommissionen skall godkänna de tilltänkta åtgärderna om de är förenliga med kommitténs yttrande.
4. Om förslaget inte är förenligt med yttrandet från kommittén eller om inget yttrande avgives, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas.
Rådet skall fatta sitt beslut med kvalificerad majoritet.
Artikel 19
1. Före den 31 december 1990 skall rådet fatta sitt beslut med kvalificerad majoritet om kommissionens förslag rörande veterinärkontroller vid handel mellan medlemsstaterna med levande djur.
Före det datum som nämns i första stycket skall rådet med kvalificerad majoritet fatta beslut, efter förslag från kommissionen, om de regler och allmänna principer som skall gälla vid de kontroller av införsel från länder utanför gemenskapen av varor som omfattas av detta direktiv. Före detta datum skall på samma sätt kontrollstationer vid de yttre gränserna inrättas och de krav fastställas som dessa gränsstationer skall uppfylla.
2. Före den 31 december 1992 skall rådet se över bestämmelserna i detta direktiv och med ledning av en rapport från kommissionen om de erfarenheter som vunnits, tillsammans med relevanta förslag, fatta beslut om dessa med kvalificerad majoritet.
Artikel 20
Fram till den 31 december 1992 får medlemsstaterna för att tillåta gradvis införande av de kontrollarrangemang som fastställs i detta direktiv, utan hinder av artikel 5.1
- upprätthålla kontroller av handlingar under transporten av kött och produkter som härrör från kött för att säkerställa att de speciella krav rörande mul- och klövsjuka och svinpest som fastställs genom gemenskapsregler uppfylls,
- verkställa kontroller av handlingar under transporten av produkter som importerats från tredje land och som är avsedda för medlemsstaterna.
Artikel 21
Rådet skall före den 1 oktober 1992, med kvalificerad majoritet efter förslag från kommissionen, bestämma vilka arrangemang som skall tillämpas när de övergångsbestämmelser som fastställs i artikel 20 upphör att gälla.
Artikel 22
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv vid ett datum som skall fastställas genom det beslut som skall fattas före den 31 december 1990, i enlighet med andra stycket i artikel 19.1, dock senast den 31 december 1991.
Dock skall Grekland ges en ytterligare ett års respit med att följa det.
Artikel 23
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 21 december 1989 om samordning av lagar och andra författningar för prövning av offentlig upphandling av varor och bygg- och anläggningsarbeten (89/665/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag (1),
i samarbete med Europaparlamentet (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
med beaktande av följande: Gemenskapens direktiv om offentlig upphandling, särskilt rådets direktiv 71/305/EEG av den 26 juli 1971 för samordning av förfarandena vid tilldelning av bygg- och anläggningsarbeten (4), senast ändrat genom direktiv 89/440/EEG (5) och rådets direktiv 77/62/EEG av den 21 december 1976 om samordningar av förfarandet vid offentlig upphandling av varor (6), senast ändrat genom direktiv 88/295/EEG (7), innehåller ej bestämmelser som säkrar deras effektiva tillämpning.
Gällande bestämmelser för tillämpning av direktiven på såväl nationell som gemenskapsnivå är inte alltid tillräckliga för att garantera efterlevnad av i sammanhanget relevanta gemenskapsregler, i synnerhet inte i ett skede, då överträdelser kan korrigeras.
Då man öppnar det offentliga upphandlingsområdet för konkurrens mellan medlemsstaterna, krävs en väsentligt större garanti för insyn och icke-diskriminering. För att detta skall ha påtaglig verkan, måste snabba och effektiva rättsmedel stå till buds i händelse av överträdelse av gemenskapsrättens regler för offentlig upphandling eller av nationell lagstiftning om genomförandet av sådana regler.
Eftersom upphandlingsförfarandet för varje särskilt kontrakt är kortvarigt, måste ett sakkunnigt prövningsorgan bl.a. vara behörigt att vidta interimistiska åtgärder i syfte att uppskjuta förfarandet hos myndigheten eller verkställigheten av dess beslut. Med hänsyn till tidsfaktorn måste vidare ges möjlighet att snabbt ingripa mot nämnda överträdelser.
Det är nödvändigt att se till att lämpliga förfaranden finns inom alla medlemsstater, så att beslut i strid mot dess bestämmelser kan upphävas och ersättning kan ges till dem som skadats av överträdelserna.
Om företagen inte begär prövning, torde rättelse i vissa fall aldrig komma till stånd, såvida man inte inrättar en särskild ordning för ändamålet.
Följaktligen bör kommissionen ges behörighet att föra ärendet inför vederbörande myndigheter i medlemslandet såväl som upphandlingsmyndigheten, så snart den anser, att en klar och konkret överträdelse har begåtts vid upphandlingsförfarandet, så att lämpliga åtgärder vidtas för skyndsam rättelse av en påstådd kränkning.
Tillämpningen av detta direktiv bör utvärderas inom en period av fyra år från genomförandet på grundval av information från medlemsstaterna om prövningsförfarandets funktion i respektive länder.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Medlemsstaterna skall vidta nödvändiga åtgärder för att garantera, att en upphandlande myndighets beslut prövas effektivt, vad beträffar upphandling inom ramen för direktiv 71/305/EEG och 77/62/EEG. I synnerhet skall prövningar göras skyndsamt enligt reglerna i följande artiklar, där särskilt uppmärksammas artikel 2.7 för de fall upphandlingsbeslut innefattar överträdelse av gemenskapsrätten för offentlig upphandling eller nationella bestämmelser om införande av sådan lag.
2. Medlemsstaterna skall förhindra diskriminering mellan företag, vilka vid upphandling gör gällande skada till följd av den åtskillnad som görs i detta direktiv mellan nationella bestämmelser om införande av gemenskapsrätten och andra nationella bestämmelser.
3. Medlemsstaterna skall se till att ett prövningsförfarande med detaljerade regler enligt medlemsstaternas bestämmande införs och att det kan åberopas av var och en, som har eller har haft intresse av att få avtal om viss offentlig upphandling av varor eller bygg- och anläggningsarbeten, och som har skadats eller riskerat att skadas av en påstådd överträdelse. Det förutses, att en medlemsstat skall kunna kräva av den person som begär prövning, att han dessförinnan meddelat den avtalsslutande myndigheten att han hävdar förekomsten av diskriminering, och att han ämnar söka prövning.
Artikel 2
1. Medlemsstaterna skall se till att införda bestämmelser om prövning enligt artikel 1 innefattar behörighet att
a) så tidigt som möjligt vidta interimistiska åtgärder för att rätta påstådda överträdelser eller förhindra ytterligare skada för berörda intressen, inklusive åtgärder för att uppskjuta eller garantera uppskjutandet av upphandlingsförfarandet liksom att förhindra verkställighet av den upphandlande myndighetens beslut,
b) antingen åsidosätta eller garantera åsidosättande av olagliga beslut, vilket innefattar undanröjandet av diskriminerande tekniska, ekonomiska eller finansiella specifikationer i anbuds- eller kontraktshandlingarna eller i varje annat dokument som har samband med upphandlingen,
c) ge ersättning åt en person, som skadats av överträdelse.
2. Behörighet enligt punkt 1 får ges till separata organ med ansvar för olika sidor av prövningsförfarandet.
3. Prövningsförfarandet i sig behöver inte automatiskt bidra till att upphandlingen skjuts upp.
5. Medlemsstaterna får bestämma att, i de fall skada görs gällande på grund av att beslut tillkommit i strid mot lag, det överklagade beslutet först skall upphävas av ett organ med nödvändig behörighet för detta.
6. Verkan av att behörighet har utövats enligt punkt 1 på ett redan slutet avtal om upphandling skall regleras i nationell lag.
Medlemsstaterna får dessutom bestämma att, utom i fall där ett beslut måste undanröjas innan ersättning ges ut, prövningsorganets behörighet sedan ett upphandlingsavtal genomförts skall begränsas till att lämna ersättning till den som lidit skada av överträdelsen.
7. Medlemsstaterna skall se till att införa bestämmelser, som garanterar, att granskningsorganens beslut verkligen åtlyds.
8. För de fall prövningsorganen ej utgörs av rättsliga instanser gäller, att skriftliga beslutsmotiveringar alltid skall ges. Dessutom gäller för dessa fall, att det måste finnas en möjlighet att pröva påstådda olagliga åtgärder vidtagna av sådana organ i en rättslig instans eller en domstol som avses i fördragets artikel 177, oberoende av såväl upphandlingsmyndigheten som prövningsorganet.
Medlemmarna i ett sådant oberoende organ skall tillsättas och frånträda på samma villkor som gäller för rättsliga instanser, tillämpade av den myndighet som utnämner och avsätter dem, samt bestämmer ämbetsperiodens längd. Åtminstone ordföranden i prövningsorganet skall ha domarkompetens. Det oberoende organet skall fatta sina beslut i ett förfarande, där båda parter hörs, och besluten skall vara lagligen bindande enligt regler bestämda av medlemsstaten.
Artikel 3
1. Kommissionen får tillgripa prövningsförfarandet enligt denna artikel, om den innan ett upphandlingskontrakt slutits anser, att en klar och konkret överträdelse av gemenskapsreglerna har ägt rum vid en offentlig upphandling inom områdena för direktiven 71/305/EEG och 77/62/EEG.
2. Kommissionen skall underrätta den berörda medlemsstaten och den upphandlande myndigheten om de skäl, som föranlett bedömningen att en klar och konkret överträdelse föreligger och kräva rättelse.
3. Inom 21 dagar från mottagandet av underrättelsen enligt punkt 2 skall medlemsstaten till kommissionen avge
a) bekräftelse på att överträdelsen har rättats till,
b) förklaring till varför rättelse ej skett, eller
c) uppgift om att upphandlingsförfarandet har avbrutits, antingen på upphandlingsmyndighetens eget initiativ, eller på grundval av maktbefogenheter som givits i artikel 2.1 a.
4. En förklaring enligt punkt 3 b kan bl.a. vila på, att den påstådda överträdelsen redan är föremål för rättslig eller annan undersökning eller prövningsförfarande enligt artikel 2.8. I sådant fall måste medlemsstaten underrätta kommissionen om resultatet av detta, så snart det blir känt.
5. Då uppgift har lämnats om att en upphandling har avbrutits enligt punkt 3 c, skall medlemsstaten underrätta kommissionen om när upphandlingsförfarandet återupptas, eller när någon annan upphandlingsprocedur med hel eller delvis anknytning till upphandlingen påbörjats. Underrättelsen skall bekräfta, att den påstådda överträdelsen har rättats eller om så inte är fallet, skälen till varför rättelse inte har skett.
Artikel 4
2. Medlemsstaterna skall årligen före den 1 mars rapportera till kommissionen om sin tillämpning av prövningsbestämmelserna under föregående kalenderår. Anvisningar om rapportens innehåll utarbetas av kommissionen i samråd med Rådgivande kommittén för offentlig upphandling.
Artikel 5
Medlemsstaterna skall före den 1 december 1991 införa de bestämmelser som är nödvändiga för att följa detta direktiv. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning och andra författningar som de antar inom det område som omfattas av detta direktiv.
Artikel 6
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av rådets förordning (EEG) nr 2658/87(1) av den 23 juli 1987, om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan, senast ändrad genom förordning (EEG) nr 20/89(2), särskilt artikel 9 i denna, och
med beaktande av följande: För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser angående klassificering av de varor som anges i bilagan till den här förordningen.
Förordning (EEG) nr 2658/87 fastställer de allmänna bestämmelserna för tolkningen av Kombinerade nomenklaturen och dessa bestämmelser gäller också varje annan nomenklatur som helt eller delvis grundar sig på denna eller som lägger ytterligare underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser med tanke på tillämpningen av tulltaxebestämmelser eller andra bestämmelser som rör varuhandeln.
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt de tillämpliga KN-nummer som anges i kolumn 2 av de skäl som anges i kolumn 3.
Nomenklaturkommittén har inte yttrat sig över förslaget inom den tid som ordföranden bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i tabellen i bilagan klassificeras nu inom Kombinerade nomenklaturen enligt de till- lämpliga KN-nummer som anges i kolumn 2 i denna tabell.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom förordning (EEG) nr 20/89(2), särskilt artikel 9 i denna, och
med beaktande av följande: För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen som är en bilaga till förordning (EEG) nr 2658/87 vad avser tulltaxeklassificering av anoraker, skidjackor, vindjackor och liknande artiklar som omfattas av bl.a. KN-nummer 6101, 6102, 6201 och 6202, är det nödvändigt att ange vissa kännetecknande egenskaper för dessa klädesplagg.
Dessa klädesplagg är av det slag som i allmänhet bärs utanpå andra kläder och som skyddar mot vind, kyla och regn.
Klädesplagg utan ärmar eller med korta ärmar ger inte detta skydd. Det är därför nödvändigt att ange att anoraker, vindjackor och liknande artiklar, som nämns ovan, måste ha långa ärmar.
Nomenklaturkommittén har inte avgivit något yttrande inom den tid som dess ordförande bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Endast klädesplagg med långa ärmar skall klassificeras som anoraker, skidjackor, vindjackor och liknande artiklar enligt KN-nummer 6101, 6102, 6201 och 6202.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska atomenergigemenskapen, särskilt artikel 31 i detta,
med beaktande av kommissionens förslag, som utformats efter yttrande av en grupp experter utsedda av Vetenskapliga och tekniska kommittén(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Bilagan till förordning (Euratom) nr 3954/87(4) innehåller rubriker för gränsvärden för livsmedel och djurfoder.
För somliga rubriker hade dock inga gränsvärden fastställts i avvaktan på beslut av rådet efter ytterligare utredning, främst av vetenskapliga experter.
Kommissionen framlade två meddelanden till rådet, den 14 juni respektive den 9 december 1988. De var avsedda som tillägg till bilagan till förordningen och hade utarbetats efter samråd med expertgruppen som avses i artikel 31 i fördraget.
Därför bör det göras tillägg till bilagan till förordningen.
Vissa andra uppgifter i denna bilaga bör också anpassas till de senaste vetenskapliga rönen inom detta område.
Därför verkar det lämpligt att sammanföra gränsvärdena och andra uppgifter i denna bilaga i en enda tabell.
Med hänsyn till det fortsatta arbetet bör det också föreskrivas att förfarandet i artikel 7 i förordning (Euratom) nr 3954/87 också tillämpas för att fastställa gränsvärden för djurfoder. Det bör därför göras lämpliga tillägg till förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (Euratom) nr 3954/87 skall ersättas med bilagan till denna förordning.
Artikel 2
Artikel 7 i förordning (Euratom) nr 3954/87 skall ersättas med följande:
"Artikel 7
Tillämpningsföreskrifter till denna förordning, en lista över mindre viktiga livsmedel tillsammans med de gränsvärden som skall tillämpas på dessa, samt gränsvärden för djurfoder, skall antas enligt artikel 30 i förordning (EEG) 804/68, som skall tillämpas på motsvarande sätt. För detta ändamål skall en kommitté tillsättas."
Artikel 3
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 64/433/EEG av den 26 juni 1964 om hygienproblem som påverkar handeln med färskt kött inom gemenskapen(1), senast ändrat genom direktiv 86/587/EEG((2), särskilt artikel 13 i detta, och
med beaktande av följande: I enlighet med artikel 13 i direktiv 64/433/EEG och i enlighet med förfarandet i artikel 16 får på begäran undantag från punkt 45 c i bilaga 1 beviljas varje medlemsstat som lämnar liknande garantier. Vid sådana undantag skall hygienkrav som lägst motsvarar kraven i nämnda bilaga fastställas.
I brev av den 26 september 1989 har myndigheterna i Spanien till kommissionen framfört en begäran om undantag från punkt 45 c i bilaga 1 till direktiv 64/433/EEG i fråga om styckning av färskt nötkött, fårkött och griskött. I begäran föreslås hygienkrav. Det är nödvändigt att de alternativa hygienkrav som fastställs i det begärda undantaget i fråga om styckning av färskt kött lägst motsvarar kraven i punkt 45 c i bilaga 1 till direktiv 64/433/EEG.
De hygienkrav som föreslås a
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 64/433/EEG av den 26 juni 1964 om hygienproblem som påverkar handeln med färskt kött inom gemenskapen(1), senast ändrat genom direktiv 88/657/EEG(2), särskilt artikel 13 i detta, och
med beaktande av följande: I enlighet med artikel 13 i direktiv 64/433/EEG och i enlighet med förfarandet i artikel 16 får på begäran undantag från punkt 45 c i bilaga 1 beviljas varje medlemsstat som lämnar liknande garantier. Vid sådana undantag skall hygienkrav som lägst motsvarar kraven i nämnda bilaga fastställas.
I brev av den 18 januari 1989 har myndigheterna i Frankrike till kommissionen framfört en begäran om undantag från punkt 45 c i bilaga 1 till direktiv 64/433/EEG i fråga om styckning av färskt nötkött, fårkött och griskött. I begäran föreslås hygienkrav. Det är nödvändigt att de alternativa hygienkrav som fastställs i det begärda undantaget i fråga om styckning av färskt kött lägst motsvarar kraven i punkt 45 c i bilaga 1 till direktiv 64/433/EEG.
De hygienkrav som föreslås a
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87(1) om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan, senast ändrad genom förordning (EEG) nr 3945/89(2), särskilt artikel 9 i denna, och med beaktande av följande:
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till förordning (EEG) nr 2658/87, är det nödvändigt att fastställa bestämmelser för klassificering av de varor som anges i bilagan till den här förordningen.
I förordning (EEG) nr 2658/87 fastställs allmänna bestämmelser för tolkningen av Kombinerade nomenklaturen och dessa gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna, eller som lägger ytterligare underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser med tanke på tillämpningen av tulltaxebestämmelser eller andra bestämmelser som rör varuhandeln.
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt de tillämpliga KN-nummer som anges i kolumn 2, av de skäl som anges i kolumn 3.
Nomenklaturkommittén har inte yttrat sig inom den tid som ordföranden bestämt vad gäller produkt nr 4 i tabellen i bilagan.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Nomenklaturkommittén vad gäller produkterna nr 1, 2, 3, 5 och 6 i tabellen i bilagan.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i tabellen i bilagan klassificeras nu inom Kombinerade nomenklaturen enligt de tillämpliga KN-nummer som anges i kolumn 2 i denna tabell.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS BESLUT av den 2 maj 1991 om erkännande av Australien som fritt från Erwinia amylovora (Burr.) Winsl. et al. (91/261/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 77/93/EEG av den 21 december om skyddsåtgärder mot att skadegörare på växter eller växtprodukter förs in till medlemsstaterna(1), senast ändrat genom kommissionens direktiv 91/27/EEG(2), särskilt bilaga 3 del B 10 i detta, och med beaktande av följande:
Enligt bestämmelserna i direktiv 77/93/EEG får växter av vissa släkten, med undantag för frukter och fröer, med ursprung i andra länder eller regioner än dem som har erkänts vara fria från Erwinia amylovora (Burr.) Winsl. et al. inte föras in till vissa medlemsstater från och med den 16 april till och med den 31 oktober om växterna har sitt ursprung på norra halvklotet samt från och med den 1 november till och med den 15 april om de har sitt ursprung på södra halvklotet.
Det framgår av officiella uppgifter som Australien har tillhandahållit att den ovan nämnda skadegöraren inte förekommer där och att landet länge har upprätthållit ett strängt förbud mot import av växter och växtprodukter som kan föra med sig denna skadegörare.
Det kan därför fastslås att det inte finns någon risk för spridning av den ovan nämnda skadegöraren.
Detta beslut inverkar inte på senare upptäckter som kan visa att den ovan nämnda organismen förekommer i landet.
Kommissionen kommer att säkerställa att Australien årligen tillhandahåller alla de tekniska uppgifter som är nödvändiga för att bedöma den ovan nämnda situationen.
De åtgärder som föreskrivs i detta beslut är förenliga medyttrandet från Ständiga kommittén för växtskydd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE. Artikel 1
Härmed förklaras att Australien erkänns vara fritt från Erwinia amylovora (Burr.) Winsl. et al. Artikel 2
Detta beslut riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 21 mars 1991 om ändring för nionde gången i direktiv 76/769/EEG om tillnärmning av medlemsstaternas lagar och andra författningar om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar) (91/173/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag(1),
i samarbete med Europaparlamentet(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Åtgärder bör vidtas för att stegvis upprätta den inre marknaden under tiden fram till den 31 december 1992. Den inre marknaden skall vara ett område utan inre gränser, inom vilket den fria rörligheten för varor, personer, tjänster och kapital är säkerställd.
Både pentaklorfenol (CAS nr 87-86-5) och dess föreningar är farliga för människan och miljön, särskilt vattenmiljön. Användningen av dessa ämnen bör regleras.
Vissa medlemsstater har redan infört begränsningar i fråga om användning eller utsläppande på marknaden av dessa ämnen eller preparat i vilka de ingår. Åtgärderna inverkar direkt på den inre marknadens upprättande och funktion. En tillnärmning av medlemsstaternas lagstiftning på detta område är således nödvändig. Bilaga 1 till direktiv 76/769/EEG(4), senast ändrat genom direktiv 89/678/EEG(5), bör därför ändras.
Kommissionen kommer att utarbeta en samordnad gemenskapskapsstrategi som avser rätten att släppa ut på marknaden och använda kemiska produkter för träskyddsändamål. Denna strategi utarbetas på grundval av uppgifter som medlemsstaterna lämnar, särskilt om hälso- och miljörisker, och med beaktande av de svårigheter som finns i medlemsstaterna på detta område.
Den gällande gemenskapslagstiftning som avser medlemsstaternas rätt att besluta om mer långtgående begränsningar för användningen av de aktuella ämnena och preparaten i arbetsmiljön berörs inte av detta direktiv.
RÅDETS DIREKTIV av den 16 december 1991 om det ömsesidiga erkännandet av båtförarcertifikat för transport av gods och passagerare på inre vattenvägar (91/672/EEG)
med beaktande av kommissionens förslag (),
Artikel 1
Vid tillämpningen av detta direktiv skall nationella båtförarcertifikat för transport av gods och passagerare på inre vattenvägar enligt bilaga 1 indelas på följande sätt:
Artikel 2
Om inte annat följer av bestämmelserna i artikel 3.5 skall båtförarcertifikat för navigering på Rhen, som utfärdas i överensstämmelse med den reviderade konventionen om sjöfarten på Rhen, gälla för alla vattenvägar inom gemenskapen.
Artikel 3
1. Båtförarcertifikat som fortfarande är giltiga och som är upptagna i grupp A i bilaga 1 skall erkännas av alla medlemsstater som giltiga för navigering på de vattenvägar av havskaraktär som är upptagna i bilaga 2, som om de själva hade utfärdat ifrågavarande båtförarcertifikat.
2. Medlemsstaterna skall ömsesidigt erkänna de båtförarcertifikat som fortfarande är giltiga och som är upptagna i grupp B i bilaga 1 som giltiga för navigering på deras inre vattenvägar, bortsett från dem för vilka behörighetsbeviset för navigering på Rhen erfordras eller sådana som är upptagna i bilaga 2, som om de själva hade utfärdat ifrågavarande båtförarcertifikat.
3. En medlemsstats erkännande av ett båtförarcertifikat enligt grupp A eller grupp B i bilaga 1 får underkastas samma villkor angående minimiålder som de villkor som fastställts i denna medlemsstat för utfärdande av ett båtförarcertifikat i samma grupp.
4. En medlemsstats erkännande av ett båtförarcertifikat får begränsas till de kategorier av fartyg för vilka detta certifikat gäller i den medlemsstat som har utfärdat det.
Medlemsstaterna skall erkänna det certifikat som utfärdas i enlighet med nummer 10 170 i ADNR (förordningen om transport av farligt gods på Rhen) som bevis på dessa kunskaper.
Artikel 4
Om så behövs skall kommissionen vidta nödvändiga åtgärder för att anpassa förteckningen över certifikat i bilaga 1 i enlighet med det förfarande som anges i artikel 7.
Artikel 5
Rådet skall senast den 31 december 1994, på grundval av ett förslag från kommissionen som skall inlämnas senast den 31 december 1993, med kvalificerad majoritet besluta om gemensamma bestämmelser för framförande på inre vattenvägar av fartyg som transporterar gods och passagerare.
Artikel 6
Artikel 7
1. Vid tillämpningen av artikel 4 skall kommissionen biträdas av en kommitté. Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till ändring av bilaga 1. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen varvid medlemsstaternas röster skall vägas enligt angivna artikel. Ordföranden får inte rösta.
Kommissionen skall själv anta ändringen av bilaga 1 om den är förenlig med kommitténs yttrande.
Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta om den föreslagna ändringen.
Artikel 8
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EEG) nr 147/91 av den 22 januari 1991 om definition och fastställande av toleranser för svinn av jordbruksprodukter i offentlig interventionslagring
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3492/90 om fastställande av de faktorer som skall beaktas i årsredovisningarna för finansiering av interventionsåtgärder i form av offentlig lagring genom garantisektionen inom Europeiska utvecklings- och garantifonden för jordbruket(1), särskilt artikel 4 i denna, och
med beaktande av följande: Den definition av toleransen som fastställs i artikel 4 i förordning (EEG) nr 3492/90 för förvaring av jordbruksprodukter i offentliga interventionslager och beräkningsmetoden för bestämning av de finansiella följderna av lagring måste anges närmare.
Denna tolerans avser den normala kvantiteten svinn i samband med normal lagring eller bearbetning av jordbruksprodukter i intervention med beaktande av kraven på riktig förvaring av produkten.
Denna tolerans skall fastställas för varje berörd produkt med hjälp av en enkel metod och mot bakgrund av den oidentifierbara kvantitet svinn som konstaterats i samband med lagring under senare år. Toleransnivån bör därför fastställas som en procentsats av det totala lagret.
För vissa produkter som bearbetas mellan uppköp och lagring skall särskilda toleranser fastställas för svinn i samband med bearbetning.
Inga lagringsåtgärder har förekommit för griskött under lång tid och denna toleransnivå bör fastställas senare om lagringsåtgärder skulle vidtas på nytt.
Tidpunkten för när de finansiella följderna av tillämpningen av toleranser skall beaktas av garantisektionen inom EUGFJ bör fastställas.
För vissa jordbruksprodukter har beräkningsmetoden för procentsatsen för normalt svinn i samband med lagring genomgått grundläggande förändringar. Dessa procentsatser bör därför revideras mot bakgrund av erfarenheten.
Toleranserna har fastställts i sektorsvisa förordningar. De bör av hänsyn till rättslig förenkling fastställas i en enda förordning.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från EUGFJ-kommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE. Artikel 1
1. För varje jordbruksprodukt som är föremål för offentlig lagring fastställs en toleransnivå för kvantiteten svinn i samband lagringsåtgärder som vidtas i enlighet med godkända regler.
2. Toleransen skall fastställas som en procentsats av den faktiska vikten utan emballage av de kvantiteter som placeras i lager och övertas under det aktuella räkenskapsåret, med tillägg för kvantiteter i lager i början av det aktuella räkenskapsåret. Den skall för varje produkt beräknas på grundval av de totala kvantiteter som lagras av ett interventionsorgan.
Den faktiska vikten vid inlagring och utlagring skall beräknas genom att från den registrerade vikten dra den standardvikt för förpackningen som fastställts i uppköpsvillkoren eller, i avsaknad av sådan, den genomsnittliga förpackningsvikt som används av myndigheten.
Artikel 2 1. Procentsatserna för normalt tillåtet svinn vid lagring fastställs härmed till följande:
- urbening av nötkött 32 %
- bearbetning av tobak i blad 19 %.
KOMMISSIONENS FÖRORDNING (EEG) nr 1026/91 av den 22 april 1991 om ändring av förordning (EEG) nr 1208/81 om fastställande av en gemenskapsskala för klassificering av slaktkroppar av fullvuxna nötkreatur
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1358/80 av den 5 juni 1980 om fastställande av orienterings- och interventionspriser för fullvuxna nötkreatur för 1980/1981 års regleringsår och om införande av en gemenskapsskala för klassificering av slaktkroppar av fullvuxna nötkreatur(1), särskilt artikel 4.1 i denna,
med beaktande av kommissionens förslag, och
med beaktande av följande: I förordning (EEG) nr 1208/81(2) fastställs gemenskapens skala för klassificering av slaktkroppar av vuxna nötkreatur.
Med tanke på de genetiska förbättringar som är ett resultat av avel med nötkreatur bör gemenskapens skala för klassificering av slaktkroppar av vuxna nötkreatur anpassas så att hänsyn tas till förekomsten av djur med dubbelmuskulatur. Det bör därför finnas en möjlighet att frivilligt kunna införa en konformationsklass utöver de existerande klasserna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE. Artikel 1
Förordning (EEG) 1208/81 ändras på följande sätt:
1. Artikel 3 skall ersättas med följande:
"Artikel 3
1. Slaktkroppar av vuxna nötkreatur skall indelas i följande kategorier:
A. Slaktkroppar av okastrerade ungdjur av hankön under två år.
B. Slaktkroppar av andra okastrerade djur av hankön.
C. Slaktkroppar av kastrerade djur av hankön.
D. Slaktkroppar av djur av honkön som har kalvat.
E. Slaktkroppar av andra djur av honkön.
Utan att det påverkar gällande interventionsbestämmeler skall bokstäverna A, B, C, D och E användas för att identifiera slaktkroppar från och med den 1 januari 1992.
Kriterier för att skilja slaktkroppskategorier åt skall fastställas i enlighet med förfarandet i artikel 27 i förordning (EEG) nr 805/68.
2. Slaktkroppar av vuxna nötkreatur skall klassificeras genom en bedömning i följdordning av
a) konformation,
b) fettgrupp
enligt definitionerna i bilagorna 1 respektive 2.
Den konformationsklass som betecknas med bokstaven S i bilaga 1 får användas av medlemsstaterna om de vid frivilligt införande av en konformationsklass över de existerande klasserna (djur med dubbelmuskulatur) önskar att ta hänsyn till egenskaperna hos eller den förväntade utvecklingen av en viss produktion.
Medlemsstater som avser att använda denna möjlighet skall meddela kommissionen och övriga medlemsstater detta.
3. Medlemsstater skall vara bemyndigade att dela upp var och en av de klasser som anges i bilagorna 1 och 2 i högst tre underklasser."
2. Bilaga 1 skall ersättas med den bilaga som finns i bilagan till denna förordning.
Artikel 2 Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EEG) nr 1781/91 av den 19 juni 1991 om ändring av förordning (EEG) nr 1014/90 om närmare tillämpningsföreskrifter för definition, beskrivning och presentation av spritdrycker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1576/89 av den 29 maj 1989 om allmänna bestämmelser för definition, beskrivning och presentation av spritdrycker(1), särskilt artikel 6.3 i denna, och med beaktande av följande:
I kommissionens förordning (EEG) nr 1014/90(2) fastställs en första omgång tillämpningsföreskrifter. Dessa behöver kompletteras.
För att ta hänsyn till hävdvunnen praxis som fanns när förordning (EEG) nr 1576/89 trädde i kraft bör det vara tillåtet att behålla vissa sammansatta namn på likörer även om inte alkoholen erhållits eller uteslutande erhållits från den spritdryck som angivits. Det är nödvändigt att specificera villkor för beteckningen för sådana likörer för att undvika varje risk för förväxling med de spritdrycker som definieras i artikel 1.4 i förordning (EEG) nr 1576/89.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för genomförande av regler om spritdrycker.
"Artikel 7b
1. I enlighet med artikel 6.1 andra strecksatsen i förordning (EEG) nr 1576/89, skall användningen av kategoribeteckningar i sammansatta beteckningar vara förbjuden vid presentation av spritdrycker såvida inte alkoholen i drycken uteslutande härrör från den spritdryck som anges.
2. I linje med situationen vid tiden för den här förordningens ikraftträdande får dock följande sammansatta beteckningar användas vid presentation av likörer som framställts i gemenskapen:
solbaerrom, även kallad blackcurrant rum.
3. Vad beträffar märkning och presentation av likörer som anges i punkt 2 skall den sammansatta termen finnas på etiketten på en enda rad med samma typsnitt och färg, och ordet "likör" skall finnas i omedelbar närhet med bokstäver som inte är mindre än det typsnittet.
Artikel 2 Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EEG) nr 2988/91 av den 11 oktober 1991 om ändring av förordning (EEG) nr 1538/91 om tillämpningsföreskrifter till förordning (EEG) nr 1906/90 om vissa handelsnormer för fjäderfäkött
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1906/90 av den 26 juni 1990 om vissa handelsnormer för fjäderfäkött(1), särskilt artikel 9 i denna, och
med beaktande av följande: I artikel 8 i kommissionens förordning (EEG) nr 1538/91(2) fastställs tillämpningsföreskrifter för den valfria klassificeringen av fryst och djupfryst fjäderfäkött i viktklasser. Den omedelbara tillämpningen av dessa bestämmelser har visat sig utgöra ett hinder för importen från tredje land av fjäderfäkött som förpackats före nämnda förordnings ikraftträdande. Tillämpningen av artikel 8 bör därför uppskjutas till den 1 mars 1992.
Förvaltningskommittén för fjäderfäkött och ägg har inte yttrat sig inom den tid som dess ordförande bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Denna förordning träder i kraft den 20 juni 1991.
Till och med den 31 december 1991 får aktörerna emellertid förpacka produkter som omfattas av denna förordning i förpackningsmaterial som är försett med de uppgifter som anges i gemenskapslagstiftningen eller i den nationella lagstiftning som tillämpades före denna förordnings ikraftträdande. Dessa produkter får sedan saluföras till och med den 31 december 1992."
RÅDETS BESLUT av den 13 juli 1992 om datorisering av veterinära förfaranden vid import (Shift-projektet), om ändring av direktiven 90/675/EEG, 91/496/EEG, 91/628/EEG och beslut 90/424/EEG och om upphävande av beslut 88/192/EEG (92/438/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, och särskilt artikel 43 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1), och
Mot bakgrund av den positiva utvecklingen i fråga om harmonisering inom veterinärområdet, bör man fastställa nya bestämmelser om datorisering av veterinärförfarandena vid import och beslut 88/192/EEG bör därför upphävas.
Dessa nya bestämmelser skall bidra till att skydda människors och djurs hälsa samtidigt som de gör det möjligt att genomföra den inre marknaden för djur och animaliska produkter.
Behovet för dessa nya bestämmelser är så mycket större eftersom kontroll vid gränserna mellan medlemsstaterna skall slopas.
Datorisering av veterinärförfarandena vid import bör erbjuda möjligheter för en officiell veterinär som skall avvisa en sändning vid en gränskontrollstation att på ett effektivt sätt förmedla relevanta upplysningar och också omfatta databaser med importvillkor och för import av djur och animaliska produkter.
Direktiv 90/675/EEG, 91/496/EEG och 91/628/EEG bör därför ändras.
Man bör därför inom ramen för rådets beslut 90/424/EEG av den 26 juni 1990 om vissa utgifter på veterinärområdet(6) fastställa att gemenskapen skall bidra till finansieringen av genomförandet av de nya åtgärderna i fråga om datorisering av veterinärförfarandena vid import.
Kommissionen bör få till uppgift att besluta om nödvändiga tillämpningsföreskrifter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Ett system för att förmedla relevant information när en officiell veterinär vid en gränskontrollstation beslutar att vidaresända en sändning.
- Organisation och drift av databaser som innehåller gemenskapens importvillkor för djur och produkter.
- Organisation och drift av databaser som innehåller import till gemenskapen av djur och produkter.
2. Den datorisering som avses i punkt 1 skall uppfylla nuvarande internationell standard.
Artikel 2
I detta beslut skall vid behov de definitioner tillämpas som återfinns i direktiv 90/675/EEG, 91/496/EEG och 91/628/EEG.
Artikel 3
1. Det informationssystem som avses i artikel 1.1 första strecksatsen skall omfatta gränskontrollstationer, medlemsstaternas centrala myndigheter och kommissionen.
2. Det informationssystem som avses i artikel 1.1 första strecksatsen skall fungera enligt principerna i bilaga 1.
Artikel 4
1. De databaser som avses i artikel 1 andra strecksatsen skall innehålla alla upplysningar om importvillkor för import till gemenskapen av djur och produkter och särskilt upplysningar om förteckningar över godkända tredje länder, godkända anläggningar, vidtagna skyddsåtgärder och godkända intygsförebilder.
2. De databaser som avses i artikel 1.1 andra strecksatsen skall organiseras och fungera enligt principerna i bilaga 2.
Artikel 5
1. De databaser som avses i artikel 1.1 tredje strecksatsen skall innehålla alla upplysningar om varje sändning av djur eller produkter som förs in till gemenskapen, särskilt om de transportvillkor för djur som fastställs i kapitel III i direktiv 91/628/EEG och resultaten av de kontroller som utförs i enlighet med direktiv 90/675/EEG och 91/496/EEG.
2. De databaser som avses i artikel 1 tredje strecksatsen skall organiseras och fungera enligt principerna i bilaga 3.
Artikel 6
Den utrustning som används vid gränskontrollstationer vid tillämpning av detta beslut kan vara den som anges i artikel 2.2 i kommissionens beslut 91/398/EEG av den 19 juli 1991 om ett datoriserat nätverk som länkar samman veterinärmyndigheterna (Animo)(7).
Artikel 7
Beslut 88/192/EEG skall härmed upphöra att gälla.
Artikel 8
Direktiv 90/675/EEG skall ändras på följande sätt:
1. Följande strecksats skall läggas till i artikel 4.1:
2. Följande skall läggas till i artikel 8.2:
"d) konsultera de databaser som avses i artikel 1, andra strecksatsen i beslut 92/438/EEG."
3. Följande mening skall läggas till i artikel 9.2 iii:
"Den officiella veterinären skall se till att uppdatering av de databaser som avses i artikel 1 tredje strecksatsen i beslut 92/438/EG utförs."
4. Artikel 11.4 b första strecksatsen skall ersättas med följande:
"- underrätta den officiella veterinären vid kontrollstället på bestämmelseorten om produkternas passage och om trolig ankomstdag via det datoriserade nätverket som länkar samman veterinärmyndigheter (Animo),".
5. Följande mening skall läggas till artikel 11.4 b:
"I så fall skall den behöriga myndigheten informeras via det datoriserade nätverket som länkar samman veterinärmyndigheter (Animo)."
6. I artikel 16.1 a skall första strecksatsen ersättas med följande:
"- aktivera det informationssystem som avses i artikel 1 första strecksatsen i beslut 92/438/EEG."
7. I artikel 16.1 a skall den tredje strecksatsen utgå.
8. Artikel 16.5 skall ersättas med följande:
"5. Bestämmelserna i beslut 92/438/EEG skall tillämpas."
Artikel 9
Direktiv 91/496/EEG ändras på följande sätt:
1. I artikel 4.1 skall följande strecksats läggas till:
"Kontrollen skall göras efter att man har konsulterat de databaser som avses i artikel 1 andra strecksatsen i beslut 92/438/EEG."
3. I artikel 6.2 skall följande mening läggas till:
"Den officiella veterinären skall se till att all uppdatering av de databaser som avses i artikel 1 tredje strecksatsen i beslut 92/438/EEG utförs."
4. I artikel 9.1 d skall orden "som avses i artikel 12.4 andra stycket" ersättas med "som avses i artikel 20 i direktiv 90/425/EEG".
5. I artikel 12.1 c skall första strecksatsen ersättas med följande:
"- aktivera det informationssystem som avses i artikel 1 första strecksatsen i beslut 92/438/EEG".
6. I artikel 12.1 c skall tredje strecksatsen utgå.
7. Artikel 12.4 skall ersättas med följande:
"4. Bestämmelserna i beslut 92/438/EEG skall tillämpas."
8. I artikel 30.2 första stycket skall orden "andra stycket" utgå.
Artikel 10
I artikel 11 i direktiv 91/628/EEG skall följande stycke läggas till:
Artikel 11
Följande artikel skall läggas till i beslut 90/424/EEG:
"Artikel 37 a
1. Ekonomiskt bidrag från gemenskapen kan beviljas för datorisering av veterinärförfarandena vid import enligt beslut 92/438/EEG(*).
Artikel 12
Tillämpningsföreskrifter för detta beslut skall vid behov antas i enlighet med det förfarande som fastställs i artikel 13.
Artikel 13
1. Kommissionen skall bistås av Ständiga veterinärkommittén som bildats genom beslut 68/361/EEG(8), hädanefter kallad 'kommittén`.
2. När det förfarande som anges i denna artikel skall tillämpas skall ordföranden utan dröjsmål hänskjuta ärendet till kommittén antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
3. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande ärendet är. Kommittén skall fatta sitt beslut med en majoritet på 54 röster, varvid medlemsstaternas röster skall vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
4. a) Kommissionen skall själv anta förslaget och tillämpa det omedelbart om det inte strider mot kommitténs yttrande.
b) Om förslaget inte är förenligt med kommitténs yttrande, eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas och tillämpa dem omedelbart.
Artikel 14
Bestämmelserna i detta beslut skall ses över före den 1 juli 1995 för att ta hänsyn till den tekniska utvecklingen och för att göra nödvändiga förbättringar särskilt med hänsyn till ny utveckling som redan kan ha konstaterats i de mest avancerade medlemsstaterna.
Artikel 15
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 25 september 1992 om fastställande av samarbetsformer mellan Animo datacentrum och medlemsstaterna (92/486/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets beslut 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden(1), senast ändrat genom direktiv 92/60/EEG(2) och särskilt artikel 20.3 i detta, och med beaktande av följande:
Kommissionen antog den 19 juli 1991 beslut 91/398/EEG om ett datoriserat system som länkar samman veterinärmyndigheterna (Animo)(3) och den 2 juli 1992 beslut 92/373/EEG om utnämnande av datacentret Animo(4).
I syfte att säkerställa att systemet Animo fungerar smidigt bör åtgärder vidtas för en harmonisering av samarbetsformerna mellan Animo datacentrum och medlemsländerna.
Bestämmelserna i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Varje medlemsstat skall i enlighet med sina nationella bestämmelser utse en myndighet som skall vara ansvarig för samordningen mellan de interna myndigheterna i varje enskild medlemsstat.
Samordningsmyndigheten skall förhandla fram ett kontrakt med Eurokom om användning av det gemensamma datacentret. Kontraktet skall undertecknas i enlighet med nationella bestämmelser.
Artikel 2
De behöriga myndigheterna i medlemsstaterna skall säkerställa det kontrakt som avses i artikel 1
- gäller till den 1 juli 1995,
- innehåller en klausul om årlig översyn,
- innehåller en klausul om uppsägning med sex månaders varsel,
- innehåller en förpliktelse från Eurokom att uppfylla alla de tekniska krav som fastställs i bilagan till kommissionens beslut 91/638/EEG(5), baserade på den tekniska lösning som Eurokom föreslog i sitt anbud. Avtal om ytterligare uppgifter för Eurokom, inklusive uppgifter i samband med införande av systemet i varje medlemsstat och projektets förvaltning, skall ingås i form av separata överenskommelser,
- anger följande taxa:
a) 300 ecu per år per lokal enhet enligt förteckningen i kommissionens beslut 92/175/EEG(6).
b) Överföringskostnader som skall variera med hänsyn till tillgång eller frånvaro av ett nationellt datacentrum och som motsvarar det fördelaktigaste pris som Eurokom har kunnat erhålla från leverantören av kommunikationsutrustning.
Artikel 3
Medlemsstaterna förpliktar sig att endast åberopa den uppsägningsklausul som avses i artikel 2 tredje strecksatsen enligt det förfarande som fastställs i artikel 20.3 i direktiv 90/425/EEG.
Artikel 4
Den sammanlagda årliga kostnaden för att delta i systemet som avses i artikel 2a femte strecksatsen och som inte skall överstiga det belopp som är fastställt för det första året, och dess fördelning mellan medlemsstaterna skall tas upp till förnyad prövning före den 1 juli 1993. Det maximala priset för varje medlemsstat under såväl det andra som tredje året skall dock inte öka med mer än 10 % av priset för det första året.
Artikel 5
Om det under införandet av systemet uppstår en situation som, särskilt vad gäller de ekonomiska aspekterna, inte ligger i linje med detta besluts mål, skall kommissionen vidta nödvändiga åtgärder i enlighet med förfarandet i artikel 42 i rådets beslut 90/424/EEG(7).
Artikel 6
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS DIREKTIV 92/4/EEG av den 10 februari 1992 om ändring i rådets direktiv 78/663/EEG om särskilda renhetskriterier för emulgerings-, stabiliserings-, förtjocknings- och geleringsmedel för användning i livsmedel
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 89/107/EEG av den 21 december 1988 om tillnärmning av medlemsstaternas lagstiftning om tillsatser som är godkända för användning i livsmedel(1), särskilt artikel 3.3 i detta, och med beaktande av följande:
Med hänsyn till de specifikationer som antagits genom Codex Alimentarius och till ny produktionsteknik är det nödvändigt att ändra rådets direktiv 78/663/EEG(2), senast ändrat genom kommissionens direktiv 90/612/EEG(3).
I enlighet med vad som föreskrivs i artikel 6 i direktiv 89/107/EEG har Vetenskapliga livsmedelskommittén rådfrågats om de föreskrifter som kan förväntas påverka folkhälsan.
De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga livsmedelskommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till direktiv 78/663/EEG ändras på det sätt som visas av bilagan till det här direktivet.
Artikel 2
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 juni 1993 och skall genast underrätta kommissionen om detta.
När en medlemsstat antar bestämmelser till följd av detta direktiv skall dessa innehålla en hänvisning till direktivet eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV 92/32/EEG av den 30 april 1992 om ändring för sjunde gången i rådets direktiv 67/548/EEG om tillnärmning av lagar och andra författningar om klassificering, förpackning och märkning av farliga ämnen
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag(1),
i samarbete med Europaparlamentet(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Olikheter mellan lagar och andra författningar om klassificering, förpackning och etikettering av farliga ämnen och anmälan av nya ämnen i medlemsstaterna kan leda till handelshinder mellan medlemsstater och skapa ojämlika konkurrensvillkor. Sådana skillnader mellan bestämmelserna i de olika medlemsstaterna påverkar direkt den inre marknadens funktion och har som följd att hälsa och miljö inte garanteras skydd på samma nivå.
Åtgärderna för en tillnärmning av de bestämmelser i medlemsstaterna som hänför sig till den inre marknadens upprättande och funktion skall, vad beträffar hälsan, säkerheten och skyddet för människan och miljön, utgå från en hög skyddsnivå.
För att skydda människan och miljön från potentiella risker som kan uppstå när nya ämnen släpps ut på marknaden är det nödvändigt att besluta om lämpliga åtgärder och särskilt att ändra och skärpa bestämmelserna i rådets direktiv 67/548/EEG(4) senast ändrat genom direktiv 90/517/EEG(5).
Alla nya ämnen som släpps ut på marknaden bör anmälas till de behöriga myndigheterna, varvid vissa uppgifter lämnas. Vad beträffar ämnen som släpps ut på marknaden i mindre kvantiteter än ett ton per år och tillverkare kan lägre krav ställas. Om å andra sidan ett ämne släpps ut på marknaden i kvantiteter som överstiger vissa gränser bör kompletterande undersökningar genomföras.
Bestämmelser bör fastställas för att införa ett anmälningsförfarande, varigenom en anmälan som gjorts i en medlemsstat gäller i hela gemenskapen. För ämnen som tillverkas utanför gemenskapen kan det vara lämpligt att tillverkaren utser en representant i gemenskapen som ensam svarar för anmälan.
För att kunna bedöma inverkan på människan och miljön bör ämnet göras till föremål för en riskbedömning. Enhetliga principer för denna riskbedömning bör fastställas.
Dessutom är det viktigt att noga följa utvecklingen och användningen av nya ämnen som släpps ut på marknaden. Det är därför nödvändigt att införa ett system varigenom alla nya ämnen tas upp i en förteckning.
Kommissionen har i enlighet med artikel 13.1 i direktiv 67/548/EEG(6) och enligt riktlinjer fastställda i kommissionens beslut 81/437/EEG gjort upp en förteckning över ämnen som fanns på marknaden i gemenskapen den 18 september 1981 (EINECS), vilken har publicerats i Europeiska gemenskapernas officiella tidning(7).
Enligt rådets direktiv 86/609/EEG av den 24 november 1986 om tillnärmning av medlemsstaternas lagar och andra författningar om skydd av djur som används för försök och andra vetenskapliga ändamål(8) är det önskvärt att nedbringa till ett minimum antalet djur som används i djurförsök. Alla lämpliga åtgärder bör vidtas för att undvika att redan gjorda djurförsök upprepas.
I rådets direktiv 87/18/EEG av den 18 december 1986 om harmonisering av lagar och andra författningar om tillämpningen av principerna för god laboratoriesed och kontrollen av och tillämpningen vid prov med kemiska ämnen(9) anges gemenskapens principer för god laboratoriesed, som skall följas vid tester av kemikalier.
För att stärka miljöskyddet och arbetarskyddet bör säkerhetsdatablad om farliga ämnen finnas tillgängliga för yrkesmässiga användare.
Till skydd för allmänheten och särskilt de arbetstagare som använder ämnena bör bestämmelser om klassificering och märkning av ämnen antas på gemenskapsnivå.
För att säkerställa en tillräckligt hög skyddsnivå för människan och miljön är det nödvändigt att vidta åtgärder som avser förpackning och provisorisk märkning av sådana farliga ämnen som inte finns upptagna i bilaga 1 till direktiv 67/548/EEG. Av samma anledning är det nödvändigt att göra tillhandahållandet av skyddsanvisningar obligatoriskt.
Enligt artikel 2 i direktiv 67/548/EEG klassificeras ämnen och preparat enligt allmänna definitioner som giftiga, hälsoskadliga, frätande eller irriterande. Erfarenheterna har visat att det är nödvändigt att förbättra denna klassificering. Exakta kriterier för klassificeringen bör anges. Enligt artikel 3 i direktivet skall också en bedömning göras av ämnets miljöfarlighet, vilket gör det nödvändigt att ange vissa kriterier och parametrar för bedömningen och införa ett undersökningsprogram i flera steg.
Det är önskvärt att införa ännu en farosymbol, "miljöfarligt", som skall anges på förpackningen.
Sekretess bör garanteras för vissa uppgifter om affärs- och driftförhållanden.
Medlemsstaterna bör i vissa fall tillåtas att vidta egna skyddsåtgärder.
Kommissionen bör ha befogenhet att anpassa samtliga bilagor till direktiv 67/548/EEG till den tekniska utvecklingen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 67/548/EEG ändras på följande sätt:
a) anmälan av ämnen,
b) utbyte av information om anmälda ämnen,
c) bedömning av de anmälda ämnenas potentiella risker för människan och miljön,
2. Direktivet skall inte gälla följande preparat i bruksfärdigt skick, avsedda för slutanvändaren:
a) Sådana farmaceutiska produkter för användning inom human- eller veterinärmedicin som avses i direktiv 65/65/EEG(1), senast ändrat genom direktiv 87/21/EEG(2).
b) Kosmetiska produkter som avses i direktiv 76/768/EEG(3), senast ändrat genom direktiv 86/199/EEG(4).
c) Ämnesblandningar som i form av avfall omfattas av direktiv 75/442/EEG(5) och 78/319/EEG(6).
d) Livsmedel.
e) Djurfoder.
f) Bekämpningsmedel.
g) Radioaktiva ämnen som avses i direktiv 80/836/EEG(7).
h) Andra ämnen eller preparat, för vilka tillämpas gemenskapsförfaranden för anmälan eller godkännande och för vilka kraven är likvärdiga med dem som föreskrivs i detta direktiv.
Kommissionen skall senast 12 månader efter anmälan av detta direktiv enligt förfarandet i artikel 29.4 a upprätta en förteckning över ovan nämnda ämnen och preparat. Förteckningen skall ses över regelbundet och vid behov ändras i enlighet med nämnda förfarande.
Detta direktiv skall inte heller gälla
- transport av farliga ämnen på järnväg, väg eller inre vattenväg, till sjöss eller med flyg,
Artikel 2
Definitioner
1. I detta direktiv används följande beteckningar med de betydelser som här anges:
a) ämnen: kemiska grundämnen och deras föreningar i naturlig eller framställd form, inklusive eventuella tillsatser nödvändiga för att bevara produkternas stabilitet och eventuella föroreningar som härrör från tillverkningsprocessen, men exklusive eventuella lösningsmedel som kan avskiljas utan att detta påverkar ämnets stabilitet eller ändrar dess sammansättning.
b) preparat: blandningar eller lösningar som består av två eller flera ämnen.
c) polymer: ett ämne bestående av molekyler, som kännetecknas av sammankoppling av en eller fler monomerenheter och utgörs av en enkel viktmajoritet molekyler som innehåller åtminstone tre monomerenheter kovalent bundna till åtminstone en annan monomerenhet eller annan reaktant, och som består av mindre än en enkel viktmajoritet molekyler med samma molekylvikt. Molekylerna skall vara fördelade över en rad molekylvikter, där skillnaden i molekylvikt främst kan hänföras till skillnader i antalet monomerenheter. I denna definition avses med "monomerenhet" en monomers form i en polymer efter reaktionen.
d) anmälan: de handlingar med föreskrivna uppgifter som lämnats till den behöriga myndigheten i en medlemsstat enligt följande:
- för ämnen framställda inom gemenskapen: av den tillverkare som släpper ut ett ämne på marknaden, ensamt eller i ett preparat,
e) släppa ut på marknaden: tillhandahållande till tredje part. I detta direktiv skall import till gemenskapens tullområde likställas med att släppa ut på marknaden.
f) vetenskaplig forskning och utveckling: vetenskapliga experiment, analyser eller kemisk forskning som utförs under kontrollerade förhållanden. Häri innefattas fastställandet av inneboende egenskaper, verkan och effektivitet såväl som vetenskapliga undersökningar i samband med produktutveckling.
g) processinriktad forskning och utveckling: vidareutvecklandet av ett ämne, varvid användningsområden för ämnet testas genom pilotförsök eller provtillverkning.
h) EINECS: (European Inventory of Existing Commercial Substances): Europeisk förteckning över befintliga marknadsförda ämnen. Denna lista utgör en fullständig förteckning över de ämnen som anses finnas på den gemensamma marknaden den 18 september 1981.
2. Med farliga avses i detta direktiv följande ämnen och preparat:
a) explosiva ämnen och preparat: fasta och flytande ämnen och ämnen i pasta- eller geléform som även utan närvaro av atmosfäriskt syre kan ge upphov till en exoterm reaktion och därvid snabbt avge gaser, och som under angivna testförhållanden detonerar, snabbt deflagrerar eller delvis inneslutna exploderar vid uppvärmning,
b) oxiderande ämnen och preparat: ämnen och preparat som i kontakt med andra ämnen, i synnerhet brandfarliga, ger upphov till en kraftig exoterm reaktion,
c) synnerligen brandfarliga ämnen och preparat: flytande ämnen och preparat som har ytterst låg flampunkt eller låg kokpunkt samt gasformiga ämnen och preparat som är antändbara i kontakt med luft av rumstemperatur och normalt lufttryck.
d) Mycket brandfarliga ämnen och preparat:
- ämnen och preparat som kan bli heta och slutligen fatta eld i kontakt med luft av rumstemperatur utan tillförsel av energi, eller
- fasta ämnen och preparat som lätt fattar eld även vid kortvarig kontakt med en antändningskälla och som fortsätter att brinna eller förbrukas även sedan kontakten med antändningskällan upphört, eller
- flytande ämnen och preparat med mycket låg flampunkt, eller
- ämnen och preparat som i kontakt med vatten eller fuktig luft utvecklar brandfarliga gaser i farliga mängder.
e) Brandfarliga ämnen och preparat: flytande ämnen och preparat med låg flampunkt.
f) Mycket giftiga ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden i mycket små mängder leder till döden eller ger akuta eller kroniska skador.
g) Giftiga ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden i små mängder leder till döden eller ger akuta eller kroniska skador.
h) Hälsoskadliga ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan leda till döden eller ge akuta eller kroniska skador.
i) Frätande ämnen och preparat: ämnen och preparat som vid kontakt med levande vävnader kan förstöra dessa.
j) Irriterande ämnen och preparat: ämnen och preparat som ej är frätande men som vid direkt, långvarig eller upprepad kontakt med hud eller slemhinnor kan orsaka inflammation.
k) Sensibiliserande ämnen och preparat: ämnen och preparat som vid inandning eller upptagning genom huden kan framkalla överkänslighet, så att karakteristiska symptom uppstår vid förnyad exponering för ämnet eller preparatet.
l) Cancerogena ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan orsaka eller öka förekomsten av cancer.
m) Mutagena ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan orsaka eller öka förekomsten av ärftliga genetiska defekter.
n) Ämnen och preparat skadliga för fortplantningen: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan orsaka eller öka förekomsten av icke ärftliga skador på avkomman eller på den manliga eller kvinnliga fortplantningsfunktionen eller -förmågan.
o) Miljöfarliga ämnen och preparat: ämnen och preparat som om de kommer ut i miljön utgör eller kan utgöra en omedelbar eller fördröjd fara för en eller flera delar av miljön.
Artikel 3
Tester och bedömning av ämnenas egenskaper
1. Tester på kemikalier som utförs inom ramen för detta direktiv skall som allmän princip utföras enligt de metoder som föreskrivs i bilaga 5. Ämnenas fysikaliskkemiska egenskaper skall bestämmas enligt de metoder som anges i bilaga 5 A. Deras toxicitet skall bestämmas enligt metoderna i bilaga 5 B och deras miljöfarlighet enligt metoderna i bilaga 5 C.
För vissa ämnen i EINECS kan det emellertid redan finnas existerande uppgifter som har tagits fram med andra metoder än de som förskrivs i bilaga 5. Huruvida dessa uppgifter är tillräckliga för att ämnet skall kunna klassificeras och märkas eller om produkten måste testas på nytt i enlighet med bilaga 5 avgörs från fall till fall, varvid bland annat beaktas att det är angeläget att begränsa antalet djurförsök med ryggradsdjur.
Laboratorieförsök skall utföras i enlighet med principerna för god laboratoriesed i direktiv 87/18/EEG och bestämmelserna i direktiv 86/609/EEG.
2. De verkliga och potentiella riskerna för människan och miljön skall bedömas enligt de principer som antagits den 30 april 1993 i enlighet med förfarandet i artikel 29.4 b. Dessa principer skall regelbundet ses över och vid behov ändras enligt samma förfarande.
Artikel 4
Klassificering
1. Ämnen skall klassificeras på grundval av sina inneboende egenskaper enligt de i artikel 2.2 fastställda kategorierna. Vid klassificering av ämnen skall hänsyn också tas till föroreningar, om dessa förekommer i koncentrationer som överstiger de koncentrationsgränser som anges i punkt 4 i denna artikel och i artikel 3 i direktiv 88/379/EEG.
2. De allmänna principerna för klassificering och märkning av ämnen och preparat skall tillämpas enligt kriterierna i bilaga 6(1), utom i fall då andra krav för farliga preparat anges i särskilda direktiv.
3. I bilaga 1(2) finns en förteckning över ämnen som klassificerats enligt principerna i punkt 1 och 2, med uppgift om deras harmoniserade klassificering och märkning. Beslutet att ta upp ett ämne i bilaga 1 med harmoniserad klassificering och märkning skall fattas enligt förfarandet i artikel 29.
Artikel 5
Medlemsstaternas förpliktelser
1. Om inte annat följer av artikel 13 skall medlemsstaterna vidta alla nödvändiga åtgärder för att säkerställa att ämnen inte kan släppas ut på marknaden, som sådana eller ingående i preparat, om de inte
- anmälts till den behöriga myndigheten i en av medlemsstaterna enligt detta direktiv,
- förpackats och märkts i enlighet med artikel 22-25, enligt kriterierna i bilaga 6 och i enlighet med resultaten av de tester som föreskrivs i bilaga 7 och 8, utom i fråga om preparat för vilka det finns särskilda bestämmelser i andra direktiv.
Dessutom skall medlemsstaterna vidta alla nödvändiga åtgärder för att säkerställa att bestämmelserna om säkerhetsdatablad i artikel 27 följs.
2. Bestämmelserna i andra strecksatsen i punkt 1 skall gälla tills ämnet upptas i bilaga 1 eller tills ett beslut att inte ta upp ämnet har fattats enligt förfarandet i artikel 29.
Artikel 6
Undersökningsplikt
Tillverkare, distributörer och importörer av i EINECS upptagna farliga ämnen som ännu inte finns med i bilaga 1 skall vara skyldiga att utföra en undersökning för att utröna vilka relevanta och tillgängliga data som finns om ämnenas egenskaper. Ämnena skall förpackas och provisoriskt märkas på grundval av denna information i enlighet med bestämmelserna i artikel 22-25 och enligt kriterierna i bilaga 6.
Artikel 7
Fullständig anmälan
1. Om inte annat följer av artikel 1.2, 8.1, 13 och 16.1 skall en anmälare av ett ämne lämna en anmälan till den behöriga myndighet som avses i artikel 16.1 i den medlemsstat där ämnet framställs eller, om tillverkaren befinner sig utanför gemenskapen, i den medlemsstat där anmälaren är verksam. Anmälan skall ha följande innehåll:
- En dokumentation med de uppgifter som krävs för att bedöma de förutsebara risker, såväl omedelbara som fördröjda, som ämnet kan medföra för människan och miljön, tillsammans med all tillgänglig information som är relevant för en sådan bedömning. Som ett minimum skall ingå de uppgifter och de undersökningsresultat som avses i bilaga 7 A, tillsammans med en detaljerad och fullständig beskrivning av de företagna undersökningarna och av de metoder som använts eller litteraturreferenser till dem.
- En redovisning av ämnets negativa effekter inom olika tänkbara användningsområden.
- Föreslagen klassificering och märkning av ämnet enligt detta direktiv.
- Endast beträffande farliga ämnen, ett förslag till säkerhetsdatablad enligt artikel 27.
- Om tillverkaren befinner sig utanför gemenskapen skall anmälaren, i enlighet med artikel 2.1 d andra strecksatsen, vid behov bifoga en förklaring från tillverkaren att anmälaren har utsetts att ensam företräda tillverkaren när det gäller att inge anmälan för ämnet i fråga.
- Anmälaren kan, om han så önskar, bifoga en motiverad begäran om att bestämmelserna i artikel 15.2 inte skall tillämpas i fråga om anmälan under en tidsperiod som inte i något fall får överstiga ett år från tidpunkten för anmälan.
Utöver ovan nämnda uppgifter kan anmälaren också tillhandahålla en preliminär riskbedömning som han gjort i enlighet med principerna i artikel 3.2.
2. Om inte annat följer av artikel 14 skall varje anmälare av ett redan anmält ämne underrätta den behöriga myndigheten
- när den mängd av ämnet som släppts ut på marknaden uppnår 10 ton per år och tillverkare, eller när den totala mängd av ämnet som släppts ut på marknaden uppnår 50 ton per tillverkare, varvid den behöriga myndigheten kan kräva att en del eller samtliga kompletterande tester/undersökningar som föreskrivs i bilaga 8 nivå 1 skall utföras inom den tid som den behöriga myndigheten bestämmer,
- när den mängd av ämnet som släppts ut på marknaden uppnår 100 ton per år och tillverkare, eller när den totala mängd av ämnet som släppts ut på marknaden uppnår 500 ton per tillverkare, varvid den behöriga myndigheten skall kräva att de kompletterande tester/undersökningar som föreskrivs i bilaga 8 nivå 1 skall utföras inom den tid som den behöriga myndigheten bestämmer, utom i fall då anmälaren kan visa att en viss test/undersökning är olämplig eller att en alternativ test/undersökning är att föredra,
- när den mängd av ämnet som släppts ut på marknaden uppnår 1000 ton per år och tillverkare, eller när den totala mängd av ämnet som släppts ut på marknaden uppnår 5000 ton per tillverkare, varvid den behöriga myndigheten skall lägga upp ett program för tester/undersökningar enligt bilaga 8 nivå 2, som skall genomföras av anmälaren inom den tid som den behöriga myndigheten bestämmer.
3. När kompletterande tester utförs, i enlighet med kraven i punkt 2 eller frivilligt, skall anmälaren meddela resultaten till den behöriga myndigheten.
Artikel 8
Begränsade anmälningskrav för ämnen som släpps ut på marknaden i mängder under ett ton per år och tillverkare
1. Om inte annat följer av artikel 1.2, 13.1 och 16.1 skall en anmälare som avser att släppa ut ett ämne på marknaden inom gemenskapen i mängder som understiger ett ton per år och tillverkare vara skyldig att till den behöriga myndighet som avses i artikel 16.1 i den medlemsstat där ämnet framställs eller, om tillverkaren befinner sig utanför gemenskapen, i den medlemsstat där anmälaren är verksam, lämna en anmälan med följande innehåll:
- En dokumentation med de uppgifter som krävs för en bedömning av de förutsebara risker, såväl omedelbara som fördröjda, som ämnet kan medföra för människan och miljön, tillsammans med all tillgänglig information som är relevant för en sådan bedömning. Som ett minimum skall i dokumentationen ingå de uppgifter och de undersökningsresultat som avses i bilaga 7 B, tillsammans med en detaljerad och fullständig beskrivning av de företagna undersökningarna och av de metoder som använts eller litteraturreferenser till dem, om den medlemsstat där anmälan lämnas så kräver.
- Alla övriga uppgifter enligt artikel 7.1.
2. Om mängden som släpps ut på marknaden understiger 100 kg per år och tillverkare kan anmälaren, om inte annat följer av artikel 16.1, begränsa uppgifterna i den ovannämnda dokumentationen till vad som föreskrivs i bilaga 7 C.
3. Om en anmälare har lämnat en begränsad dokumentation enligt punkt 2, skall han, innan den mängd av ämnet som släpps ut på marknaden uppnår 100 kg per år och tillverkare eller den totala mängd som släpps ut på marknaden per tillverkare uppnår 500 kg, förse den behöriga myndigheten med de kompletterande uppgifter som krävs för att rapporten skall motsvara kraven i bilaga 7 B.
4. Likaledes skall en anmälare som har lämnat en begränsad anmälan enligt kraven i punkt 1, lämna en fullständig anmälan enligt kraven i artikel 7 innan den mängd av ämnet som släpps ut på marknaden uppnår ett ton per år per tillverkare eller den totala mängd som släpps ut på marknaden per tillverkare uppnår fem ton
5. De ämnen som anmälts enligt punkt 1 och 2 skall, i den mån anmälaren rimligen kan förväntas känna till deras farliga egenskaper, förpackas och provisoriskt märkas i enlighet med reglerna i artikel 22-25 och enligt kriterierna i bilaga 6. Om det ännu inte är möjligt att märka dem i enlighet med principerna i artikel 23, skall utöver märkningen från de redan utförda testerna på etiketten anges "Varning - ämnet ännu inte fullständigt testat".
Artikel 9
Redan anmälda ämnen (tioårsregeln)
Om uppgifter enligt artikel 7 och 8 lämnats minst 10 år tidigare behöver en anmälare inte tillhandahålla sådana uppgifter som krävs för dokumentationen enligt bilaga 7 A 7 D, förutom uppgifterna under punkt 1 och 2 i de nämnda bilagorna.
Artikel 10
Utsläppande på marknaden av anmälda ämnen
1. Om inte annat anges av den behöriga myndigheten, får ämnen som anmälts enligt artikel 7.1 släppas ut på marknaden tidigast 60 dagar efter det att myndigheten mottagit en dokumentation som överensstämmer med kraven i detta direktiv.
Om den behöriga myndigheten anser att dokumentationen inte uppfyller kraven i direktivet och meddelar anmälaren detta enligt artikel 16.2, får ämnet släppas ut på marknaden tidigast 60 dagar efter det att myndigheten mottagit de uppgifter som behövs för att anmälan skall överensstämma med direktivet.
2. Om inte annat anges av den behöriga myndigheten, får ämnen som anmälts enligt artikel 8.1 eller 8.2 släppas ut på marknaden tidigast 30 dagar efter det att myndigheten mottagit en dokumentation som överensstämmer med kraven i detta direktiv.
Om den behöriga myndigheten anser att dokumentationen inte uppfyller kraven i direktivet och meddelar anmälaren detta enligt artikel 16.3, får ämnet släppas ut på marknaden tidigast 30 dagar efter det att myndigheten mottagit de uppgifter som behövs för att anmälan skall överensstämma med direktivets krav. Om anmälaren underrättats enligt artikel 16.3 att dokumentationen har godtagits, gäller dock att ämnet får släppas ut på marknaden tidigast 15 dagar efter det att den behöriga myndigheten mottagit dokumentationen.
Artikel 11
Ämnen som framställs utanför gemenskapen
Om det i fråga om ämnen som framställs utanför gemenskapen finns mer än en anmälan för ett ämne framställt av samma tillverkare, skall kommissionen och de nationella myndigheterna fastställa den totala årliga mängden som släpps ut på marknaden inom gemenskapen på grundval av de uppgifter som lämnats enligt artikel 7.1, 8.1 och 14. Skyldigheten att utföra kompletterande tester enligt artikel 7.2 åligger samtliga anmälare gemensamt.
Artikel 12
Polymerer
I fråga om polymerer skall särskilda bestämmelser fastställas i bilaga 7 i den form som anges i bilaga 7 D och enligt det förfarande som anges i artikel 29.4 b angående den dokumentation som enligt artikel 7.1 och 8.1 skall ingå i anmälan.
Artikel 13
Undantagsbestämmelser
1. Bestämmelserna i artikel 7, 8, 14 och 15 tillämpas inte på följande ämnen:
- Ämnen som finns upptagna i EINECS.
- Tillsatser och ämnen som endast används i djurfoder och omfattas av direktiv 70/524/EEG och 82/471/EEG(1).
- Ämnen som endast används i livsmedel och omfattas av direktiv 89/107/EEG(2), samt ämnen som endast används som smakämnen i livsmedel och omfattas av direktiv 88/388/EEG.
- Aktiva ingredienser som endast används i de farmaceutiska produkter som avses i artikel 1.2 a. Som sådana räknas inte kemiska halvfabrikat.
- Ämnen som endast används i vissa andra produktkategorier för vilka gemenskapen tillämpar anmälnings- eller godkännandeförfaranden och för vilka kraven i fråga om uppgiftslämnande är likvärdiga med dem som föreskrivs i detta direktiv. Senast 12 månader efter anmälan av detta direktiv skall kommissionen i enlighet med förfarandet i artikel 29.4 a upprätta en förteckning över sådana gemenskapsregler. Denna förteckning skall regelbundet ses över och vid behov ändras enligt samma förfarande.
2. De ämnen som anges nedan skall anses ha anmälts enligt detta direktiv om följande villkor är uppfyllda:
- Polymerer med undantag för sådana som i kombinerad form innehåller minst 2 % av ett ämne som inte finns upptaget i EINECS.
- Ämnen som släpps ut på marknaden i mindre mängder än 10 kg per år och tillverkare, förutsatt att tillverkaren/importören uppfyller de krav som uppställs av de medlemsstater där ämnet släpps ut på marknaden. Dessa krav får inte gå utöver vad som föreskrivs i bilaga 7 C, punkt 1 och 2.
- Ämnen som släpps ut på marknaden i begränsade mängder, inte i något fall över 100 kg per tillverkare och år, och som är avsedda enbart för vetenskaplig forskning och utveckling som utförs under kontrollerade förhållanden.
En tillverkare eller importör som begagnar sig av detta undantag måste föra löpande anteckningar av vilka framgår ämnets identitet, märkningsinformation, mängder samt en förteckning över kunder. Dessa uppgifter skall på begäran ställas till förfogande för den behöriga myndigheten i den medlemsstat där tillverkningen, importen eller den vetenskapliga forskningen och utvecklingen sker.
- Ämnen som säljs till ett begränsat antal registrerade kunder för användning vid processinriktad forskning och utveckling i mängder som är begränsade till vad som krävs för den processinriktade forskningen och utvecklingen. Dessa ämnen får undantas i ett år, under förutsättning dels att tillverkaren eller importören till den behöriga myndigheten i varje medlemsstat där tillverkning, import eller processinriktad forskning och utveckling sker lämnar uppgifter om ämnenas identitet, märkningsinformation, mängder, skälen varför dessa mängder behövs samt en förteckning över kunderna och deras forsknings- och utvecklingsprogram, dels att han rättar sig efter krav som dessa myndigheter eller medlemsstaterna uppställer för sådan forskning och utveckling. De krav som medlemsstaterna uppställer får inte gå utöver vad som föreskrivs i artikel 8. Efter ett år skall anmälningsskyldighet normalt gälla för dessa ämnen. Tillverkaren eller importören skall också försäkra att ämnet eller preparatet det ingår i endast kommer att hanteras av kundens personal under kontrollerade förhållanden och inte vid något tillfälle kommer att göras tillgängligt för allmänheten, som sådant eller i ett preparat. Om den behöriga myndigheten anser att en oacceptabel risk föreligger för människan eller miljön kan myndigheten vidare föreskriva att detsamma skall gälla för produkter som innehåller de nya ämnen som framställts under den processinriktade forskningen och utvecklingen.
I undantagsfall får den ovannämnda ettårsperioden förlängas med ytterligare ett år, om anmälaren på ett tillfredsställande sätt kan visa för den behöriga myndigheten att en sådan förlängning är motiverad.
3. De ämnen som avses i punkt 2 skall, i den mån anmälaren rimligen kan förväntas känna till deras farliga egenskaper, förpackas och provisoriskt märkas av tillverkaren eller dennes representant i enlighet med reglerna i artikel 22-25 och enligt kriterierna i bilaga 6.
Om det inte är möjligt att märka ämnena fullständigt och i enlighet med principerna i artikel 23 på grund av att resultaten från testerna enligt bilaga 7 A inte är tillgängliga, bör utöver märkningen från de utförda testerna på etiketten anges "Varning - ämnet ännu inte fullständigt testat".
Artikel 14
Kompletterande uppgifter
1. En anmälare av ett ämne som redan anmälts i enlighet med artikel 7.1 eller 8.1 skall vara skyldig att på eget initiativ skriftligen underrätta den behöriga myndighet till vilken anmälan ursprungligen lämnades om:
- förändringar i de årliga eller totala mängder som släpps ut på den gemensamma marknaden av honom eller, om ämnet tillverkas utanför gemenskapen och anmälaren ensam företräder denne, av honom eller någon annan,
- nya rön angående ämnets påverkan på människan eller miljön, som han rimligen kan förväntas känna till,
- nya användningsområden för vilka ämnet släpps ut på marknaden och som han rimligen kan förväntas känna till,
- alla ändringar i ämnenas sammansättning som avses i bilaga 7 A, B eller C, avsnitt 1.3,
- alla förändringar i hans ställning (tillverkare eller importör).
2. Varje importör av ett ämne framställt av en tillverkare utanför gemenskapen som importerar ämnet inom ramen för en anmälan som tidigare lämnats av en ensam företrädare i enlighet med artikel 2.1 d, skall vara skyldig att tillse att denne förses med aktuell information angående de mängder av ämnet som han släpper ut på marknaden inom gemenskapen.
Artikel 15
Ny anmälan av samma ämne och åtgärder för att undvika upprepade tester på ryggradsdjur
1. För ett ämne som redan har anmälts i enlighet med artikel 7.1 eller 8.1, kan den behöriga myndigheten medge att den som därefter anmäler ämnet vid tillämpningen av avsnitt 3-5 i bilaga 7 A och B och avsnitt 3 och 4 i bilaga 7 c åberopar de testresultat som lämnats av den förste anmälaren, förutsatt att den andre anmälaren kan visa att det nyanmälda ämnet är identiskt med det redan anmälda, också vad beträffar renhetsgrad och föroreningar. Den förste anmälaren måste ge skriftligt tillstånd till att hans testresultat får åberopas.
2. Innan försök utförs på ryggradsdjur i syfte att upprätta en anmälan i enlighet med artikel 7.1 eller 8.1, och om inte annat följer av punkt 1, skall den som avser att anmäla ett ämne fråga den behöriga myndigheten i den medlemsstat där han ämnar inlämna sin anmälan
a) om det ämne han avser att anmäla redan är anmält, och
b) om den första anmälarens namn och adress.
a) Den behöriga myndighet som mottar förfrågan finner det styrkt att den nya anmälaren ämnar släppa ut ämnet på marknaden i de uppgivna mängderna.
b) Ämnet är tidigare anmält.
c) Den första anmälaren har inte begärt och beviljats ett tidsbegränsat undantag från denna artikel.
Den första anmälaren och den nya anmälaren skall vidta alla rimliga åtgärder för att nå en överenskommelse om utbyte av information, så att upprepade tester på ryggradsdjur kan undvikas.
3. Anmälare av ett ämne som i enlighet med punkt 1 och 2 har kommit överens om utbyte av information enligt bilaga 7 skall också vidta alla nödvändiga åtgärder för att nå en överenskommelse om utbyte av information som erhållits från tester på ryggradsdjur och som lämnats i enlighet med artikel 7.2.
4. Om en anmälare och en ny anmälare av ett och samma ämne trots bestämmelserna i punkt 2 och 3 inte kan nå en överenskommelse om utbyte av information, får medlemsstaterna, i syfte att förhindra tester på ryggradsdjur, i fråga om anmälare inom deras territorier tillämpa nationella bestämmelser, som innebär att gamla och nya anmälare är skyldiga att dela på uppgiftslämnandet, och fastställa förfarandet för användningen av uppgifterna. Bestämmelserna får omfatta regler om det tidsbegränsade undantag som avses i artikel 7.1 sista strecksatsen och om en rimlig avvägning mellan berörda parters intressen.
Artikel 16
Myndigheternas rättigheter och skyldigheter
1. Medlemsstaterna skall utse en eller flera behöriga myndigheter som skall ansvara för mottagandet av uppgifter enligt artikel 7-14 och för bedömningen av huruvida uppgifterna överensstämmer med kraven i detta direktiv.
Om det visar sig nödvändigt för bedömningen av riskerna med ett ämne får de behöriga myndigheterna dessutom begära ytterligare underlag eller kompletterande tester angående ämnen eller nedbrytningsprodukter som har anmälts eller beträffande vilka uppgifter lämnats enligt detta direktiv. Därvid kan begäras att sådana uppgifter som avses i bilaga 8 skall lämnas tidigare än som anges i artikel 7.2.
Dessutom får de behöriga myndigheterna
- i kontrollsyfte ta nödvändiga prover,
- begära att anmälaren tillhandahåller ämnet i sådana mängder som anses nödvändiga för att utöva kontrolltester,
- vidta lämpliga åtgärder som hänför sig till en säker användning av ämnet, tills sådana bestämmelser införs på gemenskapsnivå.
I fråga om ämnen som anmälts i enlighet med artikel 7.1, 8.1 och 8.2 skall den behöriga myndighet som mottar anmälan göra en riskbedömning i enlighet med de allmänna principer som avses i artikel 3.2. Bedömningen skall omfatta rekommendationer om den lämpligaste metoden för att testa ämnet och, där så är lämpligt, rekommendationer om åtgärder i syfte att minska riskerna för människan och miljön i samband med att ämnet släpps ut på marknaden. Riskbedömningen skall regelbundet ses över med hänsyn till kompletterande uppgifter som lämnas i enlighet med denna artikel eller artikel 7.2, 8.3 och 14.1.
2. I fråga om anmälningar som lämnats i enlighet med artikel 7 skall myndigheterna inom 60 dagar efter mottagandet skriftligen underrätta anmälaren om huruvida anmälan anses överensstämma med detta direktiv.
Om dokumentationen godtas skall myndigheten samtidigt meddela anmälaren det officiella nummer som tilldelats hans anmälan. Om dokumentationen inte godtas skall myndigheten meddela anmälaren vilka kompletterande uppgifter som krävs för att dokumentationen skall anses överensstämma med detta direktiv.
3. I fråga om anmälningar som lämnats i enlighet med artikel 8 skall de behöriga myndigheterna senast 30 dagar efter det att anmälan kommit in avgöra om den överensstämmer med detta direktiv och, i fall då anmälan bedöms inte överensstämma med detta direktiv, upplysa anmälaren om vilka kompletterande uppgifter som krävs för att dokumentationen skall överensstämma med direktivet. Om anmälan överensstämmer med detta direktiv skall myndigheten inom samma tid meddela anmälaren det officiella nummer som tilldelats hans anmälan.
4. Beträffande ämnen som framställts utanför gemenskapen och för vilka fler än en anmälan inkommit som avser ett ämne som framställs av en och samma tillverkare, skall de behöriga myndigheterna tillsammans med kommissionen svara för beräkningen av de årliga och totala mängder som släpps ut på marknaden inom gemenskapen. Om de mängder uppnås som anges i artikel 7.2, skall den behöriga myndighet som mottagit anmälan eller anmälningarna kontakta anmälarna, meddela dem vilka de andra anmälarna är och upplysa dem om deras gemensamma ansvar enligt artikel 11.
5. Förfarandet i artikel 28 skall följas när ett förslag till klassificering och märkning fastställs eller ändras.
6. Om inte annat följer av artikel 19.1 skall medlemsstaterna och kommissionen tillse att sekretess gäller för uppgifter om kommersiell utveckling och tillverkning.
Artikel 17
Kommissionens roll i anmälningsförfarandet
När en medlemsstat mottagit den dokumentation som avses i artikel 7.1 och 8.1 eller uppgifter från kompletterande tester som utförts enligt artikel 7.2 och 8.3 eller kompletterande uppgifter som lämnats i enlighet med artikel 14, skall den till kommissionen snarast möjligt sända en kopia av dokumentationen eller av de kompletterande uppgifterna eller en sammanfattning därav.
I fråga om de kompletterande uppgifter som avses i artikel 16.1 skall den behöriga myndigheten meddela kommissionen vilka tester som valts, skälen för detta, testresultaten och, i tillämpliga fall, bedömningen av resultaten. I fråga om uppgifter som mottagits i enlighet med artikel 13.2 skall den behöriga myndigheten till kommissionen vidarebefordra sådana som kan vara av allmänt intresse för kommissionen och andra behöriga myndigheter.
Den riskbedömning som avses i artikel 16.1 eller en sammanfattning av denna bedömning skall vidarebefordras till kommissionen så snart den är tillgänglig.
Artikel 18
Kommissionens skyldigheter
1. När dokumentation och de uppgifter som avses i artikel 17 kommit in till kommissionen skall den vidarebefordra kopior till medlemsstaterna. Kommissionen kan också om den anser det lämpligt vidarebefordra annat relevant material som den har insamlat i enlighet med detta direktiv.
2. En behörig myndighet i en annan medlemsstat kan direkt samråda med den behöriga myndighet som mottog den ursprungliga anmälan eller med kommissionen om vissa punkter i de uppgifter som ingår i den dokumentation som föreskrivs i detta direktiv eller om den riskbedömning som avses i artikel 16.1. Den kan också föreslå att ytterligare tester eller uppgifter begärs eller att riskbedömningen omprövas. Om den behöriga myndighet som mottog den ursprungliga anmälan inte tillmötesgår de andra myndigheternas önskemål rörande kompletterande uppgifter, bekräftande tester eller ändringar av de undersökningsprogram som avses i bilaga 8, eller rörande riskbedömningen, skall den motivera sitt beslut för de berörda myndigheterna. Om myndigheterna inte kan enas och någon av myndigheterna med stöd av utförligt angivna skäl finner att kompletterande uppgifter, bekräftande tester, ändringar av undersökningsprogrammen eller en omprövning av riskerna verkligen krävs för att skydda människan och miljön, kan den begära att kommissionen fattar ett beslut i enlighet med förfarandet i artikel 29.4 b.
Artikel 19
Sekretess
1. Om anmälaren anser att det finns ett sekretessproblem, kan han ange vilka uppgifter enligt artikel 7, 8 och 14 som enligt hans bedömning är kommersiellt känsliga och kan medföra skada industriellt eller kommersiellt om de lämnas ut, och som därför bör hållas hemliga för alla utom för de behöriga myndigheterna och kommissionen. En fullständig motivering måste lämnas i sådana fall.
I fråga om anmälningar och uppgifter som lämnats i enlighet med artikel 7.1, 7.2 och 7.3, samt skall industriell och kommersiell sekretess inte gälla för
a) ämnets handelsnamn,
b) tillverkarens eller anmälarens namn,
c) fysikalisk-kemiska uppgifter om ämnet enligt avsnitt 3 i bilaga 7 A 7 C,
d) möjliga sätt att göra ämnet ofarligt,
e) sammanfattningen av resultaten från toxikologiska och ekotoxikologiska tester,
h) informationen som lämnas i säkerhetsdatabladet,
i) vad gäller ämnen i bilaga 1, analysmetoder som gör det möjligt att upptäcka ett farligt ämne när det kommit ut i miljön och bestämma direkt exponering hos människor.
Om anmälaren, tillverkaren eller importören själv senare offentliggör tidigare sekretessbelagda uppgifter, skall han meddela den behöriga myndigheten detta.
2. Den myndighet som mottagit anmälan eller uppgifterna skall på eget ansvar avgöra vilka uppgifter som omfattas av industriell och kommersiell sekretess i enlighet med punkt 1.
Uppgifter som godtagits som konfidentiella av den myndighet som mottagit anmälningshandlingarna från anmälaren skall behandlas som konfidentiella även av andra behöriga myndigheter och av kommissionen.
3. Ämnen som finns upptagna i förteckningen enligt artikel 21.1 och som inte är klassificerade som farliga i detta direktivs mening kan, om den behöriga myndighet som mottagit anmälan så begär, upptas under sitt handelsnamn. Normalt får sådana ämnen upptas under handelsnamnet i högst tre år. Om den behöriga myndighet som mottog anmälan anser att ett offentliggörande av det kemiska namnet i dess IUPAC-form i sig självt skulle avslöja information angående kommersiellt utnyttjande eller kommersiell framställning, kan ämnet emellertid upptas under sitt handelsnamn så länge den behöriga myndigheten anser det lämpligt.
Farliga ämnen kan på begäran från den behöriga myndighet som mottog anmälan upptas endast under sina handelsnamn tills de upptas i bilaga 1.
4. Sekretessbelagda uppgifter som kommer till kommissionens eller en medlemsstats kännedom skall hållas hemliga.
I samtliga fall gäller att sådana uppgifter
- får lämnas ut endast till de myndigheter vilkas ansvars områden anges i artikel 16.1,
- dock får röjas för sådana personer som är direkt engagerade i administrativa eller rättsliga förfaranden som innefattar sanktioner och som genomförs i syfte att kontrollera ämnen som släppts ut på marknaden, samt för personer som deltar i eller skall höras i samband med lagstiftningsarbete.
Artikel 20
Utväxling av den sammanfattade dokumentationen
1. De uppgifter som lämnats i enlighet med artikel 17 och 18.1 kan vidarebefordras till kommissionen och medlemsstaterna i sammanfattad form.
I sådana fall skall de behöriga myndigheterna i en medlemsstat och kommissionen för tillämpningen av artikel 18.2 alltid kunna ta del av anmälningshandlingarna och de kompletterande uppgifterna.
2. Kommissionen skall utforma ett gemensamt system för utväxling av de uppgifter som avses i artikel 17 och 18.1. Detta system skall antas enligt förfarandet i artikel 29.
Artikel 21
Förteckningar över existerande och nya ämnen
1. Kommissionen skall upprätta en förteckning över samtliga ämnen som anmälts enligt detta direktiv. Listan skall sammanställas i enlighet med bestämmelserna i kommissionens beslut 85/71/EEG(1).
Artikel 22
Förpackning
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att tillse att farliga ämnen endast kan släppas ut på marknaden om förpackningen uppfyller följande krav:
a) Förpackningen skall vara så utformad och konstruerad att allt läckage förhindras. Detta krav skall inte gälla om särskilda säkerhetsanordningar föreskrivs.
b) Materialet i förpackningen och förslutningen skall inte kunna angripas av innehållet eller bilda farliga föreningar med detta.
c) Förpackningen och förslutningarna skall genomgående vara starka och stadiga så att de inte kan lossna och så att de tål normal påfrestning under hanteringen.
d) Återförslutbara stängningsanordningar skall vara så konstruerade att de kan återförslutas upprepade gånger utan att innehållet kan komma ut.
e) Behållare som innehåller ämnen som säljs till eller tillhandahålls allmänheten och är märkta "mycket giftigt", "giftigt" eller "frätande" enligt detta direktiv skall, oberoende av storleken, vara försedda med barnsäkra förslutningsanordningar och en varningsmärkning som kan uppfattas vid beröring.
f) Behållare som innehåller ämnen som säljs till eller tillhandahålls allmänheten och är märkta "hälsoskadligt", "synnerligen brandfarligt" eller "mycket brandfarligt" enligt detta direktiv skall, oberoende av storleken, vara försedda med en varningsmärkning som kan uppfattas vid beröring.
2. Medlemsstaterna kan också föreskriva att förpackningarna ursprungligen skall vara förslutna och plomberade på ett sådant sätt att plomberingen bryts när förpackningen öppnas första gången.
3. Ändringar i de kategorier av ämnen vilkas förpackningar skall vara utrustade enligt punkt 1 e och 1 f skall beslutas enligt förfarandet i artikel 29.
4. Ändringar i de tekniska specifikationerna för de anordningar som avses i punkt 1 e och 1 f skall beslutas enligt förfarandet i artikel 29.4 och återfinns i punkt A och B i bilaga 9 till detta direktiv.
Artikel 23
Märkning
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att säkerställa att farliga ämnen endast släpps ut på marknaden om märkningen på förpackningen uppfyller följande krav.
2. På varje förpackning skall tydligt och outplånligt anges följande:
a) Namnet på ämnet enligt en av de benämningar som anges i bilaga 1. Om ämnet ännu inte är upptaget i bilaga 1 skall namnet anges med den internationellt vedertagna nomenklaturen.
b) Namn och fullständig adress med telefonnummer för den i gemenskapen verksamma person som är ansvarig för att ämnet släpps ut på marknaden, antingen denne är tillverkare, importör eller distributör.
c) Farosymboler, om sådana fastställts, och upplysning om typen av fara som är förenad med ämnets användning. Farosymbolens utformning och ordalydelsen i faroangivelsen skall följa vad som föreskrivs i bilaga 2(1). Symbolen skall vara tryckt i svart på orangegul botten. Farosymboler och faroangivelser skall överensstämma med dem som anges i bilaga 1. För farliga ämnen som ännu inte finns upptagna i bilaga 1 skall faroangivelser och farobeteckningar tilldelas enligt reglerna i bilaga 6.
Om mer än en farosymbol tilldelas ett ämne gäller följande:
- Om symbolen T är obligatorisk behöver inte symbolerna X och C anges, om inte annat följer av bilaga 1.
- Om symbolen C är obligatorisk behöver inte symbolen X anges.
- Om symbolen E är obligatorisk behöver inte symbolerna F och O anges.
d) Standardfraser (R-fraser) som anger särskilda risker som är förenade med användningen av ämnet. R-fraserna skall överensstämma med vad som anges i bilaga 3. De R-fraser som skall användas för varje ämne anges i bilaga 1. För farliga ämnen som ännu inte finns upptagna i bilaga 1 skall R-fraser tilldelas enligt reglerna i bilaga 6.
e) Standardfraser (S-fraser) med skyddsanvisningar för en säker användning av ämnet. S-fraserna skall överensstämma med vad som anges i bilaga 4. De S-fraser som skall användas för varje ämne anges i bilaga 1. För farliga ämnen som ännu inte finns upptagna i bilaga 1 skall S-fraser tilldelas enligt reglerna i bilaga 6.
f) EEG-nummer, när sådant tilldelats. EEG-numret erhålls från EINECS eller från den förteckning som avses i artikel 21.1.
För ämnen som finns upptagna i bilaga 1 skall dessutom ordet "EEG-märkning" anges på etiketten.
3. För irriterande, mycket brandfarliga, brandfarliga och oxiderande ämnen behöver R-fraser och S-fraser inte anges om förpackningen inte innehåller mer än 125 ml. Detta gäller också för samma mängd farliga ämnen som inte säljs av detaljister till allmänheten.
4. Information av typen "inte giftig", "inte hälsoskadlig" eller annan liknande upplysning får inte förekomma på etiketter eller förpackningar till ämnen som omfattas av detta direktiv.
Artikel 24
Tillämpningen av märkningskraven
Dessa mått är endast avsedda för den information som krävs enligt detta direktiv och vid behov för kompletterande hälso- och säkerhetsinformation.
2. Etikett krävs inte om uppgifterna är tydligt angivna på själva förpackningen i enlighet med punkt 1.
3. Etiketten - eller i fall som avses i punkt 2, förpackningen - skall ha sådan färg och utformning att farosymbolen och dess bakgrund framträder tydligt.
4. De i artikel 23 föreskrivna upplysningarna på etiketten skall framträda tydligt mot bakgrunden och skall vara tryckta i så stor stil och med så stora mellanrum att de är lätta att läsa.
Särskilda bestämmelser om de upplysningarna som avser utformning och dimensioner förs in i bilaga 6 enligt förfarandet i artikel 29.4 b.
5. Medlemsstaterna får föreskriva att farliga ämnen som släpps ut på marknaden i det egna landet skall vara märkta på landets eget eller egna språk.
6. Vid tillämpningen av detta direktiv skall märkningskraven anses vara uppfyllda i följande fall:
a) När en yttre förpackning innehåller en eller flera inre förpackningar, om den yttre förpackningen är märkt enligt internationella regler för transport av farliga ämnen och den inre förpackningen eller de inre förpackningarna är märkta i enlighet med detta direktiv.
b) När det bara finns en förpackning
- och denna förpackning är märkt i enlighet med internationella regler om transport av farliga ämnen och enligt artikel 23.2 a, b och d-f, och
- när det behövs för särskilda typer av förpackningar såsom transportabla gasflaskor, förpackningen är märkt i enlighet med de särskilda krav som anges i bilaga 6.
För farliga ämnen som inte lämnar en medlemsstats territorium får märkning ske enligt nationella regler i stället för enligt internationella regler för transport av farliga ämnen.
Artikel 25
Undantag från kraven på märkning och förpackning
1. Artikel 22-24 skall inte gälla sådana bestämmelser som avser ammunition eller explosiva varor som släpps ut på marknaden för att vid användningen ge explosioner eller pyrotekniska effekter.
Ovannämnda artiklar skall inte heller gälla bestämmelser som avser butan, propan eller gasol förrän den 30 april 1997.
2. Dessutom får medlemsstaterna
a) tillåta att märkning enligt artikel 23 anbringas på annat lämpligt sätt om förpackningen är för liten eller på annat sätt olämplig för att märkas i enlighet med artikel 24.1 och 24.2,
b) trots bestämmelserna i artikel 23 och 24 tillåta att förpackningen för farliga ämnen som inte är explosiva, mycket giftiga eller giftiga förpackas omärkta eller märks på något annat sätt, om de innehåller så små mängder att det inte finns någon anledning anta att de som hanterar ämnet eller andra kan utsättas för fara,
c) om förpackningen är för liten för märkning enligt artikel 23 och 24 och det inte finns någon anledning att anta att de som hanterar ämnet eller andra kan utsättas för fara, trots bestämmelserna i ovanstående artiklar tillåta att förpackningar med explosiva, mycket giftiga eller giftiga ämnen märks på annat lämpligt sätt.
Detta undantag innebär inte att andra symboler, faroangivelser, R-fraser eller S-fraser än dem som föreskrivs i detta direktiv får användas.
3. Om en medlemsstat tillämpar något av undantagen i punkt 2 skall den genast underrätta kommissionen.
Artikel 26
Reklam
Reklam för ett ämne som tillhör en eller flera av kategorierna i artikel 2.2 skall vara förbjuden om inte de aktuella kategorierna anges i reklamen.
Artikel 27
Säkerhetsdatablad
1. För att särskilt yrkesmässiga användare skall kunna vidta nödvändiga åtgärder till skydd för miljön samt hälsan och säkerheten på arbetsplatsen skall tillverkaren, importören eller distributören i samband med eller före den första leveransen lämna ett säkerhetsdatablad till mottagaren. Detta blad skall innehålla den information som krävs för att skydda människan och miljön.
Informationen kan lämnas på papper eller elektroniskt. Därefter skall tillverkaren, importören eller distributören till mottagaren av säkerhetsdatabladet sända sådan ny relevant information om ämnet som kommer till hans kännedom.
2. Allmänna regler för säkerhetsdatabladens utarbetande, distribution, innehåll och utformning skall fastställas i enlighet med förfarandet i artikel 29.4 a.
Artikel 28
Anpassning till den tekniska utvecklingen
Nödvändiga ändringar för att anpassa bilagorna till den tekniska utvecklingen skall beslutas i enlighet med förfarandet i artikel 29.
Artikel 29
Förfarandet vid anpassning till den tekniska utvecklingen
1. Kommissionen skall biträdas av en kommitté bestående av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Yttrandet skall beslutas med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Rösterna från medlemsstaternas företrädare i kommittén skall vägas på det sätt som föreskrivs i artikeln. Ordföranden får inte rösta.
3. Kommissionen skall själv anta förslaget om det är förenligt med kommitténs yttrande.
Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
4. a) Utom i de fall som avses i b) skall kommissionen om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits själv besluta att de föreslagna åtgärderna skall vidtas. I det fall som avses i artikel 31.2 skall tidsfristen vara sex veckor.
b) I fråga om åtgärder för anpassning till den tekniska utvecklingen som avser bilaga 2, 6, 7 och 8 skall kommissionen om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits själv besluta att de föreslagna åtgärderna skall vidtas, såvida inte rådet med enkel majoritet har avvisat förslaget.
Artikel 30
Klausul om fri rörelse
Medlemsstaterna får inte på grunder som rör anmälan, klassificering, förpackning eller märkning i detta direktivs mening förbjuda, begränsa eller hindra att ämnen som uppfyller kraven i detta direktiv släpps ut på marknaden.
Artikel 31
Skyddsklausul
1. Om en medlemsstat i ljuset av ny information på goda grunder anser att ett ämne som har bedömts uppfylla kraven i detta direktiv ändå utgör en fara för människan eller miljön på grund av att klassificeringen, förpackningen eller märkningen inte längre är riktig, kan den tillfälligt omklassificera ämnet eller, om så är nödvändigt, förbjuda att ämnet släpps ut på marknaden eller föreskriva att särskilda villkor skall gälla inom det egna territoriet. Den skall omedelbart meddela kommissionen och de andra medlemsstaterna om varje sådan åtgärd och motivera sitt beslut.
2. Kommissionen skall fatta ett beslut i enlighet med förfarandet i artikel 29.4 a.
3. Om kommissionen sedan beslut fattats i enlighet med punkt 2 anser att tekniska anpassningar av bilagorna till detta direktiv krävs för fall som avses i punkt 1 ovan, skall den fatta ett beslut i frågan i enlighet med förfarandet i artikel 29.
Artikel 32
Rapporter
1. Vart tredje år skall medlemsstaterna till kommissionen lämna en rapport om genomförandet av detta direktiv inom sina respektive territorier. Den första rapporten skall lämnas tre år efter genomförandet av detta direktiv.
2. Vart tredje år skall kommissionen på grundval av de uppgifter som avses i punkt 1 upprätta en samlad rapport som skall överlämnas till medlemsstaterna."
2. Artikel 24, 25 och 27 skall betecknas artikel 33, 34 och 35.
3. Bilaga 2, 6, 7 och 8 ändras härmed enligt följande:
- Bilaga 2 ändras genom tillägget av en symbol som betecknar miljöfara enligt bilaga 1 i detta direktiv.
- Bilaga 6 del 1 A ersätts av bilaga 2 till detta direktiv.
- Bilaga 7 ersätts av bilaga 3 till detta direktiv.
- Bilaga 8 ersätts av bilaga 4 till detta direktiv.
- I artikel 10.3 och 11 ersätts "artikel 8c" med "artikel 28".
3. Direktiv 78/631/EEG:
- I artikel 6.2 g ersätts "artikel 6" med "artikel 23".
- I artikel 10.3 och 11 ersätts "artikel 8 c" av "artikel 28".
4. Direktiv 88/379/EEG:
- I det andra och det åttonde stycket i ingressen ersätts hänvisningen till direktiv 79/831/EEG med en hänvisning till föreliggande direktiv.
- I artikel 3.3 ersätts "cancerogena, mutagena och teratogena verkningar" med "cancerogena och mutagena egenskaper samt verkningar på fortplantningen".
- I artikel 3.5 ersätts "artikel 8.2 i direktiv 67/548/EEG" med "artikel 13.3 i direktiv 67/548/EEG".
- Artikel 3.5 o skall ha följande lydelse:
"o) Preparat skall anses som skadliga för fortplantningen och tilldelas åtminstone farosymbolen och faroangivelsen "giftigt" om de innehåller ett ämne som har sådana verkningar och som tilldelas minst en av de R-fraser enligt bilaga 6 till direktiv 67/548/EEG som betecknar ämnen som skadliga för fortplantningen i kategori 1, i koncentrationer som motsvarar eller överstiger
- antingen de koncentrationer som anges i bilaga 1 till direktiv 67/548/EEG för ämnet i fråga, eller
- den koncentration som anges i punkt 6 i bilaga 1 (tabell VI) till detta direktiv, om ämnet inte är upptaget i bilaga 1 till direktiv 67/548/EEG eller förekommer där, men utan angivande av koncentrationsgränser."
- Artikel 3.5 p skall ha följande lydelse:
"p) Preparat skall anses behöva behandlas som skadliga för fortplantningen och tilldelas minst farosymbolen och faroangivelsen "giftigt" om de innehåller ett ämne som har sådana verkningar och som tilldelas minst en av de R-fraser enligt bilaga 6 till direktiv 67/548/EEG som betecknar ämnen som är skadliga för fortplantningen enligt kategori 2, i koncentrationer som motsvarar eller överstiger
- antingen de koncentrationer som anges i bilaga 1 till direktiv 67/548/EEG för ämnet i fråga, eller
- den koncentration som anges i punkt 6 i bilaga 1 (tabell VI) till detta direktiv, om ämnet inte är upptaget i bilaga 1 till direktiv 67/548/EEG eller förekommer där, men utan angivande av koncentrationsgränser."
- Artikel 3.5 q skall ha följande lydelse:
"q) Preparat skall anses behöva behandlas som skadliga för fortplantningen och tilldelas minst farosymbolen och faroangivelsen "giftigt" om de innehåller ett ämne som har sådana verkningar och som tilldelas minst en av de R-fraser enligt bilaga 6 till direktiv 67/548/EEG som betecknar ämnen som är skadliga för fortplantningen i kategori 3, i koncentrationer som motsvarar eller överstiger
- antingen de koncentrationer som anges i bilaga 1 till direktiv 67/548/EEG för ämnet i fråga, eller
- den koncentration som anges i punkt 6 i bilaga 1 (tabell VI) till detta direktiv, om ämnet inte är upptaget i bilaga 1 till direktiv 67/548/EEG eller förekommer där, men utan angivelse av koncentrationsgränser."
- I artikel 6.1 a ersätts "artikel 15.1" med "artikel 22.1".
- I artikel 6.3 ersätts "artikel 21" av "artikel 28".
- I artikel 7.1 c ii ersätts "artikel 11.4" av "artikel 19.4".
- I artikel 7.1 ersätts "artikel 16.2 c" av "artikel 23.2 c".
- Följande punkt infogas i artikel 8:
"3a De i artikel 7 föreskrivna uppgifterna på etiketten skall framträda tydligt mot bakgrunden och skall vara tryckta i så stor stil och med så stora mellanrum att de är lätta att läsa.
Särskilda bestämmelser om upplysningarnas uppställning och format förs in i bilaga 6 till direktiv 67/548/EEG i enlighet med förfarandet i artikel 28.4 b i nämnda direktiv".
- I artikel 10, 14.2 och 15 ersätts "artikel 21" med "artikel 28".
- I rubriken till bilaga 1, del 6 ersätts "teratogena verkningar" med "verkningar på fortplantningen".
- I bilaga 1 tabell 6 ersätts "teratogena ämnen" med "ämnen som är skadliga för fortplantningen".
Artikel 3
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 oktober 1993. De skall genast underrätta kommissionen om detta.
2. När dessa åtgärder beslutas av medlemsstaterna skall författningarna innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
3. Medlemsstaterna skall till kommissionen överlämna texterna till nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV 92/77/EEG av den 19 oktober 1992 med tillägg till det gemensamma systemet för mervärdesskatt och med ändring av direktiv 77/388/EEG (harmonisering av mervärdesskattesatser)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av kommissionens förslag(),
med beaktande av Europaparlamentets yttrande(),
med beaktande av ekonomiska och sociala kommitténs yttrande(), och
med beaktande av följande: Fullbordandet av den inre marknaden, vilket är ett av de grundläggande målen för gemenskapen, kräver som ett första steg att tull- och skattekontrollerna vid gränserna avskaffas.
För att snedvridningar skall undvikas förutsätter avskaffandet av dessa kontroller vad gäller mervärdesskatt inte endast en enhetlig skattebas utan även att ett flertal skattesatser och skattenivåer ligger tillräckligt nära varandra mellan medlemsstaterna. Det är därför nödvändigt att ändra direktiv 77/388/EEG().
Under övergångstiden bör vissa undantag från reglerna beträffande skatternas antal och nivå vara möjliga.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 77/388/EEG ändras på följande sätt:
1. Artikel 12.3 skall ersättas med följande:
"3. a) Från och med den 1 januari 1993 skall medlemsstaterna tillämpa en normalskattesats, vilken till och med den 31 december 1996 inte får vara lägre än 15%.
På grundval av den rapport om hur övergångsbestämmelserna har fungerat och de förslag till slutgiltiga bestämmelser som kommissionen skall lägga fram i överensstämmelse med artikel 281, skall rådet före den 31 december 1995 enhälligt besluta om den lägsta skattesatsnivå som efter den 31 december 1996 skall tillämpas såsom normalskattesats.
Medlemsstaterna får även tillämpa en eller två reducerade skattesatser. Dessa får inte vara lägre än 5 % och får endast avse tillhandahållande av sådana varor och tjänster som anges i bilaga H.
b) Medlemsstaterna får tillämpa en reducerad skattesats på tillhandahållande av naturgas och elektricitet, under förutsättning att ingen risk för snedvridande verkningar på konkurrensen föreligger. En medlemsstat som avser att tillämpa en sådan skattesats skall underrätta kommissionen innan så sker. Kommissionen skall fatta beslut beträffande förekomsten av risk för snedvridning av konkurrensen. Om kommissionen inte har gjort detta inom tre månader efter mottagandet av sådan underrättelse, anses någon risk för snedvridning av konkurrensen inte föreligga.
c) Regler om vilka skattesatser som skall tillämpas på konstverk, antikviteter och samlarföremål fastställs genom direktivet med specialbestämmelser för begagnade varor, konstverk, antikviteter och samlarföremål. Rådet skall anta detta direktiv före den 31 december 1992.
d) Regler om beskattningen av andra jordbruksprodukter än sådana som tillhör kategori 1 i bilaga H skall enhälligt antas av rådet före den 31 december 1994 på grundval av kommissionens förslag.
Intill dess kan de medlemsstater som för närvarande tillämpar reducerad skattesats fortsätta att göra det; de som för närvarande tillämpar normalskattesats kan däremot inte tillämpa reducerad skattesats. Detta medger ett tvåårigt uppskov med införandet av normalskattesatsen.
e) De regler och skattesatser som skall tillämpas på guld skall fastställas genom ett direktiv med specialbestämmelser om guld. Kommissionen skall lägga fram ett förslag härom i sådan tid att det kan enhälligt antagas av rådet före den 31 december 1992.
Medlemsstaterna kommer från och med den 1 januari 1993 att vidta alla nödvändiga åtgärder för att bekämpa bedrägeri och annan oredlighet på detta område. Dessa åtgärder får inbegripa införandet av ett system för redovisning av mervärdesskatt på tillhandahållande av guld mellan skattskyldiga personer inom samma medlemsstat, vilket låter köparen betala skatt för säljarens räkning och samtidigt ger köparen rätt till avdrag med samma belopp som ingående skatt."
2. Första meningen i artikel 12.4 skall utgå.
3. Följande stycke läggs till i artikel 12.4:
"På grundval av kommissionens rapport skall rådet vartannat år, med början 1994, granska omfattningen av de reducerade skattesatserna. Rådet kan på kommissionens förslag enhälligt besluta att ändra i förteckningen över varor och tjänster i bilaga H."
4. Artikel 28.2 ersätts med följande:
"2. Utan hinder av artikel 12.3 skall följande bestämmelser gälla under den övergångsperiod som nämns i artikel 28l:
a) Undantag med återbetalning av skatt som erlagts i föregående led, och reducerade skattesatser som är lägre än den minimiskattesats som lagts fast i artikel 12.3 vad gäller de reducerade skattesatser som var i kraft den 1 januari 1991 och som står i överensstämmelse med gemenskapslagstiftningen och uppfyller de villkor som stadgas i artikel 17 sista strecksatsen i rådets andra direktiv av den 11 april 1967, får bibehållas.
Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa bestämningen av egna resurser i samband med dessa operationer.
I händelse av att bestämmelserna i denna punkt för Irlands del skulle skapa snedvridning av konkurrensen när det gäller tillhandahållande av energiprodukter för uppvärmning och belysning, kan kommissionen på särskild begäran ge Irland rätt att tillämpa en reducerade skattesats på sådant tillhandahållande, i enlighet med artikel 12.3. I sådant fall skall Irland inlämna sin begäran till kommissionen tillsammans med alla nödvändiga upplysningar. Om kommissionen inte har fattat något beslut inom tre månader efter mottagandet av denna begäran, skall Irland anses ha fått rätt att tillämpa den föreslagna reducerade skattesatsen.
b) Medlemsstater som den 1 januari 1991 på andra varor och tjänster än sådana som anges i bilaga H i överensstämmelse med gemenskapslagstiftningen tillämpade regler om undantag med återbetalning av skatt som erlagts i föregående led eller reducerade skattesatser som var lägre än det minimum som lagts fast i artikel 12.3 vad gäller reducerade skattesatser får tillämpa den reducerade skattesatsen eller den ena av de två reducerade skattesatser som nämns i artikel 12.3 på sådana varor eller tjänster.
c) Medlemsstater som enligt villkoren i artikel 12.3 måste höja den normalskattesats som gällde den 1 januari 1991 med mer än 2 %, får tillämpa en reducerad skattesats som är lägre än det minimum som fastlagts i artikel 12.3 vad gäller den reducerade skattesatsen på sådana kategorier av varor och tjänster som specificeras i bilaga H. Vidare får dessa medlemsstater tillämpa en sådan skattesats på restaurangtjänster, barnkläder, barnskor och bostäder. Medlemsstaterna får inte med stöd av detta stycke införa regler om undantag med återbetalning av skatten i föregående led.
d) Medlemsstater som den 1 januari 1991 tillämpade en reducerad skattesats på restaurangtjänster, barnkläder, barnskor och bostäder får fortsätta att tillämpa denna på dessa områden.
e) Medlemsstater som den 1 januari 1991 tillämpade en reducerad skattesats på andra varor och tjänster än sådana som specificeras i bilaga H får tillämpa denna reducerade skattesats eller en av de två reducerade skattesatser som nämns i artikel 12.3 på dessa områden, förutsatt att skattesatsen inte understiger 12 %.
f) Grekland får tillämpa mervärdesskattesatser som är intill 30 % lägre än motsvarande skattesatser på det grekiska fastlandet i departementen Lesbos, Chios, Samos, Dodekaneserna och Cykladerna, liksom på följande öar i Egeiska havet: Thasos, Norra Sporaderna, Samothrake och Skiros.
g) Rådet skall på grundval av en rapport från kommissionen före den 31 december 1994 på nytt granska bestämmelserna i a-f ovan med särskild hänsyn till den inre marknadens riktiga funktion. I den händelse betydande snedvridning av konkurrensen uppstår, skall rådet på kommissionens förslag enhälligt besluta om lämpliga åtgärder."
5. Bilaga H i bilagan till detta direktiv skall bifogas.
Artikel 2
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 december 1992. De skall genast underrätta kommissionen härom.
När medlemsstaterna antar dessa åtgärder, skall besluten innehålla en hänvisning till detta direktiv eller åtföljas av sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EEG) nr 305/92 av den 7 februari 1992 om ändring av förordning (EEG) nr 410/90 om fastställande av kvalitetsnormer för kiwifrukt
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1035/72 av den 18 maj 1972 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom förordning (EEG) nr 1623/91(2), särskilt artikel 2.2 andra stycket i denna, och med beaktande av följande:
I kommissionens förordning (EEG) nr 410/90(3) fastställs kvalitetsnormer för kiwifrukt.
Vissa av bestämmelserna skiljer sig mellan de olika språkversionerna. Dessa bestämmelser bör därför ändras.
För att anpassa kvalitetsnormerna för kiwifrukt till de övriga EEG-normerna för frukt och grönsaker bör det göras ändringar vad avser "hållbarhet", "storlek" och "storlekssortering".
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för frukt och grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
b) Det tredje stycket under "ii) Klass I" skall i alla språkversioner ha följande lydelse:
"Den skall ha sorttypiska egenskaper. Följande smärre fel är dock tillåtna om de inte påverkar produktens allmänna utseende, kvaliteten, hållbarheten och förpackningens presentation:
- Ett mindre fel i formen (dock inte svullnader eller missbildningar).
- Ett mindre färgfel.
- Ytliga skador på skalet som täcker en yta av högst 1 cm².
- Ett mindre "Haywardmärke" i form av längsgående linjer men utan förhöjning."
c) Under "iii) Klass II" skall tredje stycket fjärde strecksatsen angående "Haywardmärken ha följande lydelse:
" - Flera mer uttalade "Hayward-märken" med mindre förhöjning."
2. Under "III. Bestämmelser angående storlekssortering" skall första stycket ha följande lydelse:
"Storleken bestäms av fruktens vikt."
3. Följande ändringar skall göras i del V. "Bestämmelser angående presentation":
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EEG) nr 762/92 av den 27 mars 1992 om ändring av bilaga V i rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), ändrad genom kommissionens förordning (EEG) nr 675/92(2), särskilt artikel 11, och med beaktande av följande:
För att uppnå en effektiv administration är det önskvärt att de upplysningar som skall ingå i en anhållan om fastställande av gränsvärde för farmakologiskt verksamma ämnen i veterinärmedicinska produkter i enlighet med förordning (EEG) nr 2377/90 så mycket som möjligt motsvarar de uppgifter som skall lämnas till medlemsstaterna i en ansökan om tillstånd att släppa ut en veterinärmedicinsk produkt på marknaden, vilken inges i enlighet med artikel 5 i rådets direktiv 81/851/EEG av den 28 september 1981 om tillnärmning av medlemsstaternas lagstiftning om veterinärmedicinska läkemedel(3), ändrat genom direktiv 90/676/EEG(4).
Det är nödvändigt att ändra bilaga V i förordning (EEG) nr 2377/90 för att beakta de ändringar som gjorts ifråga om kraven vid prövning av veterinärmedicinska produkter vilka infördes genom kommissionens direktiv 92/18/EEG av den 20 mars 1992 om ändring av bilaga till rådets direktiv 81/852/EEG om tillnärmning av medlemsstaternas lagstiftning om analytiska, farmakologiska, toxikologiska och kliniska normer och prövningsplaner för veterinärmedicinska läkemedel.
Bestämmelserna i denna förordning är förenliga med yttrandet från Kommittén för anpassning till den tekniska utvecklingen av direktiven om avlägsnande av tekniska handelshinder inom den veterinärmedicinska sektorn, inrättad genom artikel 2b i rådets direktiv 81/852/EEG(5), ändrat genom direktiv 87/20/EEG(6).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
RÅDETS FÖRORDNING (EEG) nr 1764/92 av den 29 juni 1992 om ändring av ordningen för import till gemenskapen av vissa jordbruksprodukter som har sitt ursprung i Algeriet, Cypern, Egypten, Israel, Jordanien, Libanon, Malta, Marocko, Syrien och Tunisien
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 113 i detta,
med beaktande av kommissionens förslag, och
med beaktande av följande: Inom den allmänna ramen för den förnyade medelhavspolitiken antog rådet och kommissionen en resolution om handel med icke-medlemsstater i medelhavsområdet på rådets möte den 18 och 19 december 1990, i syfte att stärka banden och öka samarbetet med länderna i regionen.
I denna resolution fastställs särskilt genomförandet av åtgärder för att främja jordbruksexport från dessa länder till gemenskapen, och närmare bestämmelser för tillämpningen av åtgärderna måste därför definieras.
För att kunna göra detta är det nödvändigt att ändra ordningen för import till gemenskapen, som omfattas av bestämmelserna i protokollen till associerings- eller samarbetsavtal med Algeriet, Cypern, Egypten, Israel, Jordanien, Libanon, Malta, Marocko, Syrien och Tunisien.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. De tullar som gäller den 31 december i gemenskapen i dess sammansättning den 31 december 1985 för de produkter som förtecknas i bilaga II till fördraget och som har sitt ursprung i de berörda icke-medlemsländerna i medelhavsområdet och för vilka tullavveckling utsträcks till tiden efter den 1 januari 1993 enligt de protokoll till associerings- eller samarbetsavtal som finns i bilaga 1 till denna förordning skall upphävas i två lika steg från och med den 1 januari 1992 och från och med den 1 januari 1993.
2. Punkt 1 tillämpas inom ramarna, om sådana finns, för tullkvoter och tidsscheman som fastställts i de protokoll som avses i den punkten och skall beakta de särskilda bestämmelser som där fastställs.
3. Som ett resultat av tillämpningen av punkt 1 skall tullarna upphävas helt när de når en nivå på 2 % eller mindre.
RÅDETS FÖRORDNING (EEG) nr 2077/92 av den 30 juni 1992 om branschorganisationer och branschavtal inom tobakssektorn
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 42 och 43 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Utvecklingen på medellång och lång sikt av gemenskapens och världens jordbruksmarknader gör det nödvändigt att ompröva vissa instrument inom den gemensamma jordbrukspolitiken för att återskapa balans på marknaden. Dessa justeringar, som principiellt syftar till att skapa mera flexibla former för marknadsstödet, förutsätter att aktörerna på marknaden ändrar sitt ekonomiska beteende och tar större hänsyn till den faktiska situationen på marknaden.
Branschorganisationer som bildats av enskilda eller grupper och som representerar en betydande del av de olika kategorier som är sysselsatta med produktion, beredning och avsättning inom tobakssektorn skulle sannolikt komma att bidra till att större hänsyn tas till situationen på marknaden liksom till att uppmuntra förändringar i det ekonomiska beteendet i syfte att förbättra kunskapen om och organisationen av produktionen, beredningen och avsättningen. Deras verksamhet skulle i vissa fall kunna bidra till att förbättra balansen på marknaden och därigenom medverka till att målen enligt artikel 39 i fördraget uppfylls. Det bör därför fastställas vilka åtgärder som skulle kunna utgöra ett sådant bidrag från branschorganisationernas sida.
Det förefaller därför lämpligt att särskilt erkänna de organisationer som kan påvisa att de är representativa på regional eller interregional nivå eller på gemenskapsnivå och som aktivt strävar efter att förverkliga de ovan nämnda målen. Ett sådant erkännande bör kunna beviljas av medlemsstaten eller av kommissionen, beroende på hur omfattande branschorganisationens verksamhet är.
För att stödja den del av branschorganisationernas verksamhet som är av särskilt intresse med tanke på de nuvarande reglerna om den gemensamma organisationen av marknaden inom tobakssektorn bör bestämmelser införas som gör det möjligt att på vissa villkor utvidga de regler som en branschorganisation antagit för sina medlemmar till att även omfatta alla producenter eller producentgrupper, även de som inte är medlemmar, i en eller flera regioner. Icke medlemmar bör också kunna vara skyldiga att betala hela eller del av den medlemsavgift som är avsedd att täcka de kostnader för nämnda verksamhet som inte avser administration. Denna ordning bör genomföras på ett sådant sätt att berörda socioekonomiska gruppers rättigheter garanteras, särskilt konsumentens rättigheter.
Andra verksamheter som de erkända branschorganisationerna bedriver kan vara av allmänt ekonomiskt eller tekniskt intresse för tobakssektorn och därmed vara värdefulla för alla som är sysselsatta inom branscherna i fråga, vare sig de är medlemmar i organisationen eller inte. I dessa fall förefaller det rimligt att icke medlemmar betalar den medlemsavgift som är avsedd att täcka andra kostnader än de rent administrativa som uppkommer som en direkt följd av verksamheten i fråga.
För att säkerställa att programmet fungerar på ett riktigt sätt bör det etableras ett nära samarbete mellan medlemsstaterna och kommissionen, varvid kommissionen bör ha en stående kontrollbefogenhet, särskilt vad gäller erkännandet av de branschorganisationer som arbetar på regional eller interregional nivå och vad gäller de avtal och de samordnade förfaranden som dessa organisationer tillämpar.
För att informera medlemsstaterna och andra intressenter bör det i början av varje år offentliggöras en lista över de organisationer som erkänts under det föregående året och en lista över de organisationer som fått sitt erkännande återkallat under samma period samt de bestämmelser som fått ett utvidgat tillämpningsområde med angivande av deras omfattning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
3. bedriver några av följande verksamheter på regional nivå i en eller flera regioner inom gemenskapen eller inom hela gemenskapen, och därvid beaktar konsumentintressena:
a) Medverkan till ökad samordning av avsättningen av tobak i blad och tobak i balar.
b) Utarbetande av standardavtal som är i överensstämmelse med gemenskapens bestämmelser.
c) Förbättrande av kunskapen om och insynen i marknaden.
d) Ökning av produkternas förädlingsvärde, särskilt genom marknadsföringsåtgärder och forskning om nya användningsområden som inte utgör ett hot mot folkhälsan.
e) Omorientering av branschen mot produkter som bättre tillgodoser marknadens behov och hänsynen till folkhälsan.
f) Forskning om metoder som gör det möjligt att begränsa användningen av växtskyddsmedel samtidigt som produktens kvalitet säkerställs och jorden skyddas.
g) Utveckling av metoder och medel för förbättring av produktkvaliteten i produktions- och beredningsledet.
2. Före erkännandet skall medlemsstaterna anmäla till kommissionen vilka branschorganisationer som ansökt om erkännande och lämna all nödvändig information om vilka näringsgrenar de omfattar, hur representativa de är, vilka verksamheter de bedriver samt den övriga information som behövs för att ta ställning till ansökan.
Kommissionen kan inom 60 dagar efter medlemsstatens anmälan motsätta sig ett erkännande.
3. Medlemsstaten skall återkalla erkännandet om
a) de krav som anges i denna förordning inte längre uppfylls,
b) branschorganisationen överträder ett eller flera av de förbud som anges i artikel 7.3, utan att det påverkar tillämpningen av rättsliga förfaranden enligt nationell lagstiftning,
c) branschorganisationen underlåter att uppfylla anmälningsplikten enligt artikel 7.2.
Medlemsstaterna skall omedelbart underrätta kommissionen om beslut om återkallande av erkännandet.
Artikel 4
1. Kommissionen skall efter ansökan erkänna branschorganisationer som
a) helt eller delvis bedriver sin verksamhet inom flera medlemsstaters territorier eller inom hela gemenskapen,
b) har bildats i överensstämmelse med en medlemsstats lagstiftning eller gemenskapsrätten
c) uppfyller föreskrifterna i artikel 3.1 b d.
2. Kommissionen skall underrätta de medlemsstater inom vilkas territorier branschorganisationen bildats och dess verksamhet bedrivs om inkomna ansökningar om erkännande. De berörda medlemsstaterna skall därefter ha två månader på sig att inkomma med synpunkter.
Kommissionen skall fatta beslut om erkännande inom tre månader efter det att den har mottagit ansökan och all information.
3. Kommissionen skall återkalla erkännandet av de organisationer som anges i punkt 1 i de fall som anges i artikel 3.3.
Artikel 5
Kommissionen skall offentliggöra namnen på de branschorganisationer som erkänts i C-serien av Europeiska gemenskapernas officiella tidning och samtidigt ange inom vilken ekonomisk sektor eller geografiskt område de är verksamma och vilka av de i artikel 2 angivna verksamheterna som de bedriver. Återkallanden av erkännanden skall också offentliggöras.
Artikel 6
Erkännandet av branschorganisationer innebär att de tillåts bedriva de verksamheter som anges i artikel 2.3 på de villkor som föreskrivs i denna förordning.
Artikel 7
1. Utan hinder av artikel 1 i förordning nr 26(4) skall artikel 85.1 i fördraget inte tillämpas på de avtal och samordnade förfaranden som de erkända branschorganisationerna ingått för genomförande av de åtgärder som anges i artikel 2.3.
2. Punkt 1 skall tillämpas endast om
- avtalen och de samordnade förfarandena anmälts till kommissionen, och
- kommissionen inom tre månader efter det att den har erhållit alla de upplysningar som behövs inte har funnit att avtalen eller de samordnade förfarandena är oförenliga med gemenskapens bestämmelser.
Avtalen och de samordnade förfarandena får inte träda i kraft förrän denna period löpt ut.
3. Avtal och samordnade förfaranden skall under alla omständigheter förklaras vara oförenliga med gemenskapens bestämmelser om de
- kan leda till någon form av uppdelning av marknaderna inom gemenskapen,
- kan medföra att den gemensamma organisationen av marknaden störs,
- kan medföra en snedvridning av konkurrensen som inte är nödvändig för att uppnå målen för den gemensamma jordbrukspolitik som branschåtgärderna syftar till.
- innebär ett fastställande av priser eller kvoter, utan att det påverkar tillämpningen av åtgärder som branschorganisationerna vidtar till följd av särskilda bestämmelser som fastställts av gemenskapen,
- kan innebära särbehandling eller sätta konkurrensen ur spel för en betydande del av produkterna i fråga.
Detta beslut får inte träda i kraft tidigare än det datum då den berörda branschorganisationen underrättats om beslutet, såvida inte branschorganisationen har lämnat felaktiga uppgifter eller missbrukat det undantag som anges i punkt 1.
Artikel 8
1. Branschorganisationerna kan begära att vissa av deras avtal eller samordnade förfaranden inom det område där de är verksamma för en begränsad tid görs bindande för enskilda och grupper inom den berörda ekonomiska sektorn som inte är medlemmar i någon organisation som ingår i branschorganisationen.
Branschorganisationerna måste för att få utvidga tillämpningsområdet för sina bestämmelser företräda minst två tredjedelar av den berörda produktionen eller handeln. Om den föreslagna utvidgningen berör flera regioner, måste branschorganisationerna påvisa att de uppnår en viss minsta nivå i fråga om representativitet inom varje näringsgren och varje region.
2. De bestämmelser, för vilka ett utvidgat tillämpningsområde begärs, skall ha tillämpats i minst ett år och avse ett av följande områden:
a) Kunskap om produktionen och marknaden.
b) Fastställande av minimikvantiteter.
c) Användande av miljövänliga odlingsmetoder.
d) Fastställande av minimistandarder för förpackning och presentation.
e) Användande av certifierat utsäde och kontroll av produktkvaliteten.
3. En utvidgad tillämpning av bestämmelserna skall godkännas av kommissionen i enlighet med det förfarande som anges i artikel 9.
Artikel 9
1. Då det gäller bestämmelser antagna av branschorganisationer som erkänts av medlemsstaterna, svarar medlemsstaterna för att berörda intressenter informeras genom offentliggörande av de avtal och samordnade förfaranden vars tillämpning avses utvidgas till att omfatta enskilda eller grupper som inte tillhör någon branschorganisation i en viss region eller grupp av regioner.
De berörda intressenterna skall ha två månader på sig att lämna sina synpunkter.
2. Vid slutet av denna period och innan beslut fattas, skall medlemsstaterna anmäla till kommissionen vilka bestämmelser de avser att göra bindande och samtidigt lämna all relevant information. I anmälan skall ingå alla de synpunkter som erhållits efter offentliggörandet enligt punkt 1 och en bedömning av ansökan om utvidgad tillämpning.
3. Kommissionen skall i C-serien av Europeiska gemenskapernas officiella tidning offentliggöra de bestämmelser för vilka utvidgad tillämpning som begärts av de branschorganisationer som den erkänt enligt artikel 4. Efter offentliggörandet skall medlemsstaterna och de berörda intressenterna ha två månader på sig att lämna sina synpunkter.
4. Om de bestämmelser för vilka utvidgad tillämpning begärs är "tekniska föreskrifter" i den betydelse som anges i direktiv 83/189/EEG(5), skall de anmälas till kommissionen i enlighet med artikel 8 i det direktivet samtidigt med den i punkt 2 angivna anmälan.
Om förutsättningarna för att avge ett detaljerat utlåtande enligt artikel 9 i det direktivet är uppfyllda, skall kommissionen, vägra godkänna de bestämmelser för vilka utvidgad tillämpning begärs, utan att detta påverkar tillämpningen av punkt 5.
5. Kommissionen skall senast tre månader efter medlemsstatens anmälan fatta beslut i enlighet med punkt 2 och, i det fall punkt 3 är tillämplig, senast fem månader efter offentliggörandet av ansökan om utvidgad tillämpning av bestämmelserna i Europeiska gemenskapernas officiella tidning.
Kommissionen skall under alla omständigheter avslå ansökan om den finner att den utvidgade tillämpningen
- förhindrar konkurrensen på en betydande del av den gemensamma marknaden,
- begränsar frihandeln, eller
- äventyrar målen för den gemensamma jordbrukspolitiken eller andra delar av gemenskapslagstiftningen.
6. De bestämmelser för vilka man ansökt om utvidgad tillämpning skall offentliggöras i Europeiska gemenskapernas officiella tidning.
7. Om bestämmelser i enlighet med denna artikel gjorts bindande för näringsidkare som inte är medlemmar i en branschorganisation, får medlemsstaten eller kommissionen, det som är lämpligast från fall till fall, besluta att enskilda eller grupper som inte är medlemmar skall betala till organisationen hela eller del av medlemsavgiften, utom för den del av avgiften som används för att täcka administrativa kostnader i samband med tillämpningen av bestämmelserna eller de samordnade förfarandena.
Artikel 10
1. När en eller flera av de i punkt 2 angivna verksamheterna bedrivs av en erkänd branschorganisation och är av allmänt ekonomiskt intresse för de personer vilkas verksamhet är knuten till en eller flera av produkterna, får medlemsstaten som beviljat erkännandet eller kommissionen, om erkännandet beviljats i enlighet med artikel 4, besluta att enskilda eller grupper som inte är medlemmar i sammanslutningen men som drar nytta av dess verksamhet skall betala till organisationen hela eller del av medlemsavgiften, i den mån medlemsavgiften är avsedd att täcka kostnader som är en direkt följd av verksamheten med undantag av varje form av administrationskostnad.
2. De verksamheter som avses i denna artikel skall anknyta till något eller några av följande områden:
- Forskning för att öka förädlingsvärdet på produkterna, särskilt genom nya användningsområden som inte utgör ett hot mot folkhälsan.
- Undersökningar om hur kvaliteten på bladtobak och tobak i balar kan förbättras.
- Forskning om odlingsmetoder som medger en minskad användning av växtskyddsmedel och garanterar att jorden och miljön skyddas.
3. De berörda medlemsstaterna skall anmäla till kommissionen vilka beslut som de avser att fatta enligt punkt 1. Dessa beslut får träda i kraft tidigast tre månader efter tidpunkten för anmälan till kommissionen. Kommissionen får inom denna tid kräva att hela eller delar av förslaget till beslut förkastas, om det allmänna ekonomiska intresse som hävdas inte förefaller välgrundat.
4. Om de verksamheter som en av kommissionen enligt artikel 4 erkänd branschorganisation bedriver är av allmänt ekonomiskt intresse, skall kommissionen anmäla sitt förslag till beslut till de berörda medlemsstaterna, som sedan har två månader på sig att lämna sina synpunkter.
Artikel 11
Varje beslut som medlemsstaterna eller kommissionen fattar om åtgärder som innebär att enskilda eller grupper som inte är medlemmar i en branschorganisation skall betala avgift skall offentliggöras i Europeiska gemenskapernas officiella tidning. Beslutet får träda i kraft tidigast två månader efter tidpunkten för offentliggörandet.
Artikel 12
Tillämpningsföreskrifter till denna förordning skall fastställas i enlighet med det förfarande som anges i artikel 23 i förordning (EEG) nr 2075/92(6).
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel
Som ett led i anpassningen av den gemensamma jordbrukspolitiken bör diversifiering av jordbruksproduktionen uppmuntras så att det blir bättre balans mellan tillgång och efterfrågan. Stimulerad efterfrågan på produkter med särskilda egenskaper skulle kunna vara till stort gagn för landsbygdens ekonomi, särskilt i mindre gynnade eller avlägset belägna trakter, genom att denna förbättras och odlarnas inkomster och avfolkning förebyggs i dessa trakter.
Det har också på senare år iakttagits att konsumenterna tenderar att fästa större vikt vid livsmedlens kvalitet än kvantitet. Intresset för speciella produkter skapar en allt större efterfrågan på jordbruksprodukter och livsmedel med känt geografiskt ursprung.
Med tanke på mångfalden av marknadsförda produkter och överflödet av information om dem måste konsumenterna för att kunna göra ett bra val få klar och koncis information om produkternas ursprung.
Märkningen av jordbruksprodukter och livsmedel är underkastad de allmänna regler som anges i rådets direktiv 79/112/EEG av den 18 december 1978 om tillnärmning av medlemsstaternas lagstiftning om märkning, presentation och reklam i fråga om livsmedel(4). Med hänsyn till den särskilda beskaffenheten hos jordbruksprodukter och livsmedel bör speciella regler införas om jordbruksprodukter och livsmedel från ett särskilt geografiskt område.
Strävan att skydda jordbruksprodukter eller livsmedel som har ett känt geografiskt ursprung har gjort att vissa medlemsstater har infört registrerade ursprungsbeteckningar. Dessa har visat sig vara till gagn för producenterna som kunnat tillförsäkra sig större inkomster genom verkliga insatser för att förbättra kvaliteten, och för konsumenterna som får möjlighet att köpa högkvalitetsprodukter med garanti beträffande produktionsmetod och ursprung.
Det finns emellertid nationella olikheter i sättet att ordna registrering av ursprungsbeteckning och geografisk beteckning. En gemenskapsmetod bör planeras. Ett gemensamt regelverk för skydd av dessa beteckningar gör det möjligt att utveckla dessa, eftersom ett sådant skydd med enhetlig metod säkerställer konkurrens på lika villkor mellan produkter med sådana beteckningar och höjer produkternas trovärdighet i konsumenternas ögon.
De planerade reglerna bör ta hänsyn till redan befintlig gemenskapslagstiftning om vin och spritdrycker som ger högre skyddsnivå.
Denna förordnings räckvidd begränsas till vissa jordbruksprodukter och livsmedel där det finns ett samband mellan egenskaperna hos produkten eller livsmedlet och det geografiska ursprunget. Räckvidden kan sedermera ökas så att också andra produkter eller livsmedel omfattas.
Nuvarande bruk gör det lämpligt att definiera två slags geografiska beskrivningar, nämligen skyddade geografiska beteckningar och skyddade ursprungsbeteckningar.
En jordbruksprodukt eller ett livsmedel som bär en sådan beteckning måste uppfylla vissa villkor som anges i en specifikation.
För att en geografisk beteckning eller en ursprungsbeteckning skall åtnjuta skydd i varje medlemsstat måste den registreras på gemenskapsnivå. Registreringen skall också ge information om produkten eller livsmedlet till dem som sysslar med handel samt till konsumenterna.
Registreringsförfarandet bör ge var och en som personligen och direkt berörs i en medlemsstat möjlighet att tillvarata sina rättigheter genom att till kommissionen framställa invändningar.
Med hänsyn till den tekniska utvecklingen bör det finnas förfaranden som gör det möjligt att ändra specifikationen efter det att registrering skett eller att ur registret avföra den geografiska beteckningen eller ursprungsbeteckningen för en jordbruksprodukt eller ett livsmedel om produkten eller livsmedlet inte längre överensstämmer med den specifikation som låg till grund när skyddet beviljades för beteckningen.
Föreskrifter bör införas för handeln med tredje land som erbjuder likvärda garantier för utfärdande och kontroll av geografiska beteckningar och ursprungsbeteckningar på deras territorium.
Föreskrifter bör införas för ett förfarande som innebär nära samverkan mellan medlemsstaterna och kommissionen genom en regleringskommitté som inrättas för ändamålet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Denna förordning fastställer regler för skydd av ursprungsbeteckningar och geografiska beteckningar för sådana jordbruksprodukter som är avsedda att förtäras av människor och som avses i bilaga 2 till fördraget och för sådana livsmedel som avses i bilaga 1 till denna förordning och de jordbruksprodukter som förtecknats i bilaga 2 till denna förordning.
Denna förordning skall dock inte tillämpas på vinprodukter och spritdrycker.
Bilaga 1 kan ändras enligt det förfarande som fastställs i artikel 15.
2. Denna förordning skall tillämpas utan att påverka andra särskilda gemenskapsregler.
3. Rådets direktiv 83/189/EEG av den 28 mars 1983 om ett informationsförfarande beträffande tekniska standarder och föreskrifter(5) skall inte tillämpas på ursprungsbeteckningar och geografiska beteckningar som omfattas av denna förordning.
- som härstammar från ifrågavarande region, ort eller land,
och - vars kvalitet eller egenskaper helt eller väsentligen beror på viss geografisk omgivning med de naturliga och mänskliga faktorer som därtill hör och vars framställning, bearbetning och beredning äger rum i det ifrågavarande geografiska området.
b) geografisk beteckning: Namn på en region, en ort eller i undantagsfall ett land, använt för att beskriva en jordbruksprodukt eller ett livsmedel
- som härstammar från ifrågavarande region, ort eller land,
och - som besitter viss kvalitet, har visst anseende eller äger viss annan egenskap som kan hänföras till detta geografiska ursprung och som framställs, bearbetas och bereds i det ifrågavarande geografiska området.
3. Vissa traditionella geografiska eller icke-geografiska namn på en jordbruksprodukt eller ett livsmedel som härstammar från en viss region eller viss ort och som uppfyller de villkor som avses i andra strecksatsen i punkt 2 a skall också betraktas som ursprungsbeteckningar.
4. Trots punkt 2 a skall vissa geografiska beteckningar behandlas som ursprungsbeteckningar när råvarorna till produkterna kommer från ett vidare geografiskt område än det område där produkterna bearbetas eller från ett annat område, om
- det område där råvarorna framställs är begränsat,
och - särskilda villkor gäller för framställningen av råvarorna,
och - kontroll har ordnats av att dessa villkor iakttas.
5. Vid tolkningen av punkt 4 får endast levande djur, kött och mjölk betraktas som råvaror. Bruk av andra råvaror kan godkännas i enlighet med det förfarande som stadgas i artikel 15.
6. För att kunna behandlas som ursprungsbeteckningar enligt punkt 4 måste beteckningarna i fråga godkännas eller redan vara godkända som ursprungsbeteckningar med nationellt skydd av ifrågavarande medlemsstat eller, om denna stat inte har ett sådant skyddssystem, ha vedertagen traditionell prägel och enastående rykte och anseende.
7. För att en beteckning skall behandlas som ursprungsbeteckning enligt punkt 4, måste ansökan om registrering inges inom två år från det att denna förordning trätt i kraft.
Artikel 3
1. Namn som har blivit generiska får inte registreras.
I denna förordning avses med namn som har blivit generiskt ett namn på en jordbruksprodukt eller ett livsmedel som, visserligen har samband med den ort eller den region där produkten eller livsmedlet från början framställdes eller marknadsfördes men har blivit den allmänna benämningen på produkten eller livsmedlet i fråga.
När det skall avgöras huruvida ett namn har blivit generiskt, skall hänsyn tas till alla faktorer, i synnerhet
- förhållandena i den medlemsstat som namnet kommer från och i de områden där produkten eller livsmedlet konsumeras,
- förhållandena i andra medlemsstater,
- berörd nationell lagstiftning och gemenskapslagstiftning.
När en ansökan om registrering avslås i enlighet med det förfarande som föreskrivs i artikel 6 och 7 av den anledningen att namnet har blivit generiskt, skall kommissionen offentliggöra beslutet i Europeiska gemenskapernas officiella tidning.
2. Ett namn får inte registreras som ursprungsbeteckning eller geografisk beteckning om det kommer i konflikt med namnet på en växtsort eller en djurras och därmed riskerar att vilseleda allmänheten om produktens verkliga ursprung.
3. Innan denna förordning träder i kraft skall rådet efter beslut med kvalificerad majoritet och på förslag av kommissionen upprätta och i Europeiska gemenskapernas officiella tidning offentliggöra en icke uttömmande vägledande förteckning över namn på jordbruksprodukter och livsmedel som omfattas av denna förordning och enligt punkt 1 skall betraktas som generiska och sålunda såsom icke registrerbara enligt denna förordning.
Artikel 4
1. För att en jordbruksprodukt eller ett livsmedel skall kunna få en skyddad ursprungsbeteckning (PDO) eller geografisk skyddad beteckning (PGI) måste produkten eller livsmedlet överensstämma med en produktspecifikation.
2. Produktspecifikationen skall omfatta bl. a. följande uppgifter:
a) Produktens eller livsmedlets benämning, inkl. ursprungsbeteckning eller geografisk beteckning.
b) En beskrivning av jordbruksprodukten eller livsmedlet, med uppgift i förekommande fall om råvarorna och de viktigaste fysiska, kemiska, mikrobiologiska och/eller organoleptiska egenskaperna hos produkten eller livsmedlet.
c) En definition av det geografiska området och i förekommande fall uppgifter som visar att kraven i artikel 2.4 är uppfyllda.
d) Uppgifter som styrker att produkten eller livsmedlet härstammar från det geografiska området, i den mening som avses i artikel 2.2 a respektive b.
e) En beskrivning av vilken metod som använts för framställning av jordbruksprodukten eller livsmedlet och i förekommande fall uppgift om den ursprungliga hävdvunna metoden i trakten.
f) Uppgifter som påvisar sambandet med den lokala omgivningen eller det geografiska ursprunget i den mening som avses i artikel 2.2 a respektive b.
g) Uppgifter om de kontrollorgan som föreskrivs i artikel 10.
h) Uppgifter om hur märkning sker med skyddad ursprungsbeteckning respektive geografisk beteckning eller jämbördiga traditionella nationella beteckningar.
i) De övriga uppgifter som föreskrivits av gemenskapen och/eller nationella stadganden.
Artikel 5
2. En grupp eller en fysisk eller juridisk person får ansöka om registrering endast av jordbruksprodukter eller livsmedel som denne själv producerar eller förädlar i den mening som avses i artikel 2.2 a eller b.
3. Ansökan om registrering skall innehålla den produktspecifikation som avses i artikel 4.
4. Ansökningen skall inges till den medlemsstat där det ifrågavarande geografiska området är beläget.
5. Medlemsstaten i fråga skall kontrollera att ansökningen uppfyller de krav som uppställts i denna förordning och om den finner att så är fallet tillställa kommissionen ansökan inklusive den produktspecifikation som avses i artikel 4 jämte de övriga handlingar varpå den byggt sitt beslut.
Om ansökningen avser ett namn på ett geografiskt område som sträcker sig in i en annan medlemsstat, skall denna senare medlemsstat tillfrågas innan beslut fattas.
1. Inom sex månader skall kommissionen genom en formell granskning kontrollera att registreringsansökningen innehåller alla de uppgifter som föreskrivs i artikel 4.
Kommissionen skall underrätta den berörda medlemsstaten om vad den därvid har funnit.
2. Om kommissionen med beaktande av vad som har framkommit vid den granskning som avses i punkt 1 finner att namnet är skyddsberättigat, skall den i Europeiska gemenskapernas officiella tidning offentliggöra sökandens namn och adress, produktens benämning, ansökningens huvudsakliga innehåll, hänvisningar till de nationella föreskrifter som kan finnas om produktens framställning och beredning och när så behövs motiveringen för sina slutsatser.
3. Om ingen invändning framställs till kommissionen i enlighet med artikel 7 skall namnet införas i ett register, "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar", som kommissionen skall föra och som skall uppta namn på de grupper och kontrollorgan som berörs.
4. Kommissionen skall i Europeiska gemenskapernas officiella tidning offentliggöra
- de namn som införts i registret,
- de ändringar i registret som företagits i enlighet med artikel 9 och 11.
5. Om kommissionen på basis av den granskning som föreskrivits i punkt 1 finner att namnet inte är skyddsberättigat, skall kommissionen i enlighet med det förfarande som föreskrivs i artikel 15 besluta att inte företa det offentliggörande som föreskrivs i punkt 2 i denna artikel.
Innan offentliggörande enligt punkt 2 och 4 och registrering enligt punkt 3 sker, får kommissionen inhämta yttrande av den kommitté som föreskrivs i artikel 15.
Artikel 7
1. Inom sex månader efter det offentliggörande i Europeiska gemenskapernas officiella tidning som avses i artikel 6.2, har varje medlemsstat rätt att framställa invändning mot registreringen.
2. Medlemsstaternas behöriga myndigheter skall se till, att alla personer som kan visa att de har ett lagligen berört ekonomiskt intresse tillåts ta del av ansökningen. Därutöver kan varje medlemsstat i enlighet med vad som eljest gäller i medlemsstaten i fråga bereda även andra parter med ett lagligen berört intresse åtkomst till ansökningen.
3. Varje lagligen berörd intresserad fysisk eller juridisk person får framställa invändning mot den begärda registreringen genom att inge en vederbörligen underbyggd skrivelse till den behöriga myndigheten i det medlemsstat där han bor eller verkar. Denna myndighet skall vidta de åtgärder som är nödvändiga för att pröva invändningen inom den fastställda tidsfristen.
4. En invändning skall upptas till behandling endast i något av följande fall:
- Invändningen visar att överträdelse skett av de villkor som avses i artikel 2.
- Invändningen visar att den föreslagna registreringen skulle äventyra överlevnaden för ett identiskt eller snarlikt namn eller varumärke eller för produkter som lagligen marknadsförs vid den tidpunkt då denna förordning offentliggörs i Europeiska gemenskapernas officiella tidning.
- Invändningen visar att det namn som registreringsansökningen avser är av generisk beskaffenhet.
5. När en invändning enligt punkt 4 är sådan att den skall tas upp till behandling, skall kommissionen uppmana de berörda medlemsstaterna att inom tre månader söka förlikning i enlighet med sina egna förfaranden. Därefter skall förfaras på endera av följande sätt.
a) Om förlikning har träffats, skall medlemsstaterna i fråga underrätta kommissionen om alla de faktorer som gjorde förlikningen möjlig jämte om sökandens och invändarens yttranden. När ingen ändring gjorts av de uppgifter som kommissionen har erhållit enligt artikel 5, skall kommissionen gå vidare i enlighet med artikel 6.4. Om någon ändring har gjorts skall kommissionen på nytt inleda det förfarande som föreskrivs i artikel 7.
b) Om ingen förlikning har träffats, skall kommissionen fatta beslut i enlighet med det förfarande som föreskrivs i artikel 15, med beaktande av traditionell skälig praxis och av den faktiska risken för förväxling. Om kommissionen beslutar att fullfölja registreringsförfarandet, skall den genomföra offentliggörande i enlighet med artikel 6.4.
Artikel 8
Beteckningarna PDO, PGI eller motsvarande traditionella nationella angivelser för skyddade ursprungsbeteckningar eller skyddade geografiska beteckningar får endast användas på jordbruksprodukter och livsmedel som uppfyller denna förordnings krav.
Artikel 9
Medlemsstaten i fråga får begära att produktspecifikationen ändras, t. ex. för att ta hänsyn till ny teknik och nya forskningsrön eller för att omdefiniera ett geografiskt område.
Artikel 6 skall därvid äga motsvarande tillämpning.
Kommissionen får dock i enlighet med det förfarande som föreskrivs i artikel 15 besluta att vid mindre ändringar inte tillämpa det förfarande som avses i artikel 6.
Artikel 10
1. Medlemsstaterna skall se till att, inom sex månader från det att denna förordning har trätt i kraft, kontrollorgan har upprättats med uppgift att säkerställa att jordbruksprodukter och livsmedel som bär en skyddad beteckning uppfyller de krav som fastställts i produktspecifikationen.
2. Ett kontrollorgan kan bestå av en eller flera för uppgiften utsedda kontrollmyndigheter och/eller privata organ som har godkänts för ändamålet av medlemsstaten. Medlemsstaterna skall tillställa kommissionen förteckningar på dessa myndigheter och/eller privata organ och deras respektive befogenheter. Kommissionen skall offentliggöra dessa uppgifter i Europeiska gemenskapernas officiella tidning.
3. Utsedda kontrollmyndigheter och godkända privata organ måste kunna garantera objektivitet och opartiskhet gentemot alla producenter och produktförädlare som underställs deras kontroll och ha ständig tillgång till den kvalificerade personal och de övriga resurser som behövs för att genomföra kontroller av jordbruksprodukter och livsmedel som bär en skyddad beteckning.
Om ett kontrollorgan anlitar ett annat organ för vissa kontrollåtgärder, måste detta senare kunna ge samma garantier. I sådana fall skall den utsedda myndigheter respektive det godkända privata organet fortfarande vara ansvarigt gentemot medlemsstaten för alla kontrollåtgärder.
Fr. o. m. den 1 januari 1988 måste ett privat organ för att kunna godkännas av en medlemsstat för de ändamål denna förordning avser, uppfylla de krav som fastställs i standarden EN 45011 av den 26 juni 1989.
4. Om en utsedd kontrollmyndighet respektive ett godkänt privat organ i en medlemsstat konstaterar att en jordbruksprodukt eller ett livsmedel som bär en skyddad ursprungsbeteckning där inte produktspecifikationens kriterier uppfylls, skall kontrollorganet vidta de åtgärder som är nödvändiga för att se till, att denna förordning följs. Kontrollorganet skall underrätta medlemsstaten om de åtgärder som vidtagits i samband med kontrollerna. Berörda parter måste underrättas om alla beslut som fattas.
5. En medlemsstat måste dra tillbaka godkännandet av ett kontrollorgan om de kriterier som avses i punkt 2 och 3 inte längre är uppfyllda. Medlemsstaten skall underrätta kommissionen härom, och denna skall i Europeiska gemenskapernas officiella tidning offentliggöra en reviderad förteckning över godkända kontrollorgan.
6. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att se till, att en producent som följer denna förordning har tillgång till kontrollsystemet.
7. Kostnaderna för de kontroller som föreskrivs i denna förordning skall bäras av de producenter som använder den skyddade beteckningen.
Artikel 11
1. Varje medlemsstat har rätt att framföra anmärkning om att ett villkor som ingår i en beteckningsskyddad jordbruksprodukts eller ett beteckningsskyddat livsmedels produktspecifikation inte är uppfylld.
2. Den medlemsstat som avses i punkt 1 skall rikta anmärkningen till den medlemsstat som är berörd. Denna skall granska anmärkningen och underrätta den klagande medlemsstaten om vad som framkommit och i förekommande fall om de åtgärder som har vidtagits.
3. Om avvikelser från produktspecifikationen upprepas och medlemsstaterna i fråga inte kunnat träffa förlikning skall en underbyggd ansökan inges till kommissionen.
4. Kommissionen skall granska denna ansökan genom att rådfråga de berörda medlemsstaterna. Kommissionen skall när så är lämpligt höra den kommitté som avses i artikel 15. Kommissionen skall därefter vidta de åtgärder som är nödvändiga. Till dessa kan höra att registreringen avförs.
Artikel 12
1. Utan att påverka tillämpningen av internationella överenskommelser kan denna förordning också tillämpas på en jordbruksprodukt eller ett livsmedel från tredje land under följande förutsättningar:
- Tredje land är berett att ge skydd likvärt det som är tillgängligt inom gemenskapen för motsvarande jordbruksprodukter eller livsmedel som härstammar från gemenskapen.
2. Om tredje lands skyddade beteckning sammanfaller med en skyddad beteckning i gemenskapen, skall registrering ske med vederbörlig hänsyn till lokalt och traditionellt språkbruk och till risken för förväxling i praktiken.
Bruk av sådana beteckningar skall vara tillåtet endast om produktens ursprungsland är klart och tydligt angivet i märkningen.
Artikel 13
1. Registrerade beteckningar skall skyddas mot följande.
a) Varje direkt eller indirekt kommersiellt bruk av den skyddade beteckningen för produkter som inte omfattas av registreringen i den mån dessa produkter är jämförbara med de produkter som har registrerats under beteckningen i fråga eller detta bruk av den skyddade beteckningen innebär att dennas anseende exploateras.
b) Varje obehörigt bruk, imitation eller anspelning, även när produktens verkliga ursprung anges eller det skyddade namnet har översatts eller åtföljs av uttryck som "stil", "typ", "metod", "sådan som tillverkas i", "imitation" eller dylikt.
c) Varje annan osann eller vilseledande uppgift om ursprung, härkomst, beskaffenhet eller väsentliga egenskaper hos produkten på dennas inre eller yttre förpackning, reklammaterial eller handlingar, liksom förpackning av produkten i behållare som är ägnad att inge en oriktig föreställning om produktens verkliga ursprung.
d) Annat beteende som är ägnat att vilseleda allmänheten om produktens verkliga ursprung.
När det i en registrerad beteckning ingår en benämning på en jordbruksprodukt eller ett livsmedel och denna benämning anses generisk, skall det inte anses strida mot reglerna i punkt a eller b ovan att använda denna generiska benämning om jordbruksprodukten eller livsmedlet i fråga.
2. Medlemsstaterna får dock låta nationella regler om rätt att bruka sådana beteckningar som avses i punkt 1 b bestå under högst fem år efter den dag denna förordning offentliggörs under förutsättning
- att produkterna lagligen har marknadsförts med användning av sådana uttryck under minst fem år före den dag denna förordning offentliggörs, och
- att märkningen klart anger produktens verkliga ursprung.
Detta undantag får dock inte leda till att produkterna fritt marknadsförs på en medlemsstats territorium där sådana uttryck är förbjudna.
3. Skyddade beteckningar får inte bli generiska.
Artikel 14
1. När en ursprungsbeteckning eller en geografisk beteckning registrerats i enlighet med denna förordning, skall ansökan om registrering av ett varumärke som svarar mot något av de fall som nämns i artikel 13 och som avser samma slags produkt, avslås om ansökningen ingivits efter dagen för det offentliggörande som avses i artikel 6.2.
Varumärkesregistrering som har skett i strid med vad som sägs i föregående stycke skall förklaras ogiltig.
Denna punkt skall också tillämpas när ansökan om registrering av varumärke ingivits före dagen för offentliggörande av den registreringsansökan som föreskrivs i artikel 6.2 under förutsättning att detta offentliggörande skedde innan varumärket registrerades.
Artikel 15
Kommissionen skall biträdas av en kommitté som skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen varvid medlemsstaternas röster skall vägas enligt nämnda artikel. Ordföranden får inte rösta.
Kommissionen skall själv anta förslaget till åtgärder om detta har tillstyrkts av kommittén.
Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte fattat något beslut inom tre månader från det att saken hänskjutits till rådet, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 16
Detaljregler för tillämpningen av denna förordning skall fastställas enligt det förfarande som föreskrivs i artikel 15.
Artikel 17
1. Inom sex månader efter det att denna förordning har trätt i kraft, skall medlemsstaterna meddela kommissionen vilka hos dem skyddade beteckningarna eller, vad gäller medlemsstater som saknar sådant skyddssystem, vilka inarbetade beteckningar de önskar registrera i enlighet med denna förordning.
2. I enlighet med det förfarande som föreskrivs i artikel 15 skall kommissionen registrera de av de beteckningar som avses i punkt 1 vilka uppfyller kraven i artikel 2 och 4. Artikel 7 skall inte vara tillämplig. Generiska beteckningar skall dock inte registrerats.
3. Medlemsstaterna får bibehålla det nationella skyddet för de beteckningar som de har meddelat i enlighet med punkt 1 intill dess att beslut om registrering i enlighet med denna förordning har fattats.
Artikel 18
Denna förordning träder i kraft tolv månader efter det att den har publicerats i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EEG) nr 2145/92 av den 29 juli 1992 om en omformulering vad avser de destinationszoner som skall användas vid fastställandet av exportbidrag, exportavgifter och vissa exportlicenser för spannmål och ris
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2727/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för spannmål(1), senast ändrad genom förordning (EEG) nr 1738/92(2), särskilt artikel 16.6 i denna,
med beaktande av rådets förordning (EEG) nr 1418/76 av den 21 juni 1976 om den gemensamma organisationen av marknaden för ris(3), senast ändrad genom förordning (EEG) nr 674/92(4), särskilt artikel 17.6 i denna, och
med beaktande av följande: I kommissionens förordning (EEG) nr 1124/77(5), senast ändrad genom förordning (EEG) nr 3049/89(6), fastställs de destinationszoner som skall användas vid fastställandet av exportbidrag och avgifter vid export av spannmål och ris.
De politiska förändringarna i östblocket, dvs. upplösningen av Sovjetunionen och Jugoslavien i oberoende stater, gör det nödvändigt att aktualisera den förteckning över destinationszoner som anges i bilagan till förordning (EEG) nr 1124/77. I den bilagan bör "Sovjetunionen" och "Jugoslavien" ersättas med namnen på de nybildade stater som tidigare ingick i Sovjetunionen och Jugoslavien. Dessutom bör det ske en omgruppering av staterna i område I, II, III och VIII när möjligheten nu bjuds.
Av hänsyn till tydligheten bör förordning (EEG) nr 1124/77 upphöra att gälla och dess bestämmelser bör införas i den här förordningen.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilagan till denna förordning anges de destinationszoner som skall användas vid fastställande av differentierade exportbidrag och exportavgifter för de produkter som förtecknas i artikel 1 punkt a, b och c i förordning (EEG) nr 2727/75 och i artikel 1 punkt a och b i förordning (EEG) nr 1418/76.
Förordning (EEG) nr 1124/77 skall upphöra att gälla.
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EEG) nr 2221/92 av den 31 juli 1992 om ändring av förordning (EEG) nr 1274/91 om tillämpningsföreskrifter för förordning (EEG) nr 1907/90 om vissa handelsnormer för ägg
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1907/90 av den 2 juni 1990 om vissa handelsnormer för ägg(1), särskilt artiklarna 10.3, 20.1 och 22.2 i denna, och med beaktande av följande:
I kommissionens förordning (EEG) nr 1274/91(2), senast ändrad genom förordning (EEG) nr 3540/91(3), fastställs de tillämpningsföreskrifter som krävs för införandet av sådana handelsnormer.
Erfarenheten har visat att bestämmelserna om frivillig angivelse av värpdagen bör ändras. Det bör entydigt klargöras att då värpdag anges, skall denna anges både på äggen och på förpackningarna. De villkor på vilka förpackningsanläggningar, som får äggen från produktionsenheter belägna på samma ställe, får ange värpdag bör bringas i överensstämmelse med de villkor som gäller för andra förpackningsanläggningar om man använder slutna behållare. Bestämmelser bör införas om märkning av ägg med värpdag då denna inte infaller på en arbetsdag.
Det valfria angivandet av produktionssystem bör begränsas till de termer som anges i förordning (EEG) nr 1274/91, med undantag för organiska eller biologiska produktionssystem. För att underlätta kontroller i hela gemenskapen bör förteckningarna över registrerade producenter utväxlas mellan medlemsstaterna och förpackningsanläggningar bör föra veckoregister över lager med klassificerade ägg.
De termer som används för livsmedelsindustrin bör harmoniseras.
Bestämmelserna om användningen av termen "extra" bör ändras i syfte att specificera villkoren för att denna term ska få förekomma på förpackningen.
En positiv vikttolerans bör införas för att säkerställa en rättvis konkurrens mellan aktörerna.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fjäderfäkött och ägg.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Artikel 1.6, andra strecksatsen, skall ersättas med följande text:
" - värpdagen skall anges på ägg vilka levereras av en produktionsenhet som är belägen på samma ställe som förpackningsanläggningen och vilka inte förpackas i slutna behållare, i vilket fall de skall klassificeras och förpackas på värpdagen, eller, om värpdagen inte infaller på en arbetsdag, den första därpå följande arbetsdagen."
1. Utöver förpackningsdagen får aktören vid förpackningstillfället ange rekommenderad sista försäljningsdag eller bäst före-dag på äggen eller på förpackningen, eller på bådadera.
2. Aktören får vid förpackningstillfället ange värpdagen på förpackningen, varvid värpdagen även skall anges på de ägg som förpackningen innehåller. Värpdagen får emellertid även stämplas på äggen på produktionsföretaget.
3. När datum som avses i denna artikel anges på ägg, och i fråga om värpdag även på förpackningen, skall en eller flera av de termer som anges i bilaga 1 användas.
4. De datum som avses i denna artikel skall anges med två siffergrupper som i följande ordning utvisar:
- dagen, från 01 till 31
- månaden, från 01 till 12."
Om värpdagen anges på ägg och äggförpackningar i enlighet med bestämmelserna i artikel 15, skall följande villkor gälla:
1 Förpackningsanläggningar skall föra separata register över
- namn och adress avseende de ägglevererande producenterna, som skall registreras efter det att den behöriga myndigheten i medlemsstaten har gjort ett kontrollbesök, och
- på begäran av denna myndighet, antalet värphönor som respektive producent håller.
2 De producenter som avses i punkt 1 skall därefter kontrolleras regelbundet. De skall föra löpande register över
- insättningsdagen, åldern vid insättning och antalet värphönor uppdelade efter hönshus,
- den dagliga äggproduktionen från varje hönshus,
- antalet ägg eller vikten på de ägg som levererats och på vilka man avser ange värpdagen, eller på vilka produktionsföretaget redan har stämplat värpdagen, uppdelade efter köpare, och med angivande av deras namn och adress samt förpackningsanläggningens nummer.
3 Ägg på vilka man avser ange värpdagen skall levereras till förpackningsanläggningar i slutna behållare, om inte produktionsenheten är belägen på samma ställe som förpackningsanläggningen. Leveranser av dessa ägg och av ägg på vilka produktionsföretaget redan har stämplat värpdagen, skall identifieras genom
- värpdagen,
- producentens namn, adress och nummer samt en kodad hänvisning till det hönshus från vilket äggen kommer,
Dessa uppgifter skall anges på behållaren och på de åtföljande dokumenten, som skall bevaras på förpackningsanläggningen i minst 6 månader.
4 De behållare som avses i punkt 3 skall öppnas på förpackningsanläggningen omedelbart innan klassificeringen påbörjas. Alla ägg från en enskild behållare skall klassificeras och förpackas utan avbrott. För ägg som skall märkas med värpdagen gäller att detta datum skall stämplas på äggen vid klassificeringen eller omedelbart efter denna.
5 För förpackningsanläggningar som får leveranser från egna produktionsenheter som är belägna på samma ställe och där äggen inte förpackats i slutna behållare, skall äggen
- stämplas med värpdagen samma dag som de värps medan ägg som värps på annan dag än arbetsdag får stämplas den första därpå följande arbetsdagen tillsammans med de ägg som värps denna dag, varvid den första dagen som inte är arbetsdag skall anges, eller
- klassificeras och förpackas i enlighet med föreskrifterna i artikel 1.6, eller
- levereras till andra förpackningsanläggningar eller industrin på värpdagen eller, om värpdagen infaller på en annan dag än arbetsdag, den första därpå följande arbetsdagen.
Om dessa förpackningsanläggningar även får ägg från externa producenter på vilka man inte avser ange värpdagen, skall dessa ägg lagras och hanteras separat. Dagligt register skall föras över uppsamling eller mottagning och klassificering av sådana ägg.
6 Förpackningsanläggningar skall föra separata register över
- de dagliga kvantiteter ägg som de mottar, uppdelade efter producenter och på vilka man avser ange värpdagen, eller på vilka produktionsföretaget redan har stämplat värpdagen, med angivande av producentens namn och adress samt registreringsnummer,
- daglig mängd ägg och äggens viktklass,
- antalet sålda ägg och/eller vikten på dessa, uppdelade efter viktklass och köpare, med angivande av köparens namn och adress.
7 De produktionsenheter och förpackningsanläggningar som avses i punkt 1 skall kontrolleras minst en gång varannan månad."
4 Artikel 18 skall ändras på följande sätt:
- I punkt 1 skall inledningsfrasen ersättas med följande:
"Inga andra termer än dem som anges här nedan får användas för att på ägg av klass 'A' och på små förpackningar innehållande sådana ägg ange de produktionssystem som avses i artikel 10.3 i förordning (EEG) nr 1907/90, med undantag för organiska och biologiska produktionssystem, och dessa termer får endast användas om de tillämpliga villkoren enligt bilaga 2 är uppfyllda."
- I punkt 1 skall det andra stycket utgå.
- Punkt 6 skall ersättas med följande:
"De förpackningsanläggningar som avses i punkt 2 skall föra separata register över den dagliga kvalitets- och viktklassificeringen samt försäljningen av ägg och små förpackningar som är märkta i enlighet med punkt 1, inbegripet köparens namn och adress, antalet förpackningar, antalet sålda ägg och/eller vikten på de ägg som sålts per viktklass och leveransdag, liksom veckoregister över lager med klassificerade ägg. I stället för att föra försäljningsregister kan de emellertid arkivera fakturor eller följesedlar på vilka finns angivet de uppgifter som avses i punkt 1."
5 Artikel 22.2 c skall ersättas med följande text:
"c) märkningen 'ÄGG TILL LIVSMEDELSINDUSTRIN', skriven med 2 cm höga bokstäver på ett eller flera av gemenskapens språk."
6 Artikel 24 skall ersättas med följande:
2. Om den banderoll eller etikett som avses i punkt 1 inte kan avlägsnas från förpackningen, skall banderollen eller förpackningen avlägsnas från försäljningsytan senast den sjunde dagen efter förpackningstillfället, varefter äggen skall förpackas på nytt.
3. Stora förpackningar som innehåller små förpackningar märks med texten `FÖRPACKNING INNEHÅLLANDE SMÅ FÖRPACKNINGAR MED "EXTRA" ÄGG`, med 2 cm höga versala bokstäver på ett eller flera av gemenskapens språk."
Med undantag för det fall som avses i artikel 13.3 i förordning (EEG) nr 1907/90, skall vid kontroll av ett parti ägg av klass `A` en tolerans medges med hänsyn till vikten per ägg. Ett sådant parti får innehålla högst 12 % ägg vars vikt gränsar till den på förpackningen angivna vikten och högst 6 % ägg av närmast lägre viktklass.
Om det kontrollerade partiet omfattar färre ägg än 180, skall ovan angivna procentsatser fördubblas."
8 Bilaga 1 skall ersättas med bilagan till denna förordning.
Artikel 2
Denna förordning träder i kraft den 1 augusti 1992. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EEG) nr 3224/92 av den 4 november 1992 om rättelse av förordning (EEG) nr 2342/92 om import av renrasiga avelsdjur av nötkreatur från tredje land och beviljande av exportbidrag för detta samt om upphävande av förordning (EEG) nr 1544/79
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött(1), senast ändrad genom förordning (EEG) nr 2066/92(2), särskilt artiklarna 10.5 och 18.6 i denna, och
med beaktande av följande: Genom kommissionens förordning (EEG) nr 2342/92(3) skärptes kontrollbestämmelserna i fråga om import från tredje land och beviljande av exportbidrag för renrasiga nötkreatur och upphävdes förordning (EEG) nr 1544/79.
Vid en genomgång visade det sig att den tyska utgåvan av förordningen inte återger de bestämmelser som förvaltningskommittén hade fått på remiss. Den tyska utgåvan bör därför ges ut i en helt ny version.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
(Berör endast den tyska utgåvan.)
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
RÅDETS BESLUT av den 8 februari 1993 om ingående av ett avtal om handel och ekonomiskt samarbete mellan Europeiska ekonomiska gemenskapen och Mongoliet (93/101/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 113 och 235 i detta,
med beaktande av kommissionens förslag,
Artikel 3
Kommissionen, biträdd av företrädare för medlemsstaterna, skall företräda gemenskapen i den gemensamma kommitté som inrättas i enlighet med artikel 13 i avtalet.
Artikel 4
Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
RÅDETS DIREKTIV 93/35/EEG av den 14 juni 1993 om ändring för sjätte gången av direktiv 76/768/EEG om tillnärmning av medlemsstaternas lagstiftning om kosmetiska produkter
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag(1),
i samarbete med Europaparlamentet(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: De juridiska oklarheterna i direktiv 76/768/EEG(4), särskilt i artiklarna 1 och 2, bör undanröjas.
Det har visat sig önskvärt att samla in uppgifter om de beståndsdelar som används i kosmetiska produkter, så att alla frågor som gäller användningen av dem och de därmed sammanhängande åtgärderna på gemenskapsnivå kan prövas på ett sätt som särskilt syftar till att upprätta en gemensam nomenklatur för beståndsdelar i kosmetiska produkter. Insamlingen av dessa uppgifter kan underlättas om kommissionen genomför en inventering av sådana beståndsdelar. Denna inventering skall vara vägledande och inte syfta till att upprätta en begränsande förteckning över ämnen för användning i kosmetiska produkter.
Större öppenhet krävs beträffande de beståndsdelar som används i kosmetiska produkter för att dessa skall kunna släppas ut på marknaden utan något föregående förfarande, för att de nödvändiga uppgifterna om slutprodukterna endast skall behövas finnas tillgängliga på tillverkningsstället eller på den plats dit de först importeras inom gemenskapen samt för att ge konsumenterna ökad information. En sådan öppenhet bör kunna uppnås om en kosmetisk produkts användningsområde och beståndsdelar anges på förpackningen. Om det av praktiska skäl är omöjligt att återge beståndsdelar och eventuella varningstexter beträffande användningen på behållaren eller den yttre förpackningen bör dessa uppgifter bifogas, så att konsumenterna får tillgång till all nödvändig information.
I fråga om färdiga kosmetiska produkter bör det fastställas vilka upplysningar som skall hållas tillgängliga för kontrollmyndigheterna på tillverkningsstället eller på den plats dit de först importerats inom gemenskapen. Dessa upplysningar skall innefatta alla nödvändiga uppgifter om identitet, kvalitet, säkerhet för människors hälsa och om de verkningar den kosmetiska produkten uppges ha.
I förebyggande syfte bör dock den behöriga myndigheten underrättas om tillverkningsplats och ges den information som är nödvändig för en snar och adekvat medicinsk behandling i händelse av betänkligheter.
Kommissionen bör ha befogenhet att ändra bilagorna 1 och 8 till direktiv 76/768/EEG med hänsyn till dessas informativa och tekniska karaktär.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 76/768/EEG ändras på följande sätt:
1. Artikel 1.1 skall ersättas med följande:
"1. Med kosmetisk produkt avses ämnen eller beredningar som är avsedda att appliceras på olika yttre partier av människokroppen (överhud, hår och hårbotten, naglar, läppar och yttre könsorgan) eller på tänder och slemhinnor i munhålan i uteslutande, eller huvudsakligt, syfte att rengöra eller parfymera dem eller förändra deras utseende och/eller korrigera kroppslukt och/eller skydda dem eller bibehålla dem i gott skick."
Kosmetiska produkter som släpps ut på marknaden inom gemenskapen får inte kunna skada människors hälsa vid normal eller rimligen förutsebar användning, varvid följande särskilt skall beaktas: presentationen av produkten, märkning, eventuella bruksanvisningar och anvisningar för kvittblivning samt eventuella andra anvisningar eller upplysningar som lämnas av tillverkaren eller hans representant eller av annan person som är ansvarig för att produkten släpps ut på gemenskapsmarknaden.
Det faktum att varningstexter av detta slag förekommer skall dock inte befria någon från skyldigheten att iaktta de övriga kraven i detta direktiv."
3. Följande led skall läggas till i artikel 4.1:
"i) beståndsdelar eller kombinationer av beståndsdelar som utprovats på djur efter den 1 januari 1998 för att uppfylla kraven i detta direktiv.
Om inte tillräckliga framsteg har uppnåtts i utvecklingen av tillfredsställande metoder som kan ersätta djurförsök, särskilt i sådana fall då alternativa provningsmetoder, trots att alla rimliga ansträngningar har gjorts, inte har kunnat valideras vetenskapligt som likvärdiga i fråga om skyddsnivån för konsumenterna med beaktande av OECD:s riktlinjer för toxicitetstester, skall kommissionen senast den 1 januari 1997 lämna förslag till åtgärder för att uppskjuta det datum då denna bestämmelse skall träda i kraft under rimlig tid, och i vart fall minst två år, i enlighet med det förfarande som fastställs i artikel 10. Kommissionen skall rådfråga Vetenskapliga kommittén för kosmetologi, innan den lämnar sådana förslag.
Kommissionen skall lämna en årlig rapport till Europaparlamentet och rådet om de framsteg som gjorts i utvecklingen, valideringen och det juridiska godkännandet av alternativa metoder som kan ersätta sådana som förutsätter djurförsök. Denna rapport skall innehålla exakta uppgifter om antal och slag av försök avseende kosmetika som utförts på djur. Medlemsstaterna skall vara skyldiga att samla in sådana uppgifter utöver den statistikinsamling som fastställs i direktiv 86/609/EEG om skydd av djur som används för försök och andra vetenskapliga ändamål. Kommissionen skall särskilt säkerställa att försöksmetoder, i vilka levande djur inte används, utvecklas, valideras och godkänns i lagstiftningen."
4. Följande artikel skall införas:
"Artikel 5a
1. Senast den 14 december 1994 skall kommissionen, med det förfarande som fastställs i artikel 10, ha sammanställt en inventering av de beståndsdelar som används i kosmetiska produkter, med stöd särskilt av information som lämnats av kosmetikaindustrin.
I denna artikel avses med beståndsdel i kosmetika varje kemiskt ämne eller beredning av syntetiskt eller naturligt ursprung, med undantag av parfym och aromatiska blandningar, som används i sammansättningen av kosmetiska produkter.
Denna inventering skall delas upp i två avdelningar: en för parfym och aromatiska råvaror och en för övriga ämnen.
2. Inventeringen skall innehålla uppgifter om
- varje beståndsdels identitet, särskilt dess kemiska benämning, CTFA-benämning, benämning i Europeiska farmakopén, den internationella generiska benämning som rekommenderas av världshälsoorganisationen, Einecs-, IUPAC-, CAS- och färgindexnummer samt den generiska benämning som avses i artikel 7.2,
- beståndsdelens normala funktion(er) i den färdiga produkten,
- då så är tillämpligt, begränsningar och villkor för användningen samt de varningstexter som skall förekomma i märkningen med hänvisning till bilagorna.
3. Kommissionen skall offentliggöra inventeringen och uppdatera den regelbundet med det förfarande som fastställs i artikel 10. Inventeringen skall vara vägledande, d. v. s. inte betraktas som en uttömmande förteckning över de ämnen som är godkända för användning i kosmetiska produkter."
5. I artikel 6.1 skall den inledande meningen ersättas med följande:
"1. Medlemsstaterna skall vidta alla de åtgärder som är nödvändiga för att försäkra sig om att kosmetiska produkter inte kan släppas ut på marknaden utan att följande information finns i outplånlig, lättläst och väl synlig skrift på behållaren och förpackningen. Den information som nämns i g behöver dock endast anges på förpackningen:"
6. Artikel 6.1 d skall ersättas med följande:
"d) Särskilda försiktighetsåtgärder som skall iakttas vid användning, i synnerhet sådana som anges i spalten "Villkor för användning och varningstexter som skall tryckas på etiketten" i bilagorna 3, 4, 6 och 7, som skall förekomma på behållare och förpackning tillsammans med eventuell information om försiktighetsåtgärder för kosmetiska produkter som används i yrkesmässig verksamhet, särskilt av frisörer. Om detta är ogörligt av praktiska skäl, skall denna information finnas på en bipacksedel, bifogad etikett, tejp eller kort och konsumenten skall hänvisas till denna information genom att antingen en förkortad upplysning eller den symbol som anges i bilaga 8 skall förekomma på behållaren och förpackningen."
7. Följande led f och g skall läggas till i artikel 6.1:
"f) Produktens funktion, om detta inte tydligt framgår av presentationen av produkten.
g) En förteckning över beståndsdelar i fallande ordning efter vikt då de tillsätts produkten. Denna förteckning skall föregås av ordet "innehåll". Om detta är ogörligt av praktiska skäl, skall uppgift om beståndsdelarna finnas på en bipacksedel, bifogad etikett, tejp eller kort och konsumenten skall hänvisas till denna information genom att antingen en förkortad upplysning eller den symbol som anges i bilaga 8 skall förekomma på behållaren och förpackningen."
Följande skall dock inte betraktas som beståndsdelar:
- Föroreningar i de använda råvarorna.
- Kompletterande tekniskt material som används vid framställningen men som inte förekommer i slutprodukten.
- Material av vilket endast oundgängligen nödvändiga kvantiteter används som lösningsmedel eller som bärare av parfym och aromatiska blandningar.
Parfym, aromatiska sammansättningar och råvaror till dessa skall betecknas med orden "parfym" eller "aromämne". Beståndsdelar som förekommer i lägre koncentrationer än 1 % får nämnas i valfri ordning efter de beståndsdelar som förekommer i högre koncentrationer. Färgämnen får upptas i valfri ordning efter övriga beståndsdelar med de färgindexnummer eller benämningar som används i bilaga 4.
I fråga om kosmetiska produkter som används i estetiskt syfte och som förekommer i flera nyanser får samtliga färgämnen som används i hela färgskalan nämnas i förteckningen, om uttrycket "kan innehålla" läggs till.
Beståndsdelar skall identifieras med den generiska benämning som avses i artikel 7.2 eller, om sådan saknas, med någon av de benämningar som avses i artikel 5a.2, första strecksatsen.
Kommissionen skall senast den 14 december 1994 i enlighet med förfarande i artikel 10 fastställa på vilka kriterier och villkor en tillverkare för att bevara affärshemligheter får ansöka om att befrias från kravet att uppta en eller flera beståndsdelar i den nämnda förteckningen."
8. Följande två stycken skall läggas till sist i artikel 6.1:
"Om det på grund av storlek eller form är ogörligt att uppta de uppgifter som avses i d och g på en bipacksedel skall dessa uppgifter förekomma på en etikett, en tejp eller ett kort som bipackas eller fästs på den kosmetiska produkten.
I fråga om tvål, kulor med badskum och andra små produkter vilkas storlek eller form gör det omöjligt att uppta de uppgifter som avses i g på en etikett, remsa, tejp eller kort eller på en bipacksedel skall dessa uppgifter skyltas i omedelbar närhet av den kosmetiska produktens säljbehållare."
9. Följande skall läggas till sist i artikel 6.3:
"Dessutom skall i varje omnämnande av djurförsök klart anges om de utförda försöken gällde slutprodukten och/eller dess beståndsdelar."
10. Artikel 7.2 skall ersättas med följande:
"2. De kan dock kräva att de uppgifter som anges i artikel 6.1 b-6.1 d och 6.1 f skall avfattas åtminstone på deras nationella eller officiella språk. De får även kräva att de uppgifter som anges i artikel 6.1 g skall avfattas på ett språk som konsumenterna kan förstå utan svårighet. Kommissionen skall därför i enlighet med förfarandet i artikel 10 fastställa en gemensam nomenklatur för beståndsdelar."
11. Artikel 7.3 skall ersättas med följande:
"3. Dessutom kan en medlemsstat kräva att snar och adekvat medicinsk behandling i händelse av betänkligheter skall göras möjlig genom att lämplig och tillräcklig information om vilka ämnen som ingår i den kosmetiska produkten finns tillgänglig för den behöriga myndigheten, som skall garantera att informationen endast används för att underlätta sådan medicinsk behandling.
Varje medlemsstat skall utse en behörig myndighet och sända uppgifter om detta till kommissionen, som skall offentliggöra denna information i Europeiska gemenskapernas officiella tidning."
12. Följande artikel skall införas:
"Artikel 7a
1. Tillverkaren eller dennes representant eller den person för vars räkning en kosmetisk produkt tillverkas eller den som är ansvarig för att en importerad kosmetisk produkt släpps ut på gemenskapsmarknaden skall i förebyggande syfte hålla följande information omedelbart tillgänglig för de behöriga myndigheterna i den medlemsstat det gäller på den adress som anges i märkningen enligt artikel 6.1 a:
a) Produktens kvalitativa och kvantitativa sammansättning. I fråga om parfymsammansättningar och parfymer: sammansättningens namn och kodnummer och uppgift om leverantören.
b) Fysikaliskkemiska och mikrobiologiska specifikationer för råvarorna och slutprodukten och renhetskriterier och kriterier för mikrobiologisk kontroll avseende den kosmetiska produkten.
c) Tillverkningsmetoden, som skall överensstämma med god tillverkningssed enligt gemenskapslagstiftning eller, om tillämplig sådan saknas, enligt lagstiftningen i den berörda medlemsstaten. Den person som är ansvarig för tillverkningen eller för den första importen till gemenskapen skall ha sådana yrkesmässiga kvalifikationer eller sådan erfarenhet som krävs i lagstiftning och praxis i den medlemsstat där tillverkningen eller den första importen sker.
d) Bedömning av slutproduktens säkerhet för människors hälsa. Tillverkaren skall därvid beakta beståndsdelens allmänna toxikologiska profil, dess kemiska struktur och dess exponeringsgrad.
Om samma produkt tillverkas på flera platser inom gemenskapen får tillverkaren välja att hålla informationen tillgänglig endast på en av dessa platser. Om så sker, samt om en begäran om detta riktas till honom i kontrollsyfte, skall han vara skyldig att ange den plats han valt till den eller de berörda tillsynsmyndigheterna.
e) Namn på och adress till den eller de experter som ansvarar för den bedömning som avses i d. Sådana experter skall ha ett examensbevis enligt definitionen i artikel 1 i direktiv 89/48/EEG i farmaci, toxikologi, dermatologi, medicin eller liknande ämne.
f) Tillgängliga uppgifter om icke önskvärda verkningar på människors hälsa som orsakas av användning av den kosmetiska produkten.
g) Bevisning för den verkan som den kosmetiska produkten uppges ha, om detta är motiverat med hänsyn till arten av denna verkan eller av produkt.
2. Den bedömning av säkerheten för människors hälsa som avses i punkt 1 d skall utföras enligt den princip om god laboratoriesed som fastställs i rådets direktiv 87/18/EEG av den 18 december 1986 om harmonisering av lagar och andra författningar om tillämpningen av principerna för god laboratoriesed och kontrollen av tillämpningen vid prov med kemiska ämnen(*).
3. Den information som avses i punkt 1 skall finnas tillgänglig på den berörda medlemsstatens nationella språk eller på ett språk som utan svårighet förstås av de behöriga myndigheterna.
4. Tillverkaren eller dennes representant eller den person för vars räkning en kosmetisk produkt tillverkas eller den som är ansvarig för att en importerad kosmetisk produkt släpps ut på gemenskapsmarknaden skall till den behöriga myndigheten i medlemsstaten meddela adressen till den plats där de kosmetiska produkterna tillverkas eller dit de först importeras inom gemenskapen, innan dessa produkter får släppas ut på gemenskapsmarknaden.
5. Medlemsstaterna skall utse de behöriga myndigheter som avses i punkterna 1 och 4 och sända uppgifter om dessa till kommissionen som skall offentliggöra denna information i Europeiska gemenskapernas officiella tidning.
13. Artikel 8.2 skall ersättas med följande:
"2. Den gemensamma nomenklaturen för beståndsdelar i kosmetiska produkter och de ändringar som, efter samråd med Vetenskapliga kosmetologikommittén, har bedömts nödvändiga för att anpassa bilagorna med hänsyn till den tekniska utvecklingen skall fastställas på lämpligt sätt med samma förfarande."
14. Bilaga 8, som återges i bilagan till detta direktiv, skall läggas till.
Artikel 2
1. Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att säkerställa att, från och med den 1 januari 1997, varken tillverkare eller importörer som är etablerade inom gemenskapen släpper ut kosmetiska produkter, som inte uppfyller kraven i detta direktiv, på marknaden.
2. Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att säkerställa att sådana produkter som avses i punkt 1 inte kan säljas eller avyttras till konsumenter efter den 31 december 1997.
Artikel 3
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 14 juni 1995. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar sådana bestämmelser skall dessa innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV 93/41/EEG av den 14 juni 1993 om upphävande av direktiv 87/22/EEG om tillnärmning av medlemsstaternas åtgärder vad gäller meddelande av försäljningstillstånd för högteknologiska läkemedel på marknaden, särskilt sådana som framställts genom bioteknologi
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag(1),
i samarbete med Europaparlamentet(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Bestämmelserna i direktiv 87/22/EEG(4) har nu ersatts med bestämmelserna i rådets förordning (EEG) nr 2309/93 av den 22 juli 1993 om gemenskapsförfaranden för godkännande för försäljning av och tillsyn över humanläkemedel och veterinärmedicinska läkemedel samt om inrättande av en europeisk läkemedelsmyndighet(5) och i rådets direktiv 88/182/EEG av den 22 mars 1988 om ändring av direktiv 83/189/EEG om ett informationsförfarande beträffande tekniska standarder och föreskrifter(6).
Direktiv 93/39/EEG(7) innehåller bestämmelser för den fortsatta administrationen av godkännanden för försäljning, som medlemsstaterna har meddelat efter yttrande från Kommittén för farmaceutiska specialiteter enligt direktiv 87/22/EEG.
Vidare innehåller direktiv 93/40/EEG(8) bestämmelser för den fortsatta administrationen av godkännanden för försäljning, som medlemsstaterna har meddelat efter yttrande från Kommittén för veterinärmedicinska läkemedel enligt direktiv 87/22/EEG.
Direktiv 87/22/EEG bör därför upphävas.
I rättssäkerhetens intresse bör bestämmelser fastställas för den fortsatta granskningen av ansökningar om godkännande för försäljning, som före den 1 januari 1995 föreläggs Kommittén för farmaceutiska specialiteter eller Kommittén för veterinärmedicinska läkemedel enligt direktiv 87/22/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 87/22/EEG skall upphöra att gälla med verkan från och med den 1 januari 1995.
Artikel 2
Ansökningar om godkännande för försäljning, som före den 1 januari 1995 har förelagts Kommittén för farmaceutiska specialiteter eller Kommittén för veterinärmedicinska läkemedel enligt artikel 2 i direktiv 87/22/EEG och beträffande vilka den berörda kommittén inte har avgivit något yttrande före den 1 januari 1995, skall anses uppfylla bestämmelserna i förordning (EEG) nr 2309/93.
Artikel 3
Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att följa detta direktiv med verkan från och med den 1 januari 1995. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av yttrandet från Ekonomiska och sociala kommittén(3), och
med beaktande av följande: I rådets direktiv 74/577/EEG(4) fastställs bestämmelser om bedövning av djur före slakt.
Den europeiska konventionen om skydd för slaktdjur godkändes på gemenskapens vägnar genom rådets beslut 88/306/EEG(5). Konventionens räckvidd är större än de befintliga gemenskapsbestämmelserna på området.
Nationella lagar om skydd av djur vid tidpunkten för slakt eller avlivning påverkar konkurrensvillkoren och följaktligen också hur den gemensamma marknaden för jordbruksprodukter fungerar.
Det är därför nödvändigt att fastställa gemensamma miniminormer för skydd av djur vid tidpunkten för slakt eller avlivning för att säkerställa en rationell utveckling av produktionen och för att underlätta genomförandet av den inre marknaden för djur och animalieprodukter.
Vid tidpunkten för slakt eller avlivning bör djur besparas onödig smärta och lidande.
Det är emellertid nödvändigt att tillåta att tekniska och vetenskapliga experiment utförs samt att ta hänsyn till de särskilda krav som vissa religiösa ceremonier ställer.
Bestämmelserna bör även säkerställa ett tillfredsställande skydd vid tidpunkten för slakt eller avlivning av djur som inte omfattas av konventionen.
I den förklaring om djurskydd som är knuten till slutakten av Fördraget om Europeiska unionen anmodar konferensen Europaparlamentet, rådet, kommissionen och medlemsstaterna att vid utformning och införande av gemenskapslagstiftning om den gemensamma jordbrukspolitiken fullt ut ta hänsyn till djurens behov av välbefinnande.
I samband med detta skall gemenskapens handlande vara i enlighet med subsidiarietsprincipen i artikel 3b i fördraget.
Direktiv 74/577/EEG bör upphöra att gälla.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Det skall inte gälla för
- tekniska eller vetenskapliga experiment i samband med förfarandena i punkt 1, vilka utförs under tillsyn av en behörig myndighet,
- djur som avlivas under kultur- eller sportarrangemang,
- vilda djur som avlivas i enlighet med artikel 3 i direktiv 92/45/EEG.
4. Fasthållning: Varje metod som tillämpas för att begränsa djurets rörelseförmåga i syfte att underlätta bedövning eller avlivning.
5. Bedövning: Varje metod som när den används på ett djur omedelbart försätter detta i ett tillstånd av medvetslöshet som varar tills döden inträder.
6. Avlivning: Varje metod som leder till att ett djur avlider.
7. Slakt: Avlivning av djur genom avblödning.
8. Behörig myndighet: Den centrala myndigheten i en medlemsstat som ansvarar för veterinärkontroller eller annan myndighet till vilken denna befogenhet har delegerats.
Den religiösa myndigheten i en medlemsstat för vars räkning slakt utförs skall emellertid ha befogenhet att tillämpa och övervaka särskilda bestämmelser i samband med slakt enligt vissa religiösa ceremonier. I fråga om dessa bestämmelser skall denna myndighet vara underställd den officiella veterinären, enligt definitionen i artikel 2 i direktiv 64/433/EEG.
Artikel 3
Djur skall skonas från all onödig upphetsning, smärta och lidande under förflyttning, uppstallning, fasthållning, bedövning, slakt eller avlivning.
KAPITEL II Krav för slakterier
Artikel 4
Slakterier, dvs. lokaler och utrustning, skall vara konstruerade på ett sådant sätt att djuren skonas från onödig upphetsning, smärta och lidande.
Artikel 5
1. Hovdjur, idisslare, svin, kaniner och fjäderfä som förs till slakterier för att slaktas skall
a) förflyttas och, om nödvändigt, uppstallas i enlighet med bilaga A,
b) fasthållas i enlighet med bilaga B,
c) bedövas före slakt eller avlivas omedelbart i enlighet med bilaga C,
d) avblödas i enlighet med bilaga D.
2. Kraven i punkt 1 c skall inte tillämpas beträffande djur som slaktas med särskilda metoder som krävs i samband med vissa religiösa ceremonier.
3. Medlemsstaternas behöriga myndigheter kan under iakttagande av fördragets allmänna bestämmelser vad gäller anläggningar som omfattas av undantag enligt artikel 4 och artikel 13 i direktiv 64/433/EEG, artikel 4 i direktiv 91/498/EEG och artikel 7 och artikel 18 i direktiv 71/118/EEG, avstå från att tillämpa punkt 1 a vad gäller kreatur, och från punkt 1 a samt metoderna för bedövning och slakt i bilaga C vad gäller fjäderfä, kaniner, svin, får och getter, under förutsättning att kraven som fastställs i artikel 3 uppfylls.
Artikel 6
1. Instrument, fasthållningsanordningar och annan utrustning och anläggningar som används vid bedövning och avlivning skall utformas, konstrueras, underhållas och användas på ett sådant sätt att bedövningen eller avlivningen sker snabbt och effektivt i enlighet med bestämmelserna i detta direktiv. Den behöriga myndigheten skall kontrollera att instrument, fasthållningsanordningar och annan utrustning som används vid bedövning eller avlivning är i överensstämmelse med ovanstående principer och skall regelbundet kontrollera att de är i gott skick och kan uppfylla denna målsättning.
2. Lämplig reservutrustning och reservinstrument skall finnas på slaktplatsen att användas i nödsituationer. De skall underhållas och besiktigas regelbundet.
Artikel 7
Förflyttning, uppstallning, fasthållning, slakt eller avlivning av djur får endast utföras av personer som har nödvändiga kunskaper och yrkesskicklighet för att utföra arbetet humant och effektivt i enlighet med kraven i detta direktiv.
Den behöriga myndigheten skall säkerställa att personer som arbetar med slaktning har nödvändig yrkesskicklighet och yrkesmässigt kunnande.
Artikel 8
Den behöriga myndigheten skall ansvara för att det utförs besiktningar och kontroller av slakterier och skall vid alla tidpunkter ha fritt tillträde till slakteriernas alla delar för att säkerställa att bestämmelserna i detta direktiv efterlevs. Besiktningarna och kontrollerna får dock genomföras samtidigt som kontroller som genomförs i andra syften.
KAPITEL III Slakt och avlivning utanför slakterier
Artikel 9
1. När de djur som avses i artikel 5.1 slaktas utanför slakterier skall artikel 5.1 b, 5.1 c och 5.1 d tillämpas.
2. Medlemsstaterna kan emellertid bevilja undantag från punkt 1 beträffande fjäderfä, kaniner, svin, får och getter som slaktas eller avlivas utanför slakterier av sin ägare för dennes personliga bruk, under förutsättning att artikel 3 efterlevs och att svin, får och getter först blir bedövade.
Artikel 10
1. När de djur som avses i artikel 5.1 skall slaktas eller avlivas vid sjukdomsbekämpning skall detta utföras i enlighet med bilaga E.
2. Djur som uppföds för pälsens skull skall avlivas i enlighet med bilaga F.
3. Dagsgamla överskottskycklingar enligt definitionen i artikel 2.3 i direktiv 90/539/EEG, och embryon i kläckningsavfall skall avlivas så snabbt som möjligt i enlighet med bilaga G.
Artikel 11
Artikel 9 och artikel 10 skall inte tillämpas beträffande djur som i en nödsituation måste avlivas omedelbart.
Artikel 12
Skadade eller sjuka djur måste slaktas eller avlivas på stället. Den behöriga myndigheten kan emellertid tillåta transport av skadade eller sjuka djur för slakt eller avlivning under förutsättning att detta inte innebär ytterligare lidande för djuren.
KAPITEL IV Slutbestämmelser
Artikel 13
1. Rådet skall, om nödvändigt, genom kvalificerad majoritet på kommissionens förslag anta andra bestämmelser om skydd av djur vid tidpunkten för slakt eller avlivning än de som omfattas av detta direktiv.
2. a) Bilagorna till detta direktiv skall ändras av rådet på förslag från kommissionen i enlighet med förfarandet i punkt 1, i synnerhet för att anpassa dem till den tekniska och vetenskapliga utvecklingen.
b) Kommissionen skall vidare senast den 31 december 1995 överlämna en rapport till rådet, som utarbetats på grundval av ett yttrande från Vetenskapliga veterinärmedicinska kommittén, tillsammans med relevanta förslag beträffande användningen av
- pistol med skarp ammunition, där kulan drivs in i hjärnan, eller andra gaser än de som avses i bilaga C eller kombinationer av dessa som används vid bedövning, särskilt koldioxid vid bedövning av fjäderfä,
- andra gaser än de som avses i bilaga C eller kombinationer av dessa som används vid avlivning,
- varje annan vetenskapligt erkänd metod för bedövning eller avlivning.
Rådet skall ta ställning till dessa förslag med kvalificerad majoritet.
c) Trots vad som sägs i a, och senast den 31 december 1995, skall kommissionen i enlighet med förfarandet i artikel 16 lämna in en rapport till Ständiga veterinärkommittén, som utarbetats på grundval av ett yttrande från Vetenskapliga veterinärmedicinska kommittén, tillsammans med relevanta förslag för fastställande av
i) nödvändig strömstyrka och varaktighet vid bedövning av de olika berörda arterna,
ii) nödvändig gaskoncentration och exponeringstid vid bedövning av de olika berörda arterna.
d) I avvaktan på att b och c skall genomföras skall nationella bestämmelser på området fortsätta att gälla under iakttagande av fördragets allmänna bestämmelser.
Artikel 14
1. Kommissionens experter får, i den mån detta är nödvändigt för att säkerställa en enhetlig tillämpning av detta direktiv, utföra kontroller på plats. De kan i detta syfte kontrollera ett representativt urval av anläggningar för att säkerställa att den behöriga myndigheten kontrollerar att dessa anläggningar uppfyller kraven i detta direktiv.
Kommissionen skall underrätta medlemsstaterna om resultaten av kontrollerna.
2. De kontroller som avses i punkt 1 skall utföras i samarbete med den behöriga myndigheten.
3. Den medlemsstat på vars område kontrollen genomförs skall ge experterna all nödvändig hjälp i deras tjänsteutövning.
4. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 16.
Artikel 15
Vid besiktning av slakterier eller anläggningar i tredje land vilka har bemyndigats eller skall bemyndigas att exportera till gemenskapen i enlighet med gemenskapsbestämmelser, skall kommissionens experter säkerställa att de djur som avses i artikel 5 har slaktats under villkor som minst garanterar samma humana behandling som den som fastställs i detta direktiv.
För att kött skall få importeras från tredje land skall det hälsointyg som åtföljer köttet kompletteras med ett intyg som visar att ovanstående krav har uppfyllts.
Artikel 16
1. Vid hänvisning till det förfarande som fastställs i denna artikel skall frågan utan dröjsmål hänskjutas till Ständiga veterinärkommittén av dess ordförande, antingen på dennes eget initiativ eller på anmodan av en representant för en medlemsstat.
2. Kommissionens representant skall förelägga kommittén ett utkast till de åtgärder som skall vidtas. Kommittén skall avge ett yttrande om utkastet inom den tid som dess ordförande fastställt beroende på hur brådskande ärendet är. Yttrandet skall avges av den majoritet som fastställs i artikel 148.2 i fördraget beträffande beslut som rådet skall anta på kommissionens förslag. Medlemsstaternas representanters röster skall vägas på det sätt som anges i samma artikel. Ordföranden skall inte delta i omröstningen.
3. a) Kommissionen skall anta de avsedda åtgärderna när de är förenliga med kommitténs yttrande.
b) Om de avsedda åtgärderna inte är förenliga med kommitténs yttrande, eller om inget yttrande avges, skall kommissionen utan dröjsmål förelägga rådet ett förslag om de åtgärder som skall vidtas. Rådet skall fatta beslut med kvalificerad majoritet.
Om rådet inte har fattat beslut före utgången av en period på tre månader från den dag då saken förelades dem, skall de föreslagna åtgärderna antas av kommissionen utom då rådet har uttalat sig mot de aktuella åtgärderna med enkel majoritet.
Artikel 17
Direktiv 74/577/EEG skall upphöra att gälla från och med den 1 januari 1995.
Artikel 18
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar, inklusive sanktionsåtgärder, som är nödvändiga för att följa detta direktiv den 1 januari 1995. De skall genast underrätta kommissionen om detta.
När medlemsstaterna antar dessa lagar och andra författningar skall de innehålla en hänvisning till detta direktiv eller vid offentliggörandet åtföljas av en sådan hänvisning. Närmare regler för denna hänvisning skall fastställas av medlemsstaterna.
2. Från och med den dag som fastställs i punkt 1 får medlemsstaterna, under iakttagande av fördragets allmänna bestämmelser, inom sina områden upprätthålla eller tillämpa mer restriktiva bestämmelser än de som omfattas av detta direktiv. De skall underrätta kommissionen om alla sådana åtgärder.
3. Medlemsstaterna skall meddela kommissionen ordalydelsen i de viktigaste nationella bestämmelserna som de antar på det område som omfattas av detta direktiv.
Artikel 19
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EEG) nr 752/93 av den 30 mars 1993 om tillämpningsföreskrifter för rådets förordning (EEG) nr 3911/92 om export av kulturföremål
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3911/92 av den 9 december 1992(1) om export av kulturföremål, särskilt artikel 7 i denna,
efter samråd med Rådgivande kommittén för kulturföremål, och
med beaktande av följande: Det är nödvändigt att anta tillämpningsföreskrifter för förordning (EEG) nr 3911/92, som bl.a. föreskriver inrättandet av en exportlicensordning för vissa kategorier av kulturföremål som anges i bilagan till den förordningen.
För att säkerställa att de exportlicenser som föreskrivs i nämnda förordning är enhetliga är det nödvändigt att fastställa regler för upprättandet, utfärdandet och användningen av formulären. Det bör därför utarbetas en förlaga till en sådan licens.
Exportlicenser måste upprättas på ett av gemenskapens officiella språk.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
AVSNITT I Formulär för licens
2. Användning av exportlicens får inte på något sätt påverka de förpliktelser som är förbundna med exportformaliteter eller därtill knutna handlingar.
Artikel 3
1. Formuläret skall tryckas på vitt träfritt skrivpapper som väger minst 55 gram per kvadratmeter.
2. Formulären skall vara 210 × 297 mm.
3. Formulären skall tryckas och fyllas i på ett av gemenskapens officiella språk, bestämt av de behöriga myndigheterna i den utfärdande medlemsstaten. De behöriga myndigheterna i den medlemsstat där formuläret uppvisas får begära att det översätts till det officiella språket eller ett av de officiella språken i den medlemsstaten. I så fall skall översättningskostnaderna bäras av innehavaren av licensen.
4. Medlemsstaterna skall vara ansvariga
- för att låta trycka formulären som skall vara försedda med tryckeriets namn och adress eller identifieringsmärke,
- för att vidta nödvändiga åtgärder för att undvika att formulären förfalskas. De sätt för identifiering som antas av medlemsstaterna för detta ändamål skall anmälas till kommissionen för att vidarebefordras till de behöriga myndigheterna i de andra medlemsstaterna.
5. Formulären skall företrädesvis fyllas i på mekanisk eller elektronisk väg. Ansökan får emellertid fyllas i läsligt för hand; i det senare fallet skall det fyllas i med bläck och med tryckbokstäver. Oavsett vilken metod som används får formulären inte innehålla raderingar, överskrivna ord eller andra ändringar. AVSNITT II
Användning av licens
Artikel 4
1. Utan att det påverkar tillämpningen av punkt 3 skall en särskild exportlicens utfärdas för varje sändning av kulturföremål.
2. I punkt 1 förstås med sändning antingen ett enda kulturföremål eller ett antal kulturföremål.
3. När en sändning innehåller ett antal kulturföremål är det de behöriga myndigheterna som skall bestämma om en eller flera exportlicenser bör utfärdas för sändningen i fråga.
Artikel 5
Formulären skall bestå av tre exemplar, varav
- ett exemplar märkt nr 1 skall utgöra ansökan,
- ett exemplar märkt nr 2 är avsett för innehavaren av licensen,
- ett exemplar märkt nr 3 skall återsändas till den utfärdande myndigheten.
Artikel 6
1. Den sökande skall fylla i fält 1, 3 -19 A och 21 och om nödvändigt 23 på ansökan och de andra exemplaren. Medlemsstaterna får emellertid föreskriva att endast ansökan behöver fyllas i.
2. Ansökan skall åtföljas av
- dokumentation som innehåller alla relevanta upplysningar om kulturföremålen och deras rättsliga status vid tidpunkten för ingivande av ansökan, i förekommande fall med hjälp av stödjande handlingar (fakturor, expertvärderingar etc),
3. De behöriga myndigheterna får för att utfärda en exportlicens kräva att de kulturföremål som skall exporteras visas upp.
4. Om tillämpningen av punkterna 2 och 3 orsakar kostnader skall dessa bäras av den som ansöker om exportlicens.
5. För att exportlicens skall beviljas skall de vederbörligen ifyllda formulären läggas fram för de behöriga myndigheter som utsetts av medlemsstaterna enligt artikel 2.2 i grundförordningen. När myndigheten har beviljat exportlicens skall exemplar 1 behållas av den myndigheten och de återstående exemplaren återsändas till innehavaren av exportlicensen eller till dennes representant.
Artikel 7
Följande skall framläggas till stöd för exportdeklarationen:
- Det exemplar som är avsett för innehavaren av licensen.
- Det exemplar som skall återsändas till den utfärdande myndigheten.
Artikel 8
2. Efter att ha fyllt i fält 19 B skall det tullkontor som är behörigt att ta emot exportdeklarationen återsända det exemplar som är avsett för innehavaren av licensen till deklaranten eller dennes representant.
3. Det exemplar av formuläret som skall återsändas till den utfärdande myndigheten skall åtfölja sändningen till kontoret vid platsen för utförsel ur gemenskapen. Tullkontoret skall om nödvändigt fylla i fält 5 i formuläret och stämpla i fält 22 och återsända det till innehavaren av exportlicensen eller dennes representant för att formuläret skall kunna sändas tillbaka till den utfärdande myndigheten.
Artikel 9
1. Exportlicensens giltighetstid får inte överstiga tolv månader räknat från utfärdandedagen.
2. I fråga om ansökan om temporär export får de behöriga myndigheterna specificera den tidsfrist inom vilken kulturföremålen skall återimporteras till den utfärdande medlemsstaten.
3. När en exportlicens löper ut utan att ha använts skall innehavaren omedelbart återsända de exemplar han har i sin ägo till den utfärdande myndigheten.
Artikel 10
Bestämmelserna i avsnitt IX i kommissionens förordning (EEG) nr 1214/92(2) och artikel 22.6 i bilaga 1 till Konventionen om ett gemensamt transiteringsförfarande som slöts den 20 maj 1987(3) mellan gemenskapen och EFTA-länderna skall gälla när varor som omfattas av denna förordning passerar genom ett EFTA-lands territorium vid förflyttning inom gemenskapen.
Artikel 11
Denna förordning träder i kraft den 1 april 1993.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EEG) nr 1785/93 av den 30 juni 1993 om de avgörande faktorerna för tillämpning av jordbruksomräkningskurser inom textilsektorn
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas avseende den gemensamma jordbrukspolitiken(1), särskilt artikel 6.2 i denna, och
med beaktande av följande: Enligt rådets förordning (EEG) nr 845/72 av den 24 april 1972 om särskilda åtgärder för att främja silkesodling(2), senast ändrad genom förordning (EEG) nr 2059/92(3), beviljas stöd för de lådor med silkesfjärilsägg som ger upphov till en lyckad maskodling. Den tidpunkt när det ekonomiska målet har uppnåtts kan därför normalt anses vara den 1 augusti varje regleringsår. Detta datum kan därför användas som den avgörande händelsen för den jordbruksomräkningskurs som skall tillämpas på stöd för odling av silkesmask.
Enligt kommissionens förordning (EEG) nr 876/75 av den 3 april 1975 om den avgörande faktorn för utbetalning av för lin och hampa samt silkesodling(4), kommissionens förordning (EEG) nr 1426/86 av den 14 maj 1986 om den avgörande faktorn för rätt till stöd för privat lagring av lin- och hampfibrer(5) och artikel 15 i kommissionens förordning (EEG) nr 1201/89 av den 3 maj 1989 om tillämpningsföreskrifter för stödsystemet för bomull(6), senast ändrad genom förordning (EEG) nr 2328/92(7), fastställs de avgörande faktorerna för jordbruksomräkningskursen på grundval av kriterier och rättsliga bestämmelser som genomgående har ändrats i samband med den nya agromonetära ordning som infördes genom förordning (EEG) nr 3813/92. I kommissionens förordning (EEG) nr 1068/93 av den 30 april 1993 om närmare föreskrifter för fastställande och tillämpning av jordbruksomräkningskurserna(8) fastställs på grundval av de nya bestämmelserna de avgörande händelserna för jordbruksomräkningskurserna, bland annat de som gäller ovannämnda belopp.
Enligt artikel 10.1 och 10.2 i förordning (EEG) nr 1068/93 skall de avgörande faktorerna för minimipriset och för stödet till bomull vara de som anges i artikel 15 i förordning (EEG) nr 1201/89. Det bör dock ges möjlighet att förutfastställa jordbruksomräkningskurserna för stödet.
Enligt artikel 11.1 i förordning (EEG) nr 1068/93 skall den jordbruksomräkningskurs som gäller i början av regleringsåret tillämpas på hektarstödet för lin och hampa. I artikel 10.3 i samma förordning fastställs att den avgörande faktorn för stöd för privat lagring av lin- och hampfibrer skall vara den dag när kontraktet för varje enskilt parti börjar gälla. Förordningarna (EEG) nr 876/75 och (EEG) nr 1426/86 kan därför upphävas.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för lin och hampa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
I artikel 15 i förordning (EEG) nr 1201/89 skall följande stycke läggas till:
Artikel 3
Förordning (EEG) nr 876/75 och förordning (EEG) nr 1426/86 skall upphöra att gälla.
Artikel 4
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EEG) nr 2040/93 av den 27 juli 1993 om fastställande av storleken på produktionsstöd för matpotatis på Madeira och storleken på produktionsstöd för sättpotatis och endiver på Azorerna, som fastställts i ecu av rådet och reducerats till följd av centralkursjusteringar
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas avseende den gemen-samma jordbrukspolitiken(1), särskilt artikel 9.1 i denna, och
med beaktande av följande: I kommissionens förordning (EEG) nr 3824/92 av den 28 december 1992 om ändring av priser och belopp fastställda i ecu till följd av centralkursjusteringarna(2), senast ändrad genom förordning (EEG) nr 1663/93(3), fastställs förteckningen över de priser och belopp som från början av regleringsåret 1993/944, skall divideras med koefficienten 1,013088, som fastställs i kommissionens förordning (EEG) nr 537/93(4), ändrad genom förordning (EEG) nr 1331/93(5), som ett led i ordningen för automatisk avveckling av negativa monetära avvikelser. I enlighet med artikel 2 i förordning (EEG) nr 3824/92 skall de sänkta priserna och beloppen fastställas och anges för varje ifrågavarande sektor.
I rådets förordning (EEG) nr 1600/92(6), ändrad genom kommissionens förordning (EEG) nr 3714/92(7), fastställs ett stöd för den lokala produktionen av matpotatis på Madeira och för sättpotatis och endiver på Azorerna. Dessa stödbelopp bör justeras enligt ovan nämnda bestämmelser.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för utsäde.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Det stöd som avses i artiklarna 16 och 27 i förordning (EEG) nr 1600/92, och som har sänkts i enlighet med artikel 2 i förordning (EEG) nr 3824/92, fastställs till 494 ecu per hektar.
Artikel 2
RÅDETS FÖRORDNING (EEG) nr 2617/93 av den 21 september 1993 om ändring av förordning (EEG) nr 1907/90 om vissa handelsnormer för ägg
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2771/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för ägg(1), särskilt artikel 2.2 i denna,
med beaktande av kommissionens förslag, och
med beaktande av följande: I förordning (EEG) nr 1907/90(2) föreskrivs vissa handels-normer för ägg.
Bestämmelserna i fråga om direkta leveranser från producenter till förpackningsanläggningar, vissa marknader och livsmedelsindustriföretag bör också gälla sådana leveranser till andra industriföretag.
Leveranser av bortsorterade ägg bör begränsas till sådana livs-medelsindustriföretag som godkänts i enlighet med rådets direktiv 89/437/EEG av den 20 juni 1989 om hygien-och hälsoproblem som påverkar tillverkningen och utsläppandet på marknaden av äggprodukter(3), för att säkerställa att sådana ägg hanteras korrekt.
Det bör klargöras att valfria märkningar på äggförpackningar avsedda som reklam får innehålla symboler och syfta på såväl ägg som andra varor.
Erfarenheten har visat att bestämmelserna om datummärkning på ägg av klass A och på de äggförpackningar som innehåller sådana ägg bör ändras så att det krävs ett obligatoriskt angivande av datum för minsta hållbarhetstid på samma sätt som för andra livsmedel, i överensstämmelse med rådets direktiv 79/112/EEG av den 18 december 1978 om tillnärmning av medlemsstaternas lagstiftning om märkning, presentation och reklam i fråga om livsmedel(4). I syfte att underlätta kontroll bör även förpackningen till importerade ägg av klass A ha en märkning som anger förpackningsdatum.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 1907/90 ändras på följande sätt:
2. Artikel 4.1 a skall ersättas med följande:
"a) ägg till någon annan än uppsamlare, förpacknings-anläggningar, de marknader som avses i artikel 2.2 a, livsmedelsindustriföretag som godkänts i enlighet med direktiv 89/437/EEG och andra företag än livsmedelsindustrin."
3. I artiklarna 6.1 och 8.3 skall ordet "livsmedelsindustri" ersättas med "livsmedelsindustriföretag som godkänts i enlighet med direktiv 89/437/EEG."
4. Artikel 7 a skall ersättas med följande:
"a) Datum för minsta hållbarhetstid 'bäst-före-datum`".
5. Artikel 10.1 a skall ersättas med följande:
"a) Namnet eller firmabeteckningen och adressen till det företag som har förpackat äggen eller låtit förpacka dem; namn, firmanamn eller varumärke som används av det företaget och som kan vara ett varumärke som används gemensamt av ett antal företag, får anges om det inte innehåller någon kommentar eller symbol som är oförenlig med denna förordning i fråga om äggens kvalitet eller färskhet, typen av produktionssystem som används vid produktionen eller äggens ursprung."
6. Artikel 10.1 e skall ersättas med följande:
"e) Datum för minsta hållbarhetstid 'bäst-före-datum` åtföljt av lämpliga förvaringsinstruktioner för ägg av klass A, och förpackningsdag för ägg av andra klasser."
7. Artikel 10.2 e skall ersättas med följande:
"e) Kommentarer eller symboler avsedda att främja försäljningen av ägg eller andra varor, under förutsättning att dessa kommentarer eller symboler är utformade på ett sådant sätt att det inte är sannolikt att de vilseleder köparen."
8. Artikel 13.2 skall ersättas med följande:
"2. När det gäller lösviktsförsäljning av ägg skall kontrollnumret på den förpackningsanläggning som klassificerade äggen anges eller, i fråga om importerade ägg, det tredje land där äggen har sitt ursprung liksom datum för minsta hållbarhetstid, åtföljt av lämpliga förvaringsinstruktioner."
9. Artikel 15 b ee skall ersättas med följande:
Kommissionen skall i enlighet med förfarandet i artikel 17 i förordning (EEG) nr 2771/75 föreskriva de övergångs-bestämmelser som behövs för genomförandet av den här förordningen, särskilt i fråga om de bestämmelser som gäller användningen av befintligt förpackningsmaterial.
Artikel 3
Denna förordning träder i kraft den 1 december 1993.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EEG) nr 2847/93 av den 12 oktober 1993 om införande av ett kontrollsystem för den gemensamma fiskeripolitiken
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag(),
med beaktande av Europaparlamentets yttrande(),
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
För att nå detta mål måste ett sådant system innehålla föreskrifter för kontroll av att åtgärderna för bevarande och förvaltning av fiskeresurserna, strukturåtgärderna och åtgärderna avseende en gemensam marknadsorganisation genomförs; det måste också innehålla vissa bestämmelser om sanktioner ifall åtgärderna inte genomförs omfattande hela fiskerisektorn, från producenten till konsumenten.
Det är bara om de berörda parterna erkänner att systemet är berättigat som det kan ge önskat resultat.
Även om det i första hand är medlemsstaterna som ansvarar för kontrollen, bör kommissionen också försöka se till att medlemsstaterna opartiskt kontrollerar och förebygger överträdelser. Kommissionen bör därför ges de finansiella medel samt rättskipnings- och lagstiftningsmedel som tillåter den att utföra detta uppdrag så effektivt som möjligt.
Erfarenheten från tillämpningen av rådets förordning (EEG) nr 2241/87 av den 23 juli 1987 om vissa åtgärder för kontroll av fisket() visar att det är nödvändigt att skärpa kontrollen av tillämpningen av föreskrifterna för bevarande av fiskeresurserna.
Det krävs att de inblandade parterna inom fiskerinäringen tar på sig ett ökat ansvar för att se till att åtgärderna för bevarande och förvaltning av fiskeresurserna genomförs.
Politiken avseende förvaltning av fiskeresurserna, som särskilt bygger på totala tillåtna fångstmängder (TAC), fångstkvoter och tekniska åtgärder bör också omfatta förvaltning av fiskeansträngningen, som innebär att fiskeverksamheten och fiskekapaciteten övervakas.
För att kunna övervaka alla fångster och landningar måste medlemsstaterna kontrollera den verksamhet som gemenskapens fiskefartyg bedriver i alla marina farvatten, samt all annan verksamhet som är förknippad med denna och har på så vis möjlighet att granska tillämpningen av bestämmelserna för den gemensamma fiskeripolitiken.
Det är av avgörande betydelse att medlemsstaterna samarbetar under inspektionerna av fiskeverksamheten ute till havs för att dessa skall bli så effektiva och ekonomiskt försvarbara som möjligt, särskilt under de inspektioner som företas i farvattnen utanför en medlemsstats jurisdiktion eller överhöghet.
I samband med införandet av den gemensamma fiskeripolitiken är det nödvändigt med åtgärder för att kontrollera de fartyg som för ett tredje lands flagg och befinner sig i gemenskapens farvatten. Det behövs särskilt ett system som gör det möjligt att följa fartygens rörelser och motta meddelanden om vilka arter som fartyget har ombord, utan att detta påverkar rätten till oskadlig genomfart genom territorialvattnet och friheten att navigera i fiskezonen om 200 sjömil.
Genom att medlemsstaterna i samarbete med kommissionen genomför pilotprojekt som kan tillämpas på vissa kategorier av fartyg, kan rådet före den 1 januari 1996 avgöra om det finns anledning att införa ett övervakningssystem via satellit eller något annat system.
Förvaltningen av fisket genom fastställande av TAC:er förutsätter en ingående kännedom om fångsternas sammansättning. En sådan kännedom behövs också för övriga förfaranden enligt förordning (EEG) nr 3760/92. Det kräver att befälhavaren på varje fiskefartyg för loggbok.
Landningsmedlemsstaten måste kunna övervaka landningarna på sitt territorium; därför bör de fiskefartyg som är registrerade i andra medlemsstater informera landningsmedlemsstaten om sin avsikt att landa på dess territorium.
Det är viktigt att vid landningen närmare klargöra och bekräfta uppgifterna i loggböckerna; de personer som har hand om landningen och avsättningen av fångsterna måste därför anmäla vilka mängder som landats, lastats om, bjudits ut till försäljning eller köpts.
För att kunna undanta små fiskefartyg från skyldigheten att föra loggbok eller fylla i en landningsdeklaration, för vilka en sådan skyldighet skulle innebära en oproportionerlig börda i förhållande till deras fiskekapacitet, är det nödvändigt att varje medlemsstat kan kontrollera dessa fartygs verksamhet genom att införa en provtagningsplan.
För att säkerställa att gemenskapens handelsåtgärder och åtgärder för bevarande respekteras bör alla fiskeprodukter som importeras till gemenskapen eller landas där, fram till dess att den första försäljningen äger rum, åtföljas av ett transportdokument som anger deras ursprung.
Begränsningar av fångsterna måste förvaltas såväl på medlemsstats- som gemenskapsnivå. Medlemsstaterna bör registrera landningarna och anmäla dem till kommissionen på elektronisk väg. Undantag från denna skyldighet måste därför kunna göras för små mängder som landas, emedan en elektronisk överföring i sådana fall skulle innebära en oproportionerligt stor administrativ och ekonomisk belastning för medlemsstaternas myndigheter.
För att säkerställa att alla de utnyttjade resurserna bevaras och förvaltas kan bestämmelserna om loggbok, landnings- och försäljningsdeklarationer samt upplysningar om omlastningar och registrering av fångster utvidgas till att omfatta sådana bestånd som inte omfattas av någon TAC eller kvot.
Medlemsstaterna måste hållas underrättade om resultaten av sina fartygs verksamhet i vatten som lyder under tredje lands jurisdiktion eller på internationellt vatten. Skyldigheten att föra loggbok och avge landnings- och omlastningsdeklaration bör därför också gälla för befälhavarna på dessa fartyg. De uppgifter som medlemsstaterna samlar in bör översändas till kommissionen.
För att hantera insamlingen och behandlingen av uppgifterna behöver databaser upprättas som särskilt gör det möjligt att samköra data. Kommissionen och dess inspektörer bör därför ha tillgång till dessa databaser på elektronisk väg för att kunna granska dem.
Om det finns nätredskap med olika maskstorlek ombord kan det inte säkert garanteras att bestämmelserna om hur fiskeredskapen får användas följs om de inte blir föremål för ytterligare kontroll. För vissa former av fiske kan det vara lämpligt att införa speciella regler som till exempel ennätsregeln.
När en medlemsstats kvot förbrukats, eller när själva TAC:en är förbrukad, måste kommissionen fatta beslut om förbud mot fiske.
Det är nödvändigt att gottgöra den skada som en medlemsstat lidit som inte har förbrukat sin kvot, tilldelning eller andel av ett bestånd eller grupp av ett bestånd när fisket stoppas till följd av att en TAC är förbrukad. Av denna anledning bör ett kompensationssystem införas.
Om de ansvariga för fiskefartygen inte följer bestämmelserna i denna förordning bör dessa fartyg bli föremål för ytterligare kontroll med hänsyn till bevarandet.
För att säkerställa att de åtgärder som vidtagits förvaltas effektivt är det nödvändigt att införa en deklarationsordning som överensstämmer med de mål och strategier som fastställs i artikel 8 i förordning (EEG) nr 3760/92, vilken är tillämplig på en medlemsstat som överskridit sin kvot.
Ett av huvudsyftena med den gemensamma fiskeripolitiken är att anpassa fångstkapaciteten till de tillgängliga resurserna. Enligt artikel 11 i förordning (EEG) nr 3760/92 är det rådets uppgift att lägga fast mål och strategier för en omläggning av fiskeansträngningen. Det är också nödvändigt att se till att åtgärderna rörande den gemensamma marknadsorganisationen respekteras, särskilt av de personer som berörs av dem. Det är därför av avgörande betydelse att varje medlemsstat, utöver de finansiella kontroller som redan finns föreskrivna i gemenskapsbestämmelserna, gör tekniska kontroller för att se till att de av rådet fastställda bestämmelserna följs.
Det är nödvändigt att fastställa allmänna regler så att gemenskapens inspektörer som utsetts av kommissionen kan se till att gemenskapsbestämmelserna tillämpas enhetligt och granska de kontroller som gjorts av medlemsstaternas behöriga myndigheter.
För att säkerställa granskningens objektivitet är det viktigt att gemenskapens inspektörer under vissa omständigheter får göra självständiga inspektioner utan att förvarna för att granska de kontroller som gjorts av de behöriga myndigheterna i medlemsstaterna. Sådana inspektioner får aldrig omfatta kontroll av privatpersoner.
De åtgärder som vidtas till följd av överträdelserna kan variera från ett land till ett annat, vilket får fiskarna att känna sig orättvist behandlade. Frånvaron av avskräckande straffpåföljder i några medlemsstater minskar kontrollernas effektivitet. Följaktligen bör medlemsstaterna vidta nödvändiga icke diskriminerande åtgärder för att förebygga och beivra oegentligheter, särskilt genom att införa ett straffsystem som effektivt berövar lagöverträdarna det ekonomiska utbytet av överträdelserna.
Om en landningsmedlemsstat inte effektivt beivrar oegentligheter kommer det att försvaga flaggmedlemsstatens möjligheter att se till att föreskrifterna för bevarande och förvaltning av fiskeresurserna följs. Det är därför nödvändigt att fastställa bestämmelser om att olovliga fångster skrivs av från landningsmedlemsstatens kvot, om denna stat underlåter att vidta effektiva åtgärder.
Medlemsstaterna bör regelbundet avlägga rapport till kommissionen om sin inspektionsverksamhet och om vilka åtgärder som vidtas vid brott mot gemenskapens bestämmelser.
För vissa åtgärder som avses i denna förordning är det lämpligt att fastställa tillämpningsföreskrifter.
Det bör säkerställas att de uppgifter som samlas in inom ramen för denna förordning behandlas konfidentiellt.
Denna förordning bör inte inverka på sådana nationella kontrollbestämmelser som, även om de hör till dennas tillämpningsområde, sträcker sig utanför förordningens minimiföreskrifter, förutsatt att de nationella bestämmelserna är förenliga med gemenskapsrätten.
Förordning (EEG) nr 2241/87 bör upphävas, med undantag av artikel 5 som fortfarande gäller fram till dess att de listor som avses i artikel 6.2 i denna förordning antagits.
Det är nödvändigt att fastställa en övergångsperiod för genomförandet av särbestämmelserna i vissa artiklar för att de behöriga myndigheterna i medlemsstaterna skall kunna införa och anpassa sina förfaranden till den nya förordningens krav.
Bestämmelserna i vissa artiklar bör träda i kraft den 1 januari 1999 i den mån de berör fisket i Medelhavet, där den gemensamma fiskeripolitiken ännu inte är helt genomförd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- åtgärderna för bevarande och förvaltning av fiskeresurserna,
- strukturåtgärderna,
- åtgärderna avseende den gemensamma organisationen av marknaden,
samt vissa bestämmelser om hur verkningsfulla de sanktioner bör vara som skall tillämpas om ovan nämnda åtgärder inte genomförs.
2. I detta syfte skall varje medlemsstat i enlighet med gemenskapsbestämmelserna vidta nödvändiga åtgärder för att säkerställa systemets effektivitet. Den skall ställa tillräckliga medel till sina behöriga myndigheters förfogande, så att de kan genomföra den inspektion och kontroll som fastställs i denna förordning.
Artikel 2
1. För att säkerställa att alla gällande föreskrifter om åtgärder för bevarande och kontroll följs skall varje medlemsstat inom sitt territorium och de marina farvatten som lyder under dess överhöghet eller jurisdiktion övervaka fisket och den därmed förbundna verksamheten. Medlemsstaten skall inspektera fiskefartygen och undersöka all verksamhet rörande landning, försäljning, transport och lagring av fisk samt registrering av landningar och försäljning, och kan på så sätt granska tillämpningen av denna förordning.
2. De fiskefartyg som kan bedriva fiske under ett tredje lands flagg och fiska i vatten som lyder under en medlemsstats överhöghet eller jurisdiktion skall ingå i ett system, där fartygets rörelser kan följas och uppgifter kan fås om vilka fångster som finns ombord.
Medlemsstaterna skall anmäla till kommissionen vilka åtgärder som vidtagits för att säkerställa att dessa förfaranden följs.
3. Varje medlemsstat skall kontrollera sina fartygs verksamhet utanför gemenskapens fiskezon, om en sådan kontroll krävs för att säkerställa att de gemenskapsbestämmelser som gäller i dessa farvatten efterlevs.
4. För att inspektionen skall bli så effektiv och ekonomisk som möjligt skall medlemsstaterna samordna sin kontrollverksamhet. De kan därför utarbeta gemensamma inspektionsprogram som gör det möjligt att kontrollera gemenskapens fiskefartyg i de i punkterna 1 och 3 nämnda farvattnen. Medlemsstaterna skall vidta sådana åtgärder som gör det möjligt för deras behöriga myndigheter och kommissionen att regelbundet och ömsesidigt hålla varandra underrättade om den erfarenhet som vunnits.
Artikel 3
1. För att åstadkomma större effektivitet i övervakningen av fiskeverksamheten skall rådet före den 1 januari 1996 i enlighet med det förfarande som fastställs i artikel 43 i fördraget besluta om i vilken utsträckning och när ett system bör införas för fortlöpande kontroll av gemenskapens fiskefartygs position från en land- eller satellitbaserad basstation med dataöverföring via satellit.
2. För att utvärdera vilken teknik som skall användas och vilka fartyg som skall omfattas av nämnda system skall medlemsstaterna i samarbete med kommissionen genomföra vissa pilotprojekt före den 30 juni 1995. Medlemsstaterna skall därför se till att ett system för fortlöpande lokalisering av vissa kategorier av fiskefartyg inom gemenskapen införs, som arbetar från en land- eller satellitbaserad basstation och använder sig av satellitkommunikation för dataöverföringen.
Medlemsstaterna får samtidigt genomföra pilotprojekt för att utvärdera användningen av automatiska anordningar för positionsregistrering.
3. När de pilotprojekt som avses i punkt 2 genomförs skall den medlemsstat vars flagg fartyget för eller i vilken fartyget är registrerat vidta nödvändiga åtgärder för att säkerställa att de data som översänds till eller inhämtas från dess fiskefartyg registreras i maskinläsbar form, oberoende av i vilka vatten fartygen fiskar eller i vilken hamn de befinner sig.
Om fiskefartygen befinner sig i farvatten som lyder under en annan medlemsstats överhöghet eller jurisdiktion skall flaggmedlemsstaten se till att de behöriga myndigheterna i den berörda medlemsstaten omgående underrättas om detta.
1. Varje medlemsstat skall själv och för egen räkning genomföra den i artikel 2 angivna inspektionen och övervakningen med hjälp av ett inspektionssystem som medlemsstaten själv fastlägger.
Medlemsstaterna skall när de utför de uppgifter som anförtrotts dem se till att de i artikel 2 angivna bestämmelserna och åtgärderna respekteras. De skall dessutom vid inspektionen undvika att göra onödiga ingrepp i den normala fiskeverksamheten. De skall också se till att ingen diskriminering sker med avseende på de sektorer och fartyg som tas ut för inspektion.
2. De ansvariga för de fiskefartyg, lokaler eller transportmedel som skall inspekteras skall medverka till att underlätta den inspektion som skall genomföras i överensstämmelse med punkt 1.
Artikel 5
I enlighet med förfarandet i artikel 36 kan tillämpningsföreskrifter antas för artiklarna 2, 3 och 4, speciellt med avseende på
a) identifiering av officiellt utsedda inspektörer, inspektionsfartyg och andra liknande inspektionsmedel som en medlemsstat kan utnyttja,
b) det förfarande som inspektörer och befälhavare på fiskefartyg skall följa när en inspektör vill göra ett besök ombord,
c) det förfarande som inspektörer som har gått ombord på ett fiskefartyg skall följa när de inspekterar fartyget, dess fiskeredskap eller fångster,
d) den rapport som inspektörerna skall sammanställa efter varje inspektion ombord,
e) märkning och identifiering av fiskefartygen och deras fiskeredskap,
f) utfärdande av intyg för fiskefartygens egenskaper avseende fiskeaktiviteter,
g) registrering av uppgifter rörande fiskefartygens position och överföring av dessa uppgifter till medlemsstaterna och kommissionen,
h) det system som skall tillämpas med avseende på de fiskefartyg som för ett tredje lands flagg för att ge upplysning om deras rörelser och vilka fiskeprodukter de har ombord.
Artikel 6
1. Befälhavarna på sådana fiskefartyg inom gemenskapen som fiskar arter ur ett bestånd eller en grupp av bestånd skall föra loggbok, i vilken de skall ange vilka fångstmängder som finns ombord av varje art, datum och plats (statistisk rektangel ICES) för dessa fångster och vilken typ av fiskeredskap som använts.
2. De arter som i enlighet med punkt 1 skall antecknas i loggboken är de arter som omfattas av TAC:er eller kvoter samt övriga arter som finns på de listor som rådet antar med kvalificerad majoritet på förslag av kommissionen.
3. Befälhavarna på gemenskapens fiskefartyg skall i loggböckerna skriva in vilka mängder som fångats i havet, datum och plats för dessa fångster samt de i punkt 2 avsedda arterna. De mängder som kastats överbord kan registreras i uppskattningssyfte.
4. Befälhavarna på gemenskapens fiskefartyg skall undantas från kraven i punkterna 1 och 3 om fartygets största längd understiger 10 m.
5. Rådet kan på kommissionens förslag med kvalificerad majoritet besluta om andra undantag än det som avses i punkt 4.
6. Varje medlemmstat skall genom stickprovskontroller kontrollera verksamheten hos de fiskefartyg som är undantagna från de krav som anges i punkterna 4 och 5 för att säkerställa att dessa fartyg följer gällande gemenskapsbestämmelser.
Varje medlemsstat skall därför utarbeta en provtagningsplan, som skall lämnas till kommissionen. Resultaten av de kontroller som görs skall regelbundet meddelas kommissionen.
7. Befälhavarna på gemenskapens fiskefartyg skall registrera de uppgifter som avses i punkterna 1 och 3, antingen i maskinläsbar form eller på papper.
8. Närmare bestämmelser skall antas för tillämpningen av denna artikel enligt det förfarande som anges i artikel 36, i vissa speciella fall med en annan geografisk grundval än den statistiska ICES-rektangeln.
Artikel 7
1. Den befälhavare på ett fiskefartyg inom gemenskapen som önskar använda landningsställen vilka är belägna i en annan medlemsstat än flaggmedlemsstaten skall minst två timmar i förväg till de behöriga myndigheterna i denna medlemsstat anmäla
- landningsplatsen eller landningsplatserna och den beräknade ankomsttiden,
- vilka mängder av varje art som skall landas.
2. Den befälhavare enligt punkt 1 som underlåter att göra anmälan kan bli utsatt för lämpliga sanktioner av de behöriga myndigheterna.
3. Kommissionen kan enligt det förfarande som anges i artikel 36 undanta vissa kategorier av fiskefartyg inom gemenskapen från den skyldighet som avses i punkt 1 under en begränsad tid, som kan förnyas, eller fastställa en annan anmälningsfrist, där hänsyn bland annat skall tas till avståndet mellan fiskebankarna, landningsplatserna och de hamnar i vilka fartygen ifråga är registrerade eller förtecknade.
Artikel 8
1. Befälhavarna på sådana fiskefartyg inom gemenskapen som har en största längd av minst 10 m, eller deras ställföreträdare, skall efter varje resa inom 48 timmar efter landningen lämna in en deklaration till de behöriga myndigheterna i den medlemsstat där landningen äger rum. Befälhavaren är ansvarig för deklarationens riktighet, som minst skall innehålla uppgift om de landade mängderna av varje art som avses i artikel 6.2 och i vilket område de fångats.
2. Rådet kan med kvalificerad majoritet på förslag av kommissionen besluta om att utsträcka den skyldighet som avses i punkt 1 till sådana fartyg som har en största längd av mindre än 10 m. Rådet kan också med kvalificerad majoritet på förslag av kommissionen besluta om undantag från skyldigheten i punkt 1 för vissa kategorier av fartyg med en största längd av minst 10 m, vilka bedriver viss typ av fiskeverksamhet.
3. Varje medlemsstat skall genom stickprovskontroller övervaka den verksamhet som bedrivs av de fiskefartyg som är undantagna från kraven i punkt 1 för att säkerställa att dessa fartyg följer gällande bestämmelser inom gemenskapen.
Varje medlemsstat skall därför utarbeta en provtagningsplan och sända den till kommissionen. Resultaten av de kontroller som görs skall regelbundet meddelas kommissionen.
4. Tillämpningsföreskrifter för denna artikel skall antas i enlighet med det förfarande som fastställs i artikel 36.
Artikel 9
1. De auktionsinrättningar eller andra av medlemsstaterna bemyndigade organ som ansvarar för den första saluföringen av de fiskeprodukter som landas i en medlemsstat skall vid första försäljningstillfället lämna in en avräkningsnota, för vars riktighet dessa organ skall ansvara, till de behöriga myndigheterna i den medlemsstat på vars territorium den första saluföringen sker. Detta ansvar omfattar bara den information som avses i punkt 3.
2. Om den första saluföringen av de fiskeprodukter som landats i en medlemsstat inte sker på det sätt som fastställs i punkt 1 får köparen inte föra bort de landade fiskeprodukterna innan en avräkningsnota lämnats in till de behöriga myndigheterna eller andra godkända organ i den medlemsstat på vars territorium saluföringen ägt rum. Köparen är ansvarig för riktigheten av de uppgifter enligt punkt 3 som avräkningsnotan innehåller.
3. De avräkningsnotor som avses i punkterna 1 och 2 skall minst innehålla följande uppgifter:
- Individuell storlek eller vikt för varje art, samt kvalitet, produktform och färskhet.
- Pris och mängd av varje art vid första försäljningstillfället och, i förekommande fall, beroende på de olika arternas storlek eller vikt, kvalitet, produktform och färskhet.
- Destinationen för de eventuella produkter som dragits tillbaka från marknaden (biprodukter, mänsklig komsumtion, förädling).
- Såväl säljarens som köparens namn.
- Dag och plats för försäljningen.
4. Dessa avräkningsnotor skall fyllas i och översändas i enlighet med landningsmedlemsstatens lagstiftning på sådant sätt och enligt sådana försäljningsvillkor att följande uppgifter kan inkluderas:
- Distriktsbeteckning och namn på det fiskefartyg som landat ifrågavarande produkter.
- Namnet på fartygets ägare eller befälhavare.
- Hamn och datum för landningen.
5. Avräkningsnotorna som avses i punkt 1 skall inom 48 timmar efter försäljningen översändas till medlemsstaternas behöriga myndigheter eller andra bemyndigade organ, antingen på elektronisk väg eller på papper.
6. De behöriga myndigheterna skall behålla ett exemplar av varje avräkningsnota under en tid av ett år räknat från början av det år som följer på året för registreringen av den information som översänts till de behöriga myndigheterna.
7. Kommissionen kan i enlighet med förfarandet i artikel 36 bevilja undantag från skyldigheten att presentera avräkningsnotan för medlemsstaternas behöriga myndigheter eller andra behöriga organ för de fiskprodukter som landats från vissa kategorier av gemenskapens fiskefartyg med en största längd av mindre än 10 m.
Dessa undantag får bara beviljas om medlemsstaten ifråga har infört ett godtagbart kontrollsystem.
8. En köpare som köper produkter som inte saluförs vidare utan endast används för privat konsumtion skall undantas från kraven i punkt 2.
9. Närmare bestämmelser för tillämpningen av denna artikel skall antas i enlighet med det förfarande som anges i artikel 36.
Artikel 10
1. a) De fiskefartyg som för ett tredje lands flagg eller är registrerade i ett tredje land, och som har tillstånd att bedriva fiske i sådana marina farvatten som lyder under en medlemsstats överhöghet eller jurisdiktion, skall föra loggbok, i vilken den i artikel 6 angivna informationen skall införas.
b) Varje medlemsstat skall se till att befälhavaren på ett fiskefartyg som för ett tredje lands flagg eller är registrerat i ett tredje land, eller dennes ställföreträdare, vid landningen lämnar in en deklaration till myndigheterna i den medlemsstat vars landningsplatser han utnyttjar med uppgift om landade mängder och datum och plats för varje fångst; för deklarationens riktighet ansvarar befälhavaren eller dennes ställföreträdare.
c) Befälhavaren på ett fiskefartyg som för ett tredje lands flagg eller är registrerat i ett tredje land skall minst 72 timmar i förväg anmäla till de behöriga myndigheterna i den medlemsstat vars landningsplatser han önskar utnyttja vid vilken tid han avser att anlöpa landningshamnen.
Befälhavaren får inte landa fångster om medlemsstatens behöriga myndigheter inte bekräftat mottagandet av förhandsanmälan.
Medlemsstaterna skall fastställa tillämpningsföreskrifter för punkt 1 c och anmäla dem till kommissionen.
2. Kommissionen får enligt förfarandet i artikel 36, under en begränsad tid som kan förlängas, undanta vissa kategorier av fiskefartyg från ett tredje land från deras förpliktelse enligt punkt 1 c, eller fastställa en annan anmälningsfrist, där hänsyn tas till bland annat avstånden mellan fiskebankarna, landningsplatserna och hamnarna i vilka fartygen ifråga är registrerade eller förtecknade.
3. Punkterna 1 och 2 skall gälla utan att de påverkar tillämpningen av de fiskeavtal som ingåtts mellan gemenskapen och vissa tredje länder.
Artikel 11
1. Utan att det påverkar tillämpningen av artiklarna 7, 8 och 9, skall befälhavaren på ett gemenskapsfartyg som
- omlastar valfria fångstmängder ur ett bestånd eller en grupp av bestånd inom en TAC eller kvot till ett annat fartyg, nedan kallat "mottagarfartyg", oberoende av omlastningsplatsen, eller
- direktlandar sådana fångstmängder utanför gemenskapens territorium,
vid omlastningen eller landningen underrätta den medlemsstat vars flagg hans fartyg för eller i vilket fartyget är registrerat om gällande arter och mängder och datumet för omlastningen eller landningen samt fångstplatsen med hänvisning till det minsta område för vilket en TAC eller kvot fastställts.
2. Senast 24 timmar innan en omlastning eller serie omlastningar som äger rum i en hamn eller i sådana marina farvatten som lyder under en medlemsstats överhöghet eller jurisdiktion inleds, eller när de avslutats, skall mottagarfartygets befälhavare underrätta denna medlemsstats behöriga myndigheter om storleken på de fångster ur ett bestånd eller en grupp av bestånd som omfattas av en TAC eller en kvot, vilka befinner sig ombord på detta fartyg.
Befälhavaren på mottagarfartyget skall förvara uppgifterna om storleken på de fångster ur ett bestånd eller en grupp av bestånd inom en TAC eller kvot vilka tagits emot vid en omlastning, datumet när de togs emot och fartyget som lastade om fångsterna till mottagarfartyget. Denna skyldighet skall anses vara uppfylld när kopior förvaras av de omlastningsdeklarationer som är utfärdade i enlighet med de närmare bestämmelserna om medlemsstaternas registrering av uppgifter om fiskefångster.
När en omlastning eller en rad omlastningar ägt rum skall mottagarfartygets befälhavare inom 24 timmar lämna in dessa uppgifter till ovannämnda behöriga myndigheter.
Befälhavaren på mottagarfartyget skall också förvara uppgifterna om vilka fångstmängder ur ett bestånd eller en grupp av bestånd inom en TAC eller kvot som mottagarfartyget lastat om till ett tredje fartyg, samt underrätta ovannämnda behöriga myndigheter om denna omlastning minst 24 timmar innan den äger rum. Efter omlastningen skall befälhavaren underrätta nämnda myndigheter om vilka mängder som lastats om.
Befälhavarna på mottagarfartyget och ovannämnda tredje fartyg skall låta de behöriga myndigheterna kontrollera riktigheten av de uppgifter som krävs enligt denna punkt.
3. Medlemsstaterna skall vidta nödvändiga åtgärder för att kontrollera riktigheten av de uppgifter som erhållits enligt punkterna 1 och 2 och i förekommande fall överlämna dessa uppgifter och resultaten av granskningen till den eller de medlemsstater där mottagarfartyget och det fartyg varifrån omlastning sker är registrerade, eller vars flagg de för.
4. Punkterna 2 och 3 skall även tillämpas på ett mottagarfartyg som för ett tredje lands flagg eller är registrerat i ett tredje land.
Artikel 12
Om omlastningen eller landningen beräknas ske mer än 15 dagar efter fångsten skall de upplysningar som krävs enligt artiklarna 8 och 11 senast 15 dagar efter fångsten överlämnas till de behöriga myndigheterna i den medlemsstat där fartyget är registrerat eller vars flagg det för.
Artikel 13
1. Alla fiskeprodukter som importeras till gemenskapen eller landas där, såväl icke beredda som beredda ombord, vilka transporteras till en annan plats än landnings- eller införselplatsen, skall åtföljas av ett dokument utfärdat av transportören fram till dess att den första försäljningen ägt rum.
2. Detta dokument skall innehålla uppgifter om
a) försändelsens ursprung (fartygets namn och distriktsbeteckning),
b) försändelsens eller försändelsernas destination och transportmedlet,
c) fiskmängderna (i kg beredd vikt) för varje transporterad art, namnet på avsändaren och platsen och datumet för lastningen.
3. Varje transportföretag skall se till att det dokument som avses i punkt 1 innehåller minst alla de uppgifter som anges i punkt 2.
4. Transportföretaget skall undantas från sin skyldighet enligt punkt 1 om något av följande villkor är uppfyllt:
a) Dokumentet enligt punkt 1 ersätts med en kopia av en av de deklarationer som avses i artiklarna 8 eller 10 i fråga om de transporterade mängderna.
b) Dokumentet enligt punkt 1 ersätts med en kopia av dokumentet T 2 M, som anger de transporterade mängdernas ursprung.
5. En medlemsstats behöriga myndigheter kan bevilja undantag från skyldigheten enligt punkt 1 om fiskmängderna transporteras innanför hamnområdet eller högst 20 km från landningsplatsen.
6. Varje medlemsstat skall göra stickprovskontroller på sitt territorium för att undersöka om förpliktelserna enligt denna artikel uppfylls.
7. Medlemsstaterna skall samordna sin kontrollverksamhet för att kontrollen skall bli så effektiv och ekonomisk som möjligt. Medlemsstaterna skall därför särskilt övervaka de varutransporter som tilldragit sig deras uppmärksamhet och som de misstänker strider mot gemenskapens föreskrifter.
Artikel 14
1. Medlemsstaterna skall se till att alla landningar som äger rum i en medlemsstat enligt artiklarna 8, 9 och 10 registreras. De kan därför kräva att den första saluföringen sker genom offentlig auktion.
2. Om den första saluföringen av landade fångster inte sker genom offentlig auktion i enlighet med bestämmelserna i artikel 9.2, skall medlemsstaterna se till att auktionsinrättningarna eller de andra organ som de bemyndigat erhåller information om ifrågavarande mängder.
3. Undantag kan göras från skyldigheten att behandla uppgifter om vilka mängder som landats av vissa kategorier av fartyg som omfattas av undantagen i artiklarna 7 och 8 eller vilka mängder som landats i hamnar som inte har en tillräckligt utvecklad administrativ struktur för att kunna registrera landningarna om en medlemsstat lämnar in en begäran om detta till kommissionen inom tolv månader efter det att denna förordning trätt i kraft. Ett sådant undantag kan beviljas om registreringen av dessa data skulle vara en oproportionerligt stor belastning för de nationella myndigheterna i förhållande till de totala mängder som landats, och om de landade arterna säljs lokalt. Varje medlemsstat skall upprätta en förteckning över de hamnar och fartyg som uppfyller kraven för ett sådant undantag och sända denna till kommissionen.
4. De medlemsstater som omfattas av undantaget i punkt 3 skall utarbeta en provtagningsplan för att bedöma storleken på de fångster som landats i de olika berörda hamnarna. Denna plan skall ha godkänts av kommissionen innan något undantag får göras. Medlemsstaten skall regelbundet sända resultaten av dessa bedömningar till kommissionen.
Artikel 15
1. Före den 15 i varje månad skall varje medlemsstat genom dataöverföring anmäla till kommissionen vilka mängder ur varje bestånd eller grupp av bestånd som omfattas av en TAC eller kvot som landats under föregående månad, samt ge kommissionen alla de upplysningar som erhållits enligt artiklarna 11 och 12.
En sådan anmälan till kommissionen skall innehålla uppgift om fångstplatsen enligt artiklarna 6 och 8 samt om de berörda fiskefartygens nationalitet.
Varje medlemsstat skall ge kommissionen en prognos över kvotutnyttjandet med angivande av det datum när kvoten beräknas vara uttömd för de arter som tagits från fiskefartyg som för denna medlemsstats flagg eller är registrerade där, när det bedöms att fångsterna av dessa arter uppgår till 70 % av den kvot, tilldelning eller andel som den staten förfogar över.
När fångsterna ur bestånd eller grupper av bestånd som omfattas av TAC:er eller kvoter riskerar att nå nivån för gällande TAC:er eller kvoter skall medlemsstaterna på kommissionens begäran lämna mer ingående upplysningar eller lämna sådana oftare än vad som krävs enligt denna punkt.
2. Kommissionen skall hålla de upplysningar som den tagit emot enligt denna artikel tillgängliga för medlemsstaterna genom dataöverföring.
3. Om kommissionen finner att en medlemsstat inte hållit den frist för överföring av uppgifter om månatliga fångster som fastställs i punkt 1 kan den fastställa ett datum när fångsterna ur ett bestånd eller en grupp av bestånd, som omfattas av en kvot eller någon annan form av mängdbegränsning, och som tas från fiskefartyg som för denna medlemsstats flagg eller är registrerade i denna medlemsstat, skall anses utgöra 70 % av den kvot, tilldelning eller andel som denna medlemsstat förfogar över, samt ett datum för när kvoten, tilldelningen eller andelen skall anses vara uttömd.
4. Varje medlemsstat skall före utgången av den första månaden i varje kvartal genom dataöverföring anmäla till kommissionen vilka mängder som landats under föregående kvartal av andra bestånd än de som avses i punkt 1.
Artikel 16
1. Utan att det påverkar tillämpningen av artikel 15 skall medlemsstaterna på den berörda medlemsstatens begäran lämna upplysning om de landningar, utbjudningar till försäljning eller omlastningar av fiskeprodukter som äger rum i deras hamnar eller i de farvatten som lyder under deras jurisdiktion från sådana fiskefartyg som för denna medlemsstats flagg eller är registrerade i denna, och som omfattar fisk ur ett bestånd eller en grupp av bestånd från en kvot som tilldelats denna medlemsstat.
Denna information skall bestå av ifrågavarande fartygs namn och distriktsbeteckning, vilka fiskmängder per bestånd eller grupp av bestånd som detta fartyg landat, bjudit ut till försäljning eller lastat om samt dagen och platsen för landningen, den första utbjudningen till försäljning eller omlastningen. Denna information skall överlämnas inom fyra arbetsdagar räknat från medlemsstatens förfrågan, eller inom en längre tidsfrist, som denna medlemsstat eller landningsmedlemsstaten kan fastställa.
2. På kommissionens anmodan skall den medlemsstat där landningen äger rum, fångsten för första gången bjuds ut till försäljning eller där omlastningen sker sända in dessa upplysningar till kommissionen, samtidigt som den sänder dem till den medlemsstat där fartyget är registrerat.
Artikel 17
1. Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa att fångsterna av sådana arter som deras fartyg tar såväl i farvatten som lyder under ett tredje lands överhöghet eller jurisdiktion som på internationellt vatten utanför zongränserna övervakas, och att omlastningar och landningar av sådana fångster granskas och registreras.
2. Kontrollåtgärderna skall säkerställa att ägarna eller befälhavarna uppfyller följande förpliktelser:
- Fiskefartygen skall ha en loggbok ombord, i vilken befälhavarna registrerar sina fångster.
- Under landning i gemenskapens hamnar skall en landningsdeklaration lämnas in till myndigheterna i den medlemsstat där landningen äger rum.
- Flaggmedlemsstaten skall närmare underrättas om alla omlastningar av fisk till fiskefartyg från tredje land och om landningar som sker direkt i tredje land.
3. Bestämmelserna i punkterna 1 och 2 skall tillämpas utan att det påverkar tillämpningen av bestämmelserna i de fiskeavtal som slutits mellan gemenskapen och tredje land, samt de internationella konventioner som gemenskapen anslutit sig till.
Artikel 18
1. Varje medlemsstat skall före utgången av den första månaden i varje kvartal på elektronisk väg anmäla till kommissionen vilka mängder som tagits i de farvatten som anges i artikel 17 och som landats under föregående kvartal, samt lämna kommissionen alla de upplysningar som erhållits i enlighet med artikel 17.2.
2. För sådana fångster som tas i ett tredje lands farvatten skall den information som lämnas i enlighet med punkt 1 anges per tredje land och bestånd med hänvisning till det minsta statistiska område som fastställts för ifrågavarande fiskeverksamhet.
Fångster som tas på internationellt vatten utanför zongränserna skall anmälas med hänvisning till det minsta statistiska område som fastställs i den internationella konventionen om fångstplats för varje art eller grupp av arter för alla bestånd som ingår i ifrågavarande fiskeverksamhet.
3. Före den 1 oktober varje år skall kommissionen se till att medlemsstaterna får tillgång till den information som den erhållit enligt denna artikel.
Artikel 19
1. För att säkerställa att de förpliktelser som fastställs i artiklarna 3, 6, 8, 9, 10, 14 och 17 uppfylls skall varje medlemsstat införa ett system för giltighetskontroll, som skall omfatta dubbelkontroller och granskning av de uppgifter som kommit in till följd av dessa förpliktelser.
2. För att underlätta denna granskning skall varje medlemsstat upprätta en elektronisk databas, där sådana data som avses i punkt 1 registreras.
Medlemsstaterna får upprätta decentraliserade databaser på villkor att dessa databaser och de metoder som används för insamling och registrering av data är standardiserade, så att de är kompatibla med varandra på en medlemsstats hela territorium.
3. Om en medlemsstat inte omedelbart kan uppfylla kraven i punkt 2 med avseende på delar av eller hela sitt fiske kan kommissionen på denna medlemsstats begäran besluta att i enlighet med förfarandet i artikel 36 bevilja den en övergångsperiod på högst tre år räknat från den dag denna förordning träder i kraft.
4. En medlemsstat som beviljats sådana undantag skall under en tid av tre år föra ett icke elektroniskt register över de uppgifter som avses i punkt 1 och upprätta en provtagningsplan, som skall godkännas av kommissionen, så att en kontroll av uppgifternas riktighet skall kunna göras på platsen. Kommissionen skall på eget initiativ kunna företa granskningar på platsen för att kunna utvärdera provtagningsplanens effektivitet.
5. Inom tolv månader efter det att denna förordning trätt i kraft skall varje medlemsstat lämna in en rapport till kommissionen, i vilken det beskrivs hur uppgifterna samlas in och kontrolleras och hur tillförlitliga de är. Kommissionen skall i samarbete med medlemsstaterna göra en sammanfattning av rapporterna, som den skall delge medlemsstaterna.
6. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 36.
Artikel 20
1. Alla fångster som bevaras ombord på ett fiskefartyg inom gemenskapen skall vara i överensstämmelse med den artsammansättning som fastställs för nätredskapen ombord på fartyget i fråga i rådets förordning (EEG) nr 3094/86 av den 7 oktober 1986 om vissa tekniska åtgärder för bevarande av fiskeresurserna().
Nätredskap som finns ombord men inte används skall stuvas undan så att de inte kan användas utan vidare i enlighet med följande bestämmelser:
a) Nätredskapen, vikterna och liknande utrustning skall lösgöras från trålborden, sveplinorna, trålvarpen och repen.
b) Nätredskapen som finns på däck eller ovanför däck skall vara säkert fastgjorda vid någon del av överbyggnaden.
2. Om fångsterna ombord på något av gemenskapens fiskefartyg tagits med nät med olika minsta maskstorlek under samma resa skall artsammansättningen beräknas för varje del av den fångst som tagits under olika förhållanden.
Varje ändring av en tidigare använd maskstorlek, liksom av fångstsammansättningen ombord vid tidpunkten för denna ändring skall därför skrivas in i loggboken och landningsdeklarationen. I speciella fall skall närmare bestämmelser om hur en stuvningsplan över bearbetade produkter för varje art skall utarbetas och hållas uppdaterad antas i enlighet med det förfarande som fastställs i artikel 36, med angivande av produkternas placering under däck.
3. Trots bestämmelserna i punkterna 1 och 2 kan rådet på grundval av en rapport utarbetad av kommissionen på dennas förslag med kvalificerad majoritet besluta att
a) inget av gemenskapens fiskefartyg som deltar i speciella typer av fiske får medföra nät med olika minsta maskstorlek under samma resa,
b) speciella regler skall gälla för användningen av nät med olika maskstorlek vid speciella typer av fiske.
Artikel 21
1. Alla fångster ur ett kvoterat bestånd eller en kvoterad grupp av bestånd, som tas av gemenskapens fiskefartyg skall skrivas av från den kvot som tilldelats flaggmedlemsstaten för gällande bestånd eller grupp av bestånd, oberoende av landningsplatsen.
2. Varje medlemsstat skall fastställa ett datum när fångsterna ur ett kvoterat bestånd eller en kvoterad grupp av bestånd, som tagits av sådana fiskefartyg som för dess flagg eller är registrerade i den staten skall anses ha förbrukat den kvot som den tilldelats för detta bestånd eller denna grupp av bestånd. Från detta datum skall den tills vidare förbjuda nämnda fartyg att fiska ur detta bestånd eller denna grupp av bestånd och att bevara ombord, omlasta och landa fisk som fångats efter detta datum, och fastställa ett datum fram till vilket det är tillåtet att lasta om och landa fångster eller lämna in de senaste fångstdeklarationerna. Denna åtgärd skall omgående anmälas till kommissionen, som sedan skall informera de övriga medlemsstaterna om den.
3. Efter en anmälan i enlighet med punkt 2, eller på eget initiativ, skall kommissionen på grundval av tillgänglig information fastställa ett datum för när de fångster ur ett bestånd eller en grupp av bestånd som omfattas av en TAC, kvot eller någon annan form av mängdbegränsning, som de fiskefartyg tagit som för en medlemsstats flagg eller är registrerade i en medlemsstat, skall anses ha förbrukat den kvot, tilldelning eller andel som står till denna medlemsstats eller, eventuellt, gemenskapens förfogande.
I samband med bedömningen av den situation som avses i första stycket skall kommissionen informera de berörda medlemsstaterna om sannolikheten av ett fiskestopp till följd av att en TAC är förbrukad.
Gemenskapens fiskefartyg skall upphöra med att fiska en art ur ett bestånd eller en grupp av bestånd som omfattas av en kvot eller TAC den dag när den kvot som tilldelats denna stat för beståndet eller gruppen av bestånd ifråga anses vara förbrukad, eller den dag när TAC:en för de arter som utgör detta bestånd eller denna grupp av bestånd anses vara förbrukad; dessa fartyg skall också upphöra med att bevara ombord, lasta om, landa eller låta lasta om eller landa fångster ur de bestånd eller grupper av bestånd som tagits efter denna dag.
4. När kommissionen i enlighet med punkt 3 första stycket har stoppat fiskeverksamheten på grund av att den TAC, kvot, tilldelning eller andel som står till gemenskapens förfogande antas vara förbrukad, och det visar sig att en medlemsstat i själva verket inte har förbrukat den kvot, tilldelning eller andel som den förfogar över av ifrågavarande bestånd eller grupp av bestånd, skall följande bestämmelser tillämpas.
Om den skada som en medlemsstat lidit genom att fisket förbjudits innan dess kvot förbrukats inte avhjälpts i enlighet med artikel 9.2 i förordning nr 3760/92, skall åtgärder beslutas på det sätt som anges i artikel 36 i syfte att på ett lämpligt sätt reparera den skada som förorsakats. Dessa åtgärder kan innebära att det görs avdrag för den medlemsstat som överskridit sin kvot, tilldelning eller andel, och att de mängder som dras av på ett lämpligt sätt delas ut till de medlemsstater vars fiske stoppats innan deras kvot förbrukats. Dessa avdrag och efterföljande tilldelningar skall göras med hänsyn till i första hand de arter och zoner för vilka kvoterna, tilldelningarna eller de årliga andelarna fastställts. Dessa avdrag eller tilldelningar kan göras under det år skadan uppstår eller under något av de följande åren.
Tillämpningsföreskrifter för denna punkt skall fastställas i enlighet med det förfarande som anges i artikel 36, särskilt beträffande bestämningen av ifrågavarande mängder.
Artikel 22
1. Om en medlemsstats behöriga myndigheter finner att ett av gemenskapens fiskefartyg allvarligt eller upprepade gånger brutit mot denna förordning kan flaggmedlemsstaten underkasta fartyget ytterligare kontroll.
Flaggmedlemsstaten skall meddela kommissionen och de övriga medlemsstaterna namnet och distriktsbeckningen på det fartyg som underkastats sådan ytterligare kontroll.
Artikel 23
1. Om kommissionen konstaterat att en medlemsstat överskridit sin kvot, tilldelning eller andel av ett bestånd eller en grupp av bestånd skall kommissionen göra avdrag från den årliga kvot, tilldelning eller andel som den medlemsstaten förfogar över. Dessa avdrag skall fastställas i enlighet med förfarandet i artikel 36.
2. Rådet skall på kommissionens förslag med kvalificerad majoritet anta avdragsbestämmelser i enlighet med de mål och förvaltningsstrategier som anges i artikel 8 i förordning (EEG) nr 3760/92, och skall då i första hand ta hänsyn till följande parametrar:
- Överfiskets omfång.
- Eventuella fall av överfiske av samma bestånd under de föregående åren.
- De berörda beståndens biologiska tillstånd.
Artikel 24
För att säkerställa att de mål och strategier som fastläggs av rådet i enlighet med artikel 11 i förordning (EEG) nr 3760/92 följs, särskilt mängdmålen avseende fiskekapaciteten hos gemenskapens fiskeflotta och anpassningen av fiskeflottans verksamhet, skall varje medlemsstat på sitt territorium och i de farvatten som lyder under dess överhöghet eller jurisdiktion göra regelbundna kontroller hos alla dem som berörs av genomförandet av ovan nämnda mål.
Artikel 25
1. Varje medlemsstat skall anta bestämmelser för att kontrollera att de mål som avses i artikel 24 uppfylls. Den skall därför företa tekniska kontroller, särskilt på följande områden:
a) Omstrukturering, förnyelse och modernisering av fiskeflottan.
b) Anpassning av fiskekapaciteten genom temporärt eller definitivt stopp.
c) Begränsning av vissa fiskefartygs verksamhet.
d) Begränsning av fiskeredskapens utformning och antal, samt deras användningssätt.
e) Utveckling av vattenbruket och kustområdena.
2. Utan att det påverkar tillämpningen av artikel 169 i fördraget kan kommissionen, om den finner att en medlemsstat inte följt bestämmelserna i punkt 1, lägga fram förslag till rådet om att anta lämpliga allmänna åtgärder. Rådet skall fatta beslut med kvalificerad majoritet.
Artikel 26
1. Tillämpningsföreskrifter för artikel 25 kan antas i enlighet med det förfarande som anges i artikel 36, särskilt med avseende på kontrollen av
a) fiskefartygens maskinstyrka,
b) fiskefartygens registertonnage,
c) fiskefartygens stillaliggandeperiod,
d) fiskeredskapens karakteristika och deras antal per fiskefartyg.
2. Medlemsstaterna skall omgående meddela kommissionen vilka kontrollmetoder som används samt namn och adress till de organ som svarar för kontrollen.
Artikel 27
1. För att underlätta den kontroll som avses i artikel 25 skall medlemsstaterna införa ett system för giltighetskontroll, som särskilt skall omfatta en korsvis kontroll av uppgifterna om fiskeflottans kapacitet och verksamhet i bl.a.
- den loggbok som avses i artikel 6,
- den landningsdeklaration som avses i artikel 8,
- gemenskapens förteckning över fiskefartyg, som avses i kommissionens förordning (EEG) nr 163/89().
2. För detta ändamål skall medlemsstaterna upprätta databaser eller bygga ut redan existerande databaser med relevant information om fiskeflottans kapacitet och verksamhet.
3. De åtgärder som avses i artikel 19.3, 19.4 och 19.5 skall tillämpas.
4. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som anges i artikel 36.
Artikel 28
1. För att säkerställa att de tekniska aspekterna av de föreskrifter om åtgärder som fastställs i förordning (EEG) nr 3759/92 av den 17 december 1992 om den gemensamma organisationen av marknaden för fiske- och vattenbruksprodukter() följs skall varje medlemsstat på sitt territorium organisera regelbundna kontroller av alla dem som berörs av tillämpningen av dessa åtgärder.
2. Dessa kontroller skall gälla de tekniska aspekterna av tillämpningen av
a) handelsstandarder, särskilt minsta storlekar,
b) prisreglering, särskilt vid
- återtagande av produkter från marknaden för andra ändamål än mänsklig konsumtion,
- lagring och/eller bearbetning av produkter som återtagits från marknaden.
Medlemsstaterna skall göra jämförelser mellan dokumenten avseende den första saluföringen av de mängder som anges i artikel 9 och de landade mängder som dokumenten anger, särskilt med avseende på deras vikt.
3. Medlemsstaterna skall ge kommissionen upplysningar om utförda kontroller, behöriga kontrollmyndigheter, konstaterade överträdelser och vilka åtgärder som dessa föranlett.
Kommissionen och medlemsstaternas behöriga myndigheter, samt tjänstemän och andra ombud, får inte sprida sådan information som samlas in genom tillämpningen av denna artikel som omfattas av tystnadsplikt.
4. Denna artikel skall inte inverka på de nationella bestämmelserna om sekretess vid rättsligt förfarande.
Artikel 29
1. Kommissionen skall kontrollera att medlemsstaterna tillämpar denna förordning genom att granska dokument och göra besök på platsen. Om kommissionen finner det lämpligt kan den företa granskningar utan förvarning.
Inför besök på platsen skall kommissionen utfärda skriftliga instruktioner åt sina inspektörer med angivande av deras befogenhet och ändamålet med deras uppdrag.
2. Närhelst kommissionen anser det nödvändigt kan dess inspektörer närvara vid de nationella tillsynsmyndigheternas kontroller och inspektioner. Inom ramen för detta uppdrag skall kommissionen upprätta lämpliga kontakter med medlemsstaterna för att om möjligt utarbeta ett inspektionsprogram som kan godtas av båda parter.
a) Medlemsstaterna skall samarbeta med kommissionen för att underlätta för denna att genomföra sina uppdrag. De skall särskilt vidta alla nödvändiga åtgärder för att inspektionerna inte skall offentliggöras, vilket skulle kunna störa genomförandet av inspektionen och kontrollen.
Om kommissionen eller dess ombud stöter på svårigheter under genomförandet av sina uppdrag, skall medlemsstaterna ställa medel till kommissionens förfogande så att den kan slutföra sin uppgift, och de skall ge inspektörerna möjlighet att utvärdera kontrollerna ifråga.
b) Om förhållandena på platsen gör det omöjligt att genomföra den inspektion och kontroll som planerats i det ursprungliga inspektionsprogrammet skall kommissionens inspektörer i samarbete med den behöriga tillsynsmyndigheten, och med dess samtycke, ändra den ursprungligen planerade inspektionen och kontrollen.
c) Vid inspektion till havs eller från luften skall medlemsstaternas myndigheter i de fall de nationella behöriga organen skall tillvarata andra viktiga uppgifter, särskilt i samband med försvaret eller säkerheten till sjöss, ha rätt att skjuta upp eller omdirigera de inspektioner som kommissionen planerat att närvara vid. I sådana fall skall medlemsstaten samarbeta med kommissionen för att vidta alternativa åtgärder.
Vid inspektioner till havs eller från luften är fartygets eller flygplanets befälhavare ensam ansvarig för inspektionen med hänsyn till dennes myndigheters skyldighet att tillämpa denna förordning. De av kommissionens inspektörer som deltar i inspektionen skall följa de regler och den praxis som befälhavaren fastställer.
3. Kommissionen kan vid behov, särskilt om gemenskapens inspektörer i enlighet med punkt 2 avslöjat att oegentligheter kan ha begåtts vid tillämpningen av denna förordning, anmoda medlemsstaterna att lämna närmare uppgifter om vilket inspektions- och kontrollprogram som de behöriga nationella myndigheterna planerat eller fastställt för en viss period och fiskeverksamhet samt vissa områden. Efter mottagandet av denna information skall kommissionens inspektörer, om denna anser det nödvändigt, göra egna inspektioner för att granska hur en medlemsstats behöriga myndigheter genomfört detta program.
När gemenskapens inspektörer granskar tillämpningen av detta program är medlemsstatens ombud alltid ansvariga för dess genomförande. Gemenskapens inspektörer kan inte på eget initiativ använda sig av de inspektionsbefogenheter som anförtrotts de nationella ombuden. Dessa inspektörer har bara tillgång till fartyg eller lokaler om de ledsagas av en medlemsstats ombud.
Efter denna kontroll skall kommissionen sända en utvärderingsrapport om programmet till den berörda medlemsstaten och eventuellt rekommendera den att vidta åtgärder för att förbättra genomförandet av kontrollerna.
4. Vid inspektioner från luften, till havs eller till lands, får de behöriga inspektörerna inte företa någon kontroll av fysiska personer.
5. Inom ramen för de besök som nämns i punkterna 2 och 3 skall kommissionens behöriga inspektörer i de ansvariga organens närvaro på platsen få tillträde till hela eller delar av informationen i de specificerade databaserna och få granska alla de dokument som är relevanta för tillämpningen av denna förordning.
Om de nationella bestämmelserna föreskriver sekretess under förundersökningen får denna information inte lämnas ut utan tillstånd från den behöriga juridiska instansen.
Artikel 30
1. Medlemsstaterna skall till kommissionen på dennas begäran överlämna all information om tillämpningen av denna förordning. Om kommissionen begär information skall den ange en rimlig tid inom vilken denna skall lämnas.
2. Om kommissionen finner att oegentligheter begåtts vid tillämpningen av denna förordning eller att de existerande kontrollmetoderna och kontrollbestämmelserna inte är effektiva, skall den meddela den eller de berörda medlemsstaterna, som då skall sätta igång en administrativ undersökning, i vilken tjänstemän från kommissionen kan delta.
Den eller de berörda medlemsstaterna skall informera kommissionen om undersökningens förlopp och resultat och lämna kommissionen en kopia av undersökningsrapporten och de centrala bevismaterial som legat till grund för utarbetandet av rapporten.
För att kunna delta i de inspektioner som avses i denna punkt skall kommissionens tjänstemän visa fram en skriftlig fullmakt, av vilken deras identitet och tjänstebeteckning framgår.
3. När kommissionens inspektörer deltar i en undersökning skall denna alltid ledas av medlemsstatens tjänstemän. Kommissionens tjänstemän får inte på eget initiativ använda sig av de inspektionsbefogenheter som tilldelats de nationella inspektörerna. Men de skall ha tillgång till samma lokaler och handlingar som dessa inspektörer.
Om det enligt nationell lagstiftning är förbehållet vissa i lagen angivna tjänstemän att utföra vissa handlingar på det straffrättsliga området skall kommissionens tjänstemän avhålla sig från att medverka i dessa handlingar. De skall särskilt avhålla sig från att delta i husrannsakningar och formella förhör av personer enligt nationell straffrätt. De skall dock ha tillträde till den information som fås på detta sätt.
4. Denna artikel påverkar inte de nationella bestämmelserna om sekretess vid rättsligt förfarande.
Artikel 31
1. Medlemsstaterna skall se till att lämpliga åtgärder vidtas mot ansvariga fysiska eller juridiska personer, även sådana förvaltnings- eller straffrättsliga åtgärder som överensstämmer med nationell lagstiftning, när det, särskilt efter en kontroll eller inspektion som utförts enligt denna förordning, står klart att den gemensamma fiskeripolitikens bestämmelser inte följts.
2. De rättsliga åtgärder som vidtas med stöd av punkt 1 skall vara av sådan art att de i enlighet med tillämpliga bestämmelser i den nationella lagstiftningen effektivt berövar de ansvariga det ekonomiska utbytet av överträdelsen eller framkallar effekter som står i proportion till överträdelsens allvar, i syfte att avskräcka från ytterligare överträdelser av samma slag.
3. Påföljderna av det rättegångsförfarande som avses i punkt 2 kan beroende på brottets allvar omfatta
- böter,
- beslag av förbjudna fiskeredskap och fångster,
- beslag av fartyget,
- tillfällig indragning av licensen,
- återkallande av licensen.
4. Bestämmelserna i denna artikel får inte hindra landnings- eller omlastningsmedlemsstaten från att överlåta den rättsliga uppföljningen av en överträdelse på de behöriga myndigheterna i registreringsmedlemsstaten, om denna samtycker till det, förutsatt att en sådan överlåtelse skapar bättre förutsättningar för att uppnå det resultat som avses i punkt 2. Landnings- eller omlastningsmedlemsstaten skall anmäla varje sådan överlåtelse till kommissionen.
Artikel 32
1. Om de behöriga myndigheterna i landnings- eller omlastningsmedlemsstaten konstaterar att en överträdelse skett mot denna förordning skall de vidta lämpliga åtgärder i enlighet med artikel 31 mot ifrågavarande fartygs befälhavare eller mot någon annan person som är ansvarig för överträdelsen.
2. Om landnings- eller omlastningsmedlemsstaten inte är densamma som flaggmedlemsstaten, och de behöriga myndigheterna inte i enlighet med sin nationella lagstiftning vidtar lämpliga åtgärder, inbegripet förvaltnings- eller straffrättsliga åtgärder mot de ansvariga fysiska eller juridiska personerna, eller inte överlåter den rättsliga uppföljningen i enlighet med artikel 31.4, får den mängd fisk som olovligen landats eller lastats om skrivas av från den medlemsstatens kvot.
Vilken fiskmängd som skall skrivas av från den medlemsstatens kvot skall fastställas på det sätt som anges i artikel 36, när kommissionen har hört de två berörda medlemsstaterna.
Om landnings- eller omlastningsmedlemsstaten inte längre har motsvarande kvot till sitt förfogande skall artikel 21.4 också tillämpas, och de olovligen landade eller omlastade fiskmängderna anses motsvara omfånget av den skada som registreringsmedlemsstaten lidit på det sätt som anges i den artikeln.
Artikel 33
1. Medlemsstaternas behöriga myndigheter skall omgående i enlighet med den nationella lagstiftningens förfarande till flagg- eller registreringsmedlemsstaten anmäla alla överträdelser av de gemenskapsbestämmelser som avses i artikel 1, med angivande av det berörda fartygets namn och distriktsbeteckning, befälhavarens och ägarens namn, omständigheterna kring överträdelsen och de förvaltnings- eller straffrättsliga påföljderna, eller andra åtgärder som vidtagits samt alla slutgiltiga avgöranden i samband med sådana överträdelser. I speciella fall skall medlemsstaterna efter anmodan överlämna denna information till kommissionen.
2. Efter en överlåtelse av den rättsliga uppföljningen i enlighet med artikel 31.4 skall flagg- eller registreringsmedlemsstaten vidta varje sådan lämplig åtgärd som avses i artikel 31.
3. Flagg- eller registreringsmedlemsstaten skall omgående anmäla till kommissionen vilka åtgärder som vidtagits i enlighet med punkt 2, samt det berörda fartygets namn och distriktsbeteckning.
Artikel 34
1. Medlemsstaterna skall till kommissionen anmäla vilka lagar och andra författningar de antagit för att förebygga och beivra lagöverträdelser.
De skall varje år anmäla alla ändringar av böternas minimi- och maximibelopp för varje typ av överträdelse, samt alla andra slag av tillämpliga påföljder.
2. Medlemsstaterna skall regelbundet underrätta kommissionen om resultaten av de inspektioner eller kontroller som görs med stöd av denna förordning, särskilt vilken mängd och typ av överträdelse som konstaterats och vilka åtgärder som vidtagits. Medlemsstaterna skall på kommissionens anmodan till denna anmäla vilka bötesbelopp som tillämpats i de konkreta fallen av överträdelse.
3. Kommissionen skall förse medlemsstaterna med ett sammandrag av de upplysningar som den erhållit i enlighet med punkterna 1 och 2.
Artikel 35
Medlemsstaterna skall före den 1 juni varje år överlämna en rapport till kommissionen om tillämpningen av denna förordning under föregående kalenderår; denna skall innehålla en utvärdering av de tekniska och mänskliga insatserna och ange vilka åtgärder som skulle kunna bidra till att mildra de brister som eventuellt kunnat konstateras. På grundval av medlemsstaternas rapporter och de egna observationerna skall kommissionen sammanställa en årlig rapport och till varje medlemsstat överlämna de delar av rapporten som berör denna. Efter att ha tagit vederbörlig hänsyn till medlemsstaternas svar skall kommissionen offentliggöra hela rapporten med medlemsstaternas svar och eventuella förslag till åtgärder i syfte att avhjälpa de konstaterade bristerna.
Artikel 36
När förfarandet i denna artikel skall tillämpas, skall ordföranden hänskjuta ärendet till Förvaltningskommittén för fiske och vattenbruk som inrättats genom förordning (EEG) nr 3760/92, nedan kallad "kommittén", antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen, varvid medlemsstaternas röster skall vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
Kommissionen skall besluta med omedelbar verkan. Om beslutet inte är förenligt med kommitténs yttrande skall kommissionen emellertid genast underrätta rådet. I sådana fall får kommissionen uppskjuta verkställandet av de beslutade åtgärderna under en tid som inte överstiger en månad från dagen då rådet underrättats.
Rådet får fatta ett annat beslut med kvalificerad majoritet inom den tid som anges i föregående stycke.
Artikel 37
1. Medlemsstaterna och kommissionen skall vidta alla nödvändiga åtgärder för att säkerställa att de uppgifter som tas emot inom ramen för denna förordning behandlas konfidentiellt.
2. Namnen på de fysiska eller juridiska personerna skall bara meddelas kommissionen eller en annan medlemsstat i de fall det uttryckligen anges i denna förordning, eller om det är nödvändigt för att förebygga eller beivra överträdelser eller granska uppenbara överträdelser.
Uppgifterna i punkt 1 skall bara föras vidare om de är så införlivade med andra uppgifter att de berörda fysiska eller juridiska personerna inte direkt eller indirekt kan identifieras.
3. Uppgifterna som utväxlas mellan medlemsstaterna och kommissionen får bara lämnas vidare till de personer i medlemsstaternas och gemenskapens institutioner vars uppgifter kräver att de har tillgång till dem; om de lämnas till andra personer skall de medlemsstater som lämnat uppgifterna uttryckligen ha givit sitt samtycke till det.
4. De uppgifter som lämnas eller tas emot i en eller annan form med stöd av denna förordning omfattas av tystnadsplikt och skall åtnjuta samma skydd som liknande uppgifter åtnjuter, såväl genom den nationella lagstiftningen i de medlemsstater som tar emot uppgifterna som genom motsvarande bestämmelser som är tillämpliga på gemenskapens institutioner.
5. Uppgifterna i punkt 1 får inte användas för något annat ändamål än det som anges i denna förordning, om inte de myndigheter som lämnar dem uttryckligen samtycker till det, och gällande bestämmelser i den medlemsstat vars myndighet tar emot uppgifterna inte förbjuder en sådan användning eller utlämning av uppgifter.
6. Bestämmelserna i punkt 1 5 får inte tolkas som ett hinder mot att de uppgifter som erhålls genom tillämpningen av denna förordning används inom ramen för sådana rättsliga åtgärder som vidtas senare på grund av att gemenskapens fiskelagstiftning inte följts. De behöriga myndigheterna i den medlemsstat som lämnar uppgifterna skall informeras om alla de fall i vilka uppgifterna används i detta syfte.
Denna artikel påverkar inte de skyldigheter som följer av internationella konventioner om ömsesidigt bistånd i straffrättsliga frågor.
7. Varje gång en medlemsstat meddelar kommissionen att den efter en slutförd undersökning funnit att en fysisk eller juridisk person, vars namn meddelats den i kraft av bestämmelserna i denna förordning, inte varit inblandad i en överträdelse, skall kommissionen omedelbart underrätta alla dem som den lämnat ut den berörda personens namn till om utgången av undersökningen eller de rättsliga åtgärderna. Personen ifråga skall inte längre behandlas som om han eller hon vore inblandad i de oegentligheter som det första meddelandet innehöll uppgift om. De uppgifter som bevaras på ett sådant sätt att den berörda personen kan identifieras skall omgående förstöras.
8. Bestämmelserna i punkt 1 5 får inte tolkas som ett hinder mot att allmänna upplysningar eller undersökningar offentliggörs, som inte nämner enskilda fysiska eller juridiska personer.
9. Uppgifterna i denna förordning skall bevaras på ett sådant sätt att de berörda personerna bara kan identifieras under den tid som behövs för ändamålet ifråga.
10. De upplysningar som tas emot inom ramen för denna förordning skall på begäran ställas till de berörda fysiska eller juridiska personernas förfogande.
Artikel 38
Denna förordning skall gälla utan att det påverkar tillämpningen av eventuella nationella kontrollåtgärder som sträcker sig utanför minimikraven, under förutsättning att de är förenliga med gemenskapsrätten och den gemensamma fiskeripolitiken.
De nationella åtgärder som avses i första stycket skall anmälas till kommissionen i enlighet med artikel 2.2 i rådets förordning (EEG) nr 101/76 av den 19 januari 1976 om en gemensam strukturpolitik för fiskerisektorn().
Artikel 39
1. Förordning (EEG) nr 2241/87 skall upphöra att gälla den 1 januari 1994 med undantag för artikel 5, som skall fortsätta att gälla till dess förordningarna om utarbetande av de förteckningar som avses i artikel 6.2 i denna förordning har trätt i kraft.
2. Hänvisningar till den i punkt 1 upphävda förordningen skall anses som hänvisningar till denna förordning.
Artikel 40
Denna förordning träder i kraft den 1 januari 1994.
Medlemsstaterna skall fram till den 1 januari 1996 undantas från skyldigheten att tillämpa bestämmelserna i artiklarna 9, 15 och 18 i fråga om dataöverföring av avräkningsnotor och registrering av landningar.
Medlemsstaterna skall fram till den 1 januari 1999 undantas från skyldigheten att tillämpa bestämmelserna i artiklarna 6, 8 och 19 i fråga om fiske i Medelhavet.
KOMMISSIONENS FÖRORDNING (EEG) nr 3063/93 av den 5 november 1993 om tillämpningsföreskrifter för rådets förordning (EEG) nr 2019/93 angående stödordningen för produktion av kvalitetshonung
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2019/93 av den 19 juli 1993 om införandet av särskilda bestämmelser för de mindre Egeiska öarna rörande vissa jordbruksprodukter(1) särskilt artikel 12.4 i denna,
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas avseende den gemen-samma jordbrukspolitiken(2), särskilt artikel 6 i denna, och
med beaktande av följande: I artikel 12 i förordning (EEG) nr 2019/93 föreskrivs att stöd skall beviljas de mindre Egeiska öarna för produktion av kvalitetshonung som innehåller en stor andel timjanhonung. Tillämpningsföreskrifter bör antas för förvaltning av ord-ningen och för kontroll av de villkor som rådet har uppställt.
För att uppmuntra honungsproducenter som är medlemmar av organisationer, som överensstämmer med definitionen i rådets förordning (EEG) nr 1360/78 av den 19 juni 1978 om producentgrupper och sammanslutningar av dessa(3), senast ändrad genom förordning (EEG) nr 746/93(4) att förbättra sina saluföringssystem för att tillmötesgå marknadens krav och att främja kvalitetsprodukter, är beviljande av stöd avhängigt att producenterna genomför årliga initiativprog-ram, som godkänns av de myndigheter som Grekland har utsett. För att uppnå målen bör programmet vara inriktat dels på genetiska förbättringar, omställning av bikupor, mekanisering och löpande utbildning för biodlare i ny produktionsteknik, dels på marknadsundersökningar, forskning om nya förpacknings-metoder och säljfrämjande åtgärder.
Tillämpningsföreskrifterna bör också omfatta fastställande av ansökningstid för stödet, vilka uppgifter ansökan minst bör innehålla, den behöriga myndighetens tidsgränser för behandling av ansökan och utbetalning av stöd, samt anmälan till kommissionen om utbetalt stöd. Det bör också fastställas bestämmelser om den kontroll som är nödvändig för att säkerställa att stödordningen tillämpas på ett korrekt sätt, och om vilka åtgärder som skall vidtas vid underlåtenhet att uppfylla bestämmelserna.
Med hänsyn till genomförandet av denna stödordning bör undantag fastställas vad gäller sista ansökningsdag och sista utbetalningsdag för stöd för 1993 års produktion.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommitttén för ägg.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Stödet till produktion av den kvalitetshonung som är specifik för de mindre Egeiska öarna och som innehåller en stor andel timjanhonung, betalas ut till grupper av honungsproducenter som är erkända enligt förordning (EEG) nr 1360/78, och som genomför initiativprogram för att förbättra villkoren för saluföring och marknadsföring av kvalitetshonung.
Fram till slutet av 1994 skall stödet dock även betalas ut till alla biodlare som har minst tio fasta producerande bikupor som är registrerade hos den behöriga myndigheten.
Artikel 2
1. Initiativprogrammet skall ha följande mål:
- Förbättring av saluföringen genom införande av teknik, mekaniserad slungning, rening och filtrering, samt yrkesutbildning.
- Upprätthållande av avkastningen genom att gamla drottningar två gånger om året byts ut mot hybrider som är anpassade till området.
- Främjande av försäljningen av kvalitetshonung genom marknadsundersökningar, utveckling av nya förpackningsmetoder, samt anordnande av och deltagande i varumässor och andra säljfrämjande åtgärder.
2. Sammanslutningarna av honungsproducenter skall förelägga den behöriga myndigheten sina program för god-kännande. Myndigheten skall, senast två månader efter prog-rammets inlämnande, besluta om godkännande eller avslag, efter att i förekommande fall ha anmodat om nödvändiga förändringar.
Artikel 3
1. Stödansökan skall lämnas in till den behöriga myndigheten under den period som dessa fastställer, dock senast den 30 september varje år, när det gäller produktionen för följande år. Vid för sen inlämning sänks stödet med 20 %, utom i fall av force majeure. Om ansökan inlämnas mer än 20 dagar efter den ansökningsperiod som fastställts av den behöriga myndigheten, skall inget stöd betalas ut.
För år 1993 kan emellertid stödansökningar lämnas in senast den 15 december 1993.
2. Stödansökan skall minst innehålla följande uppgifter:
- Sammanslutningens eller biodlarens namn och adress.
- Antal fasta bikupor i produktion och det registrerings-nummer som den behöriga myndigheten tilldelat dem.
- Den mängd honung med stor andel timjanhonung som producerats under den period för vilken det ansöks om stöd.
3. När det totala antalet bikupor för vilka det ansöks om stöd överstiger det högsta tillåtna antalet bikupor enligt artikel 12.3 i förordning (EEG) nr 2019/93, skall den behöriga myndigheten fastställa en schablonmässig koefficient för sänkning av alla stödbelopp.
Artikel 4
Grekland skall betala ut stödet senast den 31 december under den period för vilken stöd beviljas, i proportion till den faktiska graden av genomförande av initiativprogrammet. Stöd skall inte utbetalas om genomförandegraden under-stiger 50 %.
För år 1993 får emellertid stödet betalas ut senast den 28 februari 1994.
Artikel 5
Grekland skall, senast den 31 januari varje år, meddela kommissionen följande:
- Antal producentsammanslutningar och antal individuella biodlare som inkommit med stödansökningar.
- Antal bikupor för vilka producentsammanslutningar och individuella biodlare ansökt om och beviljats stöd.
- Den sänkningskoefficient som eventuellt tillämpas.
- De initiativprogram som blivit godkända.
- Antal oegentligheter som konstaterats och de bikupor som de gäller.
För år 1993 får dessa uppgifter emellertid överlämnas senast den 15 mars 1994.
Artikel 6
1. Grekland skall, genom kontroller på plats, säkerställa att uppgifterna som lämnats i stödansökan är korrekta, samt att villkoren för utbetalning av stöd uppfylls.
- Genomförandet av inititativprogrammet.
Artikel 7
2. Om stöd måste indrivas på grund av oegentligheter som kan tillskrivas sökanden, oavsett om dessa orsakats avsiktligt eller genom grov försumlighet, skall den behöriga myndigheten driva in utbetalda belopp med en höjning på 20 % samt ränta enligt punkt 1. Sökanden skall inte vara berättigad till stöd det följande året.
RÅDETS FÖRORDNING (EEG) nr 3089/93 av den 29 oktober 1993 om ändring av förordning (EEG) nr 2299/89 om en uppförandekod för datoriserade bokningssystem
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 84.2 i detta,
med beaktande av kommissionens förslag (),
med beaktande av Europaparlamentets yttrande (),
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
med beaktande av följande: Förordning (EEG) nr 2299/89 () utgör ett viktigt led i avskaffandet av snedvriden konkurrens mellan lufttrafikföretag och mellan datoriserade bokningssystem, och skyddar därigenom konsumenternas intressen.
Det är nödvändigt att utvidga tillämpningen av förordning (EEG) nr 2299/89 och klargöra dess bestämmelser, och dessa åtgärder bör vidtas på gemenskapsnivå för att säkerställa att förordningens syften uppnås i alla medlemsstater.
Denna förordning inskränker inte tillämpningen av artiklarna 85 och 86 i fördraget.
Enligt kommissionens förordning (EEG) nr 83/91 () är fördragets artikel 85.1 inte tillämplig på överenskommelser om gemensamma inköp, gemensam utveckling och drift av datoriserade bokningssystem.
Icke-regelbunden lufttrafik är av stor betydelse i gemenskapens territorium.
Huvuddelen av dessa resor är paketresor eller kombinerade produkter, där lufttransport bara utgör en del i hela produkten.
I princip konkurrerar "seat-only" eller separata lufttransportprodukter på icke-regelbunden lufttrafik direkt med de lufttransportprodukter som erbjuds på regelbundna flygningar.
Det är önskvärt att likadana produkter behandlas på samma sätt och att säkerställa en rättvis konkurrens mellan de båda typerna av lufttransportprodukter samt en opartisk spridning av information till konsumenten.
Alla frågor som rör användningen av datoriserade bokningssystem för alla typer av lufttransportprodukter bör behandlas i en och samma förordning, som beslutas av rådet.
De konsumenter som söker efter olika produkter bör ges möjlighet att begära textbilder för enbart regelbunden eller icke-regelbunden lufttrafik.
Det bör klargöras att förordning (EEG) nr 2299/89 bör tillämpas på de datoriserade bokningssystem som erbjuds till eller används av alla slutkonsumenter, antingen de är enskilda personer eller företag.
De lufttrafikföretag som använder ett datoriserat bokningssystem i sina egna klart markerade kontor eller diskar bör inte omfattas av bestämmelserna om primär textbild.
Det är lämpligt med en klar åtskillnad mellan ett avtal om deltagande i eller som tillåter användning av ett system och leveransen av den tekniska utrustningen, varvid leveransen omfattas av sedvanlig avtalsrätt vilket ger systemleverantören rätt att kräva att få sina direkta kostnader täckta i de fall då ett avtal om deltagande eller abonnemang sägs upp enligt bestämmelserna i denna förordning.
Om moderföretag vägrar att ge samma information om tidtabeller, biljettpriser och platstillgång till andra system än deras eget och vägrar ta emot bokningar från dessa system kan det allvarligt snedvrida konkurrensen mellan datoriserade bokningssystem.
Att de datoriserade bokningssystemen är konkurrensmässigt neutrala i förhållande till lufttrafikföretag måste säkerställas vad gäller likhet i funktion och datasäkerhet, särskilt genom lika tillträde till funktioner, information/data och gränssnitt samt en klar åtskillnad mellan lufttrafikföretagens egna tjänster och distributionstjänster.
Konkurrensmässig likhet kommer att ökas genom att man säkerställer att de datoriserade bokningssystemen har separat juridisk identitet.
Ett moderföretag kan i konkurrensen mellan lufttrafikföretag få orättvisa fördelar av att det kontrollerar sitt datoriserade bokningssystem. Därför är det nödvändigt med en fullständigt lika behandling av moderföretag respektive deltagande lufttrafikföretag i den utsträckning som ett moderföretag använder de tjänster i dess eget system som omfattas av denna förordning.
I konsumenternas intresse är det önskvärt att en primär textbild ges för varje transaktion som begärs av en konsument.
Det är önskvärt att utförliga upplysningar om avsättning, bokning och försäljning görs tillgängliga för deltagande lufttrafikföretag på ett icke diskriminerande sätt och med samma skyndsamhet. Identifiering av eller personlig information om en passagerare eller ett företag måste förbli konfidentiell. Därför skall en systemleverantör genom tekniska hjälpmedel och lämpliga säkerhetskrav, åtminstone vad gäller mjukvara, säkerställa att otillåtet tillträde till information inte kan äga rum.
Fakturorna bör innehålla tillräckligt med information för att deltagande lufttrafikföretag och abonnenter skall kunna kontrollera sina kostnader. För att underlätta en sådan kontroll bör sådan information göras tillgänglig på magnetiska medier.
I konsumenternas intresse är det önskvärt att klargöra att en flygning eller kombination av flygningar inte skall visas mer än en gång på den primära textbilden, utom i de fall där genom ett konsortium eller någon annan form av uppgörelse varje lufttrafikföretag som bedriver lufttrafik tar på sig separat ansvar för erbjudandet och försäljningen av lufttransportprodukter på de berörda flygningarna.
Systemleverantören skall säkerställa att principerna om teknisk överensstämmelse med bestämmelserna om likhet i funktion och datasäkerhet övervakas av en oberoende kontrollant.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 2299/89 ändras på följande sätt:
Denna förordning skall gälla för datoriserade bokningssystem i den utsträckning som de omfattar lufttransportprodukter som erbjuds eller används inom gemenskapens territorium, oavsett
P systemleverantörens status eller nationalitet,
P varifrån den utnyttjade informationen kommer eller var den centrala databehandlingsanläggningen i fråga är belägen,
P den geografiska belägenheten av de flygplatser mellan vilka lufttransporten äger rum.
Artikel 2
I denna förordning används följande beteckningar med de betydelser som här anges:
a) separat lufttransportprodukt: lufttrafik för befordran av passagerare mellan två flygplatser, inklusive bitjänster och ytterligare förmåner som erbjuds till försäljning och/eller säljs som en integrerad del av lufttransporttjänsten.
b) kombinerad lufttransportprodukt: en på förhand avtalad kombination av en separat lufttransportprodukt med andra tjänster som inte är bitjänster till lufttransport, och som erbjuds till försäljning och/eller säljs till ett totalpris.
c) lufttransportprodukt: både separata lufttransportprodukter och kombinerade lufttransportprodukter.
d) regelbunden lufttrafik: en serie flygningar, där varje flygning uppfyller följande kriterier:
P Den utförs med luftfartyg för befordran av passagerare eller passagerare och gods och/eller post mot vederlag på ett sådant sätt att det på varje flygning finns platser att köpa för enskilda personer (antingen direkt av lufttrafikföretaget eller av dess auktoriserade agenter).
P Den bedrivs så att den betjänar trafiken mellan samma, två eller flera, orter antingen
1. enligt en utgiven tidtabell, eller
2. med flygningar som är så regelbundna eller täta att de utgör en igenkännlig planmässig serie.
e) biljettpris: det pris som skall betalas för separata lufttransportprodukter och villkoren för när detta pris är tillämpligt.
f) datoriserat bokningssystem: ett datoriserat system som innehåller information om bland annat lufttrafikföretags
P tidtabeller,
P platstillgång,
P biljettpriser, och
P tjänster i samband med flygbefordran,
med eller utan möjligheter till
P att reservera platser eller
P att utställa biljetter
av sådan omfattning att några av eller samtliga dessa tjänster ställs till förfogande för abonnenterna.
g) distributionstjänster: tjänster som en systemleverantör ställer till en abonnents eller konsuments förfogande för att förmedla information om lufttrafikföretags tidtabeller, platstillgång, biljettpriser och tjänster i samband med flygbefordran samt för att reservera platser och/eller utställa biljetter och för att tillhandahålla andra tjänster i samband härmed.
h) systemleverantör: varje företag och dess filialer som har ansvaret för driften eller marknadsföringen av ett datoriserat bokningssystem.
i) moderföretag: ett lufttrafikföretag som direkt eller indirekt, ensamt eller tillsammans med andra, äger eller effektivt kontrollerar en systemleverantör, såväl som varje lufttrafikföretag som det äger eller effektivt kontrollerar.
j) effektiv kontroll: ett förhållande som bygger på rättigheter, avtal eller andra grunder, som antingen var för sig eller tillsammans och med hänsyn till faktiska omständigheter och berörda rättsregler, ger en möjlighet att direkt eller indirekt utöva ett avgörande inflytande över ett företag, i synnerhet genom
P rättigheten att förfoga över alla eller en del av företagets tillgångar,
P rättigheter eller avtal som ger ett avgörande inflytande över sammansättningen hos företagets organ, omröstning eller andra beslut, eller som på annat sätt ger ett avgörande inflytande över driften av ett företag.
k) deltagande lufttrafikföretag: ett lufttrafikföretag som har ett avtal med en systemleverantör om förmedling av sina lufttransportprodukter genom ett datoriserat bokningssystem. I den utsträckning som ett moderföretag använder tjänsterna i sitt eget datoriserade bokningssystem, som omfattas av denna förordning, betraktas det som ett deltagande lufttrafikföretag.
l) abonnent: en person eller ett företag som inte är ett deltagande lufttrafikföretag och som enligt avtal eller annan överenskommelse med en systemleverantör använder ett datoriserat bokningssystems distributionstjänster för försäljning av lufttransportprodukter.
m) konsument: varje person som önskar upplysning om eller har för avsikt att köpa en lufttransportprodukt.
n) primär textbild: en textbild som ger omfattande och opartisk information om flygförbindelser mellan två orter inom en angiven tidsperiod.
o) restid: skillnaden mellan tidtabellsenlig avgångs- och ankomsttid.
p) serviceförbättring: varje produkt eller tjänst som inte är en distributionstjänst och som en systemleverantör på egna vägnar erbjuder abonnenter i anslutning till ett datoriserat bokningssystem.
Artikel 3
knyta oskäliga villkor till ett avtal med ett deltagande lufttrafikföretag,
fordra att tilläggsvillkor godtas, som genom sin karaktär eller enligt affärssed inte har något samband med deltagandet i leverantörens datoriserade bokningssystem, och skall tillämpa samma villkor för samma servicenivå.
b) En systemleverantör får inte ställa som villkor för att få delta i leverantörens datoriserade bokningssystem att ett deltagande lufttrafikföretag inte samtidigt deltar i ett annat system.
c) Ett deltagande lufttrafikföretag skall ha rätt att säga upp sitt avtal med en systemleverantör med en uppsägningstid som inte behöver överstiga sex månader, dock att den tidigast får löpa ut vid utgången av det första avtalsåret.
I sådana fall skall en systemleverantör bara ha rätt att få tillbaka de direkta kostnaderna för uppsägningen av avtalet.
4. Om en systemleverantör avser att förbättra de distributionstjänster han erbjuder eller den utrustning som används i samband med att dessa tjänster erbjuds, skall han erbjuda samtliga deltagande lufttrafikföretag, inklusive moderföretag, information om och möjlighet att få del av dessa förbättringar med samma skyndsamhet, på samma villkor och under samma förutsättningar med förbehåll för de tekniska begränsningar som ligger utanför systemleverantörens kontroll, och på ett sådant sätt att det inte är någon skillnad i tidsförloppet för genomförandet av de nya förbättringarna mellan moderföretag och deltagande lufttrafikföretag."
2. Följande artikel skall läggas till:
"Artikel 3a
1. a) Ett moderföretag får inte diskriminera ett konkurrerande datoriserat bokningssystem genom att vägra att ge det senare, på begäran och med samma skyndsamhet, samma information om tidtabeller, biljettpriser och platstillgång avseende dess egna flygförbindelser, som det ger sitt eget datoriserade bokningssystem, eller att vägra distribuera sina lufttransportprodukter genom ett annat datoriserat bokningssystem, eller att vägra acceptera eller med samma skyndsamhet bekräfta en bokning som görs från ett konkurrerande datoriserat bokningssystem avseende dess egna lufttransportprodukter som det distribuerar genom sitt eget datoriserade bokningssystem. Moderföretaget skall bara vara förpliktat att acceptera och bekräfta de bokningar som överensstämmer med dess biljettpriser och villkor.
1. b) Moderföretaget skall inte vara förpliktat att acceptera några kostnader i samband med detta utom för återgivande av den information som skall ges och för accepterade bokningar.
1. c) Moderföretaget skall ha rätt att utföra kontroller för att säkerställa att artikel 5.1 respekteras av det konkurrerande datoriserade bokningssystemet.
2. Skyldigheten enligt denna artikel skall inte gälla till förmån för ett konkurrerande datoriserat bokningssystem när, det enligt förfarandena i artikel 6.5 eller 7.3 och 7.4 har konstaterats att det datoriserade bokningssystemet bryter mot artikel 4a eller att en systemleverantör inte kan ge tillräckliga garantier för att skyldigheterna enligt artikel 6 om moderföretags obehöriga tillgång till information uppfylls."
3. Artikel 4 skall ersättas med följande:
"Artikel 4
2. En systemleverantör får inte reservera någon specifik dataladdnings- eller databehandlingsmetod eller någon annan distributionstjänst för ett eller flera av sina moderföretag.
3. En systemleverantör skall säkerställa att dess distributionstjänster är avskilda på ett klart och verifierbart sätt från varje lufttrafikföretags privata tjänster rörande platstillgång, företagsledning och avsättning. Åtskillnaden får ske antingen logiskt genom mjukvara eller fysiskt på ett sådant sätt att varje förbindelse mellan distributionstjänsterna och de privata tjänsterna bara uppnås genom ett gränssnitt mellan två tillämpningar. Oavsett metoden för åtskillnad skall ett sådant gränssnitt göras tillgängligt för alla moderföretag och deltagande lufttrafikföretag utan diskriminering samt ge lika behandling avseende procedurer, protokoll, inmatning och utmatning. När relevanta och allmänt accepterade standarder för lufttransportsektorn finns tillgängliga skall systemleverantörerna erbjuda tjänster som är kompatibla med dessa."
1. a) Ett datoriserat bokningssystem skall ge en textbild som är klar och som inte är diskriminerande.
1. b) En systemleverantör får inte avsiktligt eller av oaktsamhet visa oriktig eller vilseledande information i sitt datoriserade bokningssystem.
2. a) En systemleverantör skall via sitt datoriserade bokningssystem tillhandahålla en eller flera primära textbilder för varje enskild transaktion som visar data som inlevererats av deltagande lufttrafikföretag, om tidtabeller, biljettpriser och tillgången på platser för enskilda köpare på ett klart och tillräckligt omfattande sätt som inte är diskriminerande eller partiskt, i synnerhet vad gäller den ordning i vilken informationen presenteras.
1. b) En konsument skall ges möjlighet att begära primära textbilder för enbart regelbunden eller icke-regelbunden lufttrafik.
1. c) Vid presentation på en primär textbild får vid sammanställning och val av flygningar mellan två givna orter ingen diskriminering göras mellan flygplatser som betjänar samma ort.
1. d) Ordningsföljden mellan olika flygmöjligheter på den primära textbilden skall vara den som framgår av bilagan.
1. e) De normer som används för att rangordna informationen får inte baseras på någon faktor som direkt eller indirekt har samband med lufttrafikföretagets identitet och inte tillämpas på ett sätt som diskriminerar något deltagande lufttrafikföretag.
3. När en systemleverantör lämnar information om biljettpriser skall textbilden vara opartisk och icke-diskriminerande och minst innehålla biljettpriserna för alla deltagande lufttrafikföretags flygningar som visas i den primära textbilden. Källan för sådan information skall vara godtagbar för de berörda deltagande lufttrafikföretagen och systemleverantörerna.
4. Information om kombinerade produkter avseende bl.a. vem som organiserar resan, platstillgång och priser skall inte visas i den primära textbilden.
5. Ett datoriserat bokningssystem anses inte bryta mot bestämmelserna i denna förordning i den utsträckning som det förändrar en textbild för att tillmötesgå en konsuments specifika förfrågningar.
Artikel 6
1. Följande bestämmelser skall styra tillgängligheten av den information i form av statistik eller av annat slag, som en systemleverantör erbjuder från sitt datoriserade bokningssystem:
a) Information om enskilda bokningar skall ställas till förfogande på lika villkor för det eller de lufttrafikföretag som deltar i utförandet av den tjänst som bokningen avser och för de abonnenter som berörs av bokningen.
b) Varje upplysning om avsättning, bokningar och försäljning skall ske på grundval av följande:
i) Att uppgifterna erbjuds med samma skyndsamhet och på ett icke-diskriminerande sätt till alla deltagande lufttrafikföretag, inklusive moderföretag.
ii) Att sådana uppgifter får, och skall på begäran, omfatta alla deltagande lufttrafikföretag och abonnenter, men skall inte identifiera eller ge personlig information om en passagerare eller ett företag.
iii) Att alla förfrågningar om sådana uppgifter skall behandlas med samma omsorg och skyndsamhet, med förbehåll för den överföringsmetod som det enskilda lufttrafikföretaget väljer.
2. Personlig information om en passagerare som kommer från ett datoriserat bokningssystem får bara med passagerarens medgivande göras tillgänglig för andra som inte är berörda av transaktionen.
3. Systemleverantören skall säkerställa att bestämmelserna i punkt 1 och 2 uppfylls genom tekniska medel eller lämpliga säkerhetskrav avseende åtminstone mjukvara, på ett sådant sätt att ett eller flera av moderföretagen inte på något sätt kan få tillgång till information som ges av eller skapas för lufttrafikföretag, utom vad som tillåts enligt denna artikel.
4. Systemleverantören skall inom tre månader efter denna förordnings ikraftträdande på begäran ställa till förfogande för alla deltagande lufttrafikföretag en utförlig beskrivning av de tekniska och administrativa åtgärder som han vidtagit för att uppfylla bestämmelserna i denna artikel.
5. Efter att ha mottagit den utförliga beskrivningen av de tekniska och administrativa åtgärder som vidtagits av systemleverantören, skall kommissionen inom tre månader fatta beslut om huruvida åtgärderna är tillräckliga för att uppfylla säkerhetskraven enligt denna artikel. Om så inte är fallet får kommissionen i sitt beslut tillämpa artikel 3a.2. Kommissionen skall genast informera medlemsstaterna om ett sådant beslut. Om rådet, på begäran av en medlemsstat, inte inom två månader efter kommissionens beslut beslutar annorlunda, skall kommissionens beslut träda i kraft."
6. I artikel 7 skall punkterna 1 och 2 ersättas med följande:
"1. Förpliktelserna för en systemleverantör enligt artikel 3 och 4 P6 gäller inte mot ett moderföretag i ett tredje land, i den mån det företagets datoriserade bokningssystem utanför gemenskapens territorium inte erbjuder EG-lufttrafikföretag en behandling som är likvärdig med den som tillämpas enligt denna förordning och enligt kommissionens förordning (EEG) nr 83/91 ().
7. I artikel 7 skall följande punkt läggas till:
"5. a) När det konstateras allvarlig diskriminering enligt punkterna 1 och 2 får kommissionen besluta om att de datoriserade bokningssystemen skall instrueras att ändra sina metoder så att diskrimineringen upphör. Kommissionen skall genast informera medlemsstaterna om ett sådant beslut.
"5. b) Om rådet, på begäran av en medlemsstat, inte inom två månader efter kommissionens beslut beslutar annorlunda, skall kommissionens beslut träda i kraft."
1. Ett moderföretag får inte till en abonnents användning av något visst datoriserat bokningssystem direkt eller indirekt knyta någon provision eller annan förmån eller någon avskräckande åtgärd för att sälja företagets lufttransportprodukter som är tillgängliga på dess flygningar.
2. Ett moderföretag får varken direkt eller indirekt kräva att en abonnent använder ett visst datoriserat bokningssystem för att sälja eller utställa biljetter för en lufttransportprodukt som företaget självt direkt eller indirekt levererar.
3. Ett lufttrafikföretags villkor för att godkänna en resebyrå som sin agent med rätt att sälja och utställa biljetter för företagets lufttransportprodukter skall inte påverka tillämpningen av punkterna 1 och 2."
9. Artikel 9.4, 9.5 och 9.6 skall ersättas med följande:
"4. a) En systemleverantör får inte ställa upp oskäliga villkor i ett avtal med en abonnent om användning av dess datoriserade bokningssystem, och i synnerhet får en abonnent alltid säga upp sitt avtal med en systemleverantör med en uppsägningstid som inte behöver överstiga tre månader, dock att den tidigast får löpa ut vid utgången av det första avtalsåret.
I sådana fall skall en systemleverantör bara ha rätt att få tillbaka de direkta kostnaderna för uppsägningen av avtalet.
"4. b) Med förbehåll för punkt 2 skall leverans av teknisk utrustning inte omfattas av villkoren enligt a.
5. En systemleverantör skall i varje abonnentavtal fastställa
a) att en primär textbild tillhandahålls för varje enskild transaktion enligt artikel 5, utom när en konsument begär information om endast ett lufttrafikföretag, eller när en konsument begär information om endast kombinerade lufttransportprodukter,
b) att abonnenten inte behandlar det material som levereras av de datoriserade bokningssystemen på ett sätt som skulle leda till att konsumenterna får oriktig, vilseledande eller diskriminerande information.
6. En systemleverantör får inte ålägga en abonnent någon skyldighet att acceptera ett erbjudande om teknisk utrustning eller mjukvara, men får kräva att en utrustning eller mjukvara som är kompatibel med hans eget system används."
10. I artikel 10 skall punkterna 1 och 2 ersättas med följande:
"1. De avgifter som begärs av en systemleverantör får inte vara diskriminerande och skall vara rimligt strukturerade och stå i ett rimligt förhållande till anskaffningskostnaden för den tjänst som tillhandahålls och utnyttjas och skall i synnerhet vara desamma för samma servicenivå.
Fakturorna för det datoriserade bokningssystemets tjänster skall vara tillräckligt informativa för att de deltagande lufttrafikföretagen och abonnenterna skall kunna se exakt vilka tjänster de utnyttjat och avgifterna för dem. Fakturor för bokningsavgifter skall minst innehålla följande uppgifter för varje sträcka:
P Typ av bokning i det datoriserade bokningssystemet.
P Passagerarens namn.
P Stat.
P Identifieringskod för IATA/ARC agentur.
P Ortkod.
P De två orterna eller sträckan.
P Bokningsdatum (transaktionsdatum).
P Resdatum.
P Linjenummer.
P Statuskod (bokningsstatus).
P Bokningsnummer (PNR-nummer).
P Boknings-/avbokningsindikator.
Fakturainformationen skall erbjudas på magnetiska medier.
Ett deltagande lufttrafikföretag skall erbjudas möjligheten att bli informerat när det sker en bokning/transaktion för vilken en bokningsavgift kommer att debiteras. Om företaget väljer att bli informerat skall det erbjudas möjligheten att kunna annullera en sådan bokning/transaktion, såvida den inte redan har accepterats.
2. En systemleverantör skall på begäran lämna intresserade parter uppgifter om tillämpade metoder och avgifter, om erbjudna systemtjänster, inklusive gränssnitt, samt om de kriterier för redigering och textbildspresentation som används. Denna bestämmelse förpliktar emellertid inte en systemleverantör att lämna information som är äganderättsligt skyddad, till exempel programvara."
11. Artikel 21 skall ersättas med följande:
"Artikel 21
Bestämmelserna i artikel 5, artikel 9.5 och i bilagan till denna förordning skall inte tillämpas på ett datoriserat bokningssystem som används av ett lufttrafikföretag eller en grupp av lufttrafikföretag i dess eget (deras egna) klart markerade kontor och försäljningsdiskar."
12. Följande artikel skall införas:
"Artikel 21a
1. Systemleverantören skall säkerställa att en oberoende kontrollant övervakar att dess datoriserade bokningssystem är tekniskt förenligt med artiklarna 4a och 6. För detta ändamål skall kontrollanten vid varje tidpunkt beviljas tillträde till de program, metoder, förfaranden och säkerhetskrav som används i de datorer eller datorsystem genom vilka systemleverantören erbjuder sina distributionstjänster. Varje systemleverantör skall minst en gång per år till kommissionen lämna sin kontrollants inspektionsrapport och slutsatser. Denna rapport skall granskas av kommissionen för att utröna om det behöver vidtas åtgärder enligt artikel 11.1.
2. Systemleverantören skall informera deltagande lufttrafikföretag och kommissionen om kontrollantens identitet minst tre månader innan utnämningen bekräftas och minst tre månader före varje årlig återutnämning. Om något av de deltagande lufttrafikföretagen inom en månad efter detta meddelande ifrågasätter kontrollantens förmåga att genomföra sina uppgifter enligt denna artikel, skall kommissionen inom ytterligare två månader och efter samråd med kontrollanten, systemleverantören och varje annan part som hävdar ett legitimt intresse besluta om kontrollanten skall ersättas."
13. Artikel 22 skall ersättas med följande:
"Artikel 22
1. Denna förordning inskränker inte tillämpningen av nationell lagstiftning om säkerhet, allmän ordning eller dataskydd.
2. De som har rättigheter enligt artikel 3.4, 4a, 6 och 21 a får inte avsäga sig dessa rättigheter genom avtal eller på annat sätt."
14. Artikel 23 skall ersättas med följande:
"Artikel 23
1. Rådet skall besluta om revidering av denna förordning senast den 31 december 1997 på grundval av ett förslag från kommissionen vilket skall överlämnas senast den 31 mars 1997 tillsammans med en redogörelse för tillämpningen av denna förordning.
2. Rådet skall se över tillämpningen av artiklarna 4a och 6.3 på grundval av en rapport som kommissionen skall lämna senast vid utgången av 1994."
15. Bilagan skall ersättas med bilagan till denna förordning.
Artikel 2
1. Denna förordning träder i kraft den trettionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
2. De nya artiklarna 3.1 och 5.2 b i förordning (EEG) nr 2299/89 skall inte tillämpas förrän sex månader efter den dag som anges i punkt 1. Kommissionen får bevilja ytterligare 12 månaders uppskov till de datoriserade bokningssystem som av objektiva skäl inte kan uppfylla bestämmelserna i artiklarna 3.1 och 5.2 b.
3. Skyldigheten enligt punkt 9 c i bilagan att visa anslutande flygtrafik med en linje per sträcka skall tillämpas från och med den 1 januari 1995.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
av den 14 december 1993
VERKSTÄLLANDE KOMMITTÉN HAR FATTAT DETTA BESLUT
med beaktande av artikel 132 i konventionen om tillämpning a
RÅDETS BESLUT av den 20 december 1994 om ingående av tilläggsprotokollet till interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Rumänien, å andra sidan, och till Europaavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan (94/48/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113 i förening med artikel 228.2 i detta,
med beaktande av Europeiska rådets slutsatser från mötet i Köpenhamn den 21 och 22 juni 1993,
med beaktande av kommissionens förslag, och
med beaktande av följande: Kommissionen har på gemenskapens vägnar förhandlat fram ett tilläggsprotokoll till interimsavtalet om handel och handelsfrågor och till Europaavtalet med Rumänien.
Detta tilläggsprotokoll bör godkännas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Tilläggsprotokollet till interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Rumänien, å andra sidan, och till Europaavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan, godkänns på Europeiska gemenskapens vägnar.
Texten till tilläggsprotokollet bifogas detta beslut.
Artikel 2
Rådets ordförande bemyndigas att utse den person som skall ha befogenhet att underteckna tilläggsprotokollet på Europeiska gemenskapens vägnar.
Rådets ordförande skall på Europeiska gemenskapens vägnar göra den anmälan som fastställs i artikel 8 i tilläggsprotokollet.
KOMMISSIONENS BESLUT av den 7 februari 1994 om ändring av rådets beslut 90/424/EEG om vissa utgifter på veterinärområdet (84/77/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets beslut 90/424/EEG av den 26 juni 1990 om vissa utgifter på veterinärområdet(1), senast ändrat genom beslut 93/439/EEG(2), särskilt artikel 24.1 i detta, och med beaktande av följande:
Enligt artikel 24 i beslut 90/424/EEG införs möjligheten att vidta en gemenskapsfinansierad åtgärd för att utrota och övervaka de sjukdomar som finns angivna i förteckningen i bilagan till detta beslut.
Heartwater, babesios och anaplasmos, som överförs av smittbärande insekter, förekommer i de franska utomeuropeiska departementen.
Med hänsyn till den särskilda hälsosituationen i de franska utomeuropeiska departementen är det motiverat att lägga till nämnda sjukdomar i bilagan till beslut 90/424/EEG.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande strecksatser skall läggas till under Grupp 1 i förteckningen i bilagan till beslut 90/424/EEG:
"- Heartwater, som överförs av smittbärande insekter i de franska utomeuropeiska departementen,
- Babesios, som överförs av smittbärande insekter i de franska utomeuropeiska departementen,
- Anaplasmos, som överförs av smittbärande insekter i de franska utomeuropeiska departementen".
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 8 februari 1994 om ändring av rådets direktiv 89/556/EEG om djurhälsovillkor för handel inom gemenskapen med och import från tredje land av embryon från tamdjur av nötkreatur (Text av betydelse för EES) (94/113/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 89/556/EEG av den 25 september 1989 om djurhälsovillkor för handel inom gemenskapen med och import från tredje land av embryon från tamdjur av nötkreatur(1), senast ändrat genom direktiv 93/52/EEG(2), särskilt artikel 16 i detta, och med beaktande av följande:
Genom artikel 1 i direktiv 89/556/EEG utesluts från direktivets räckvidd embryon som är resultatet av vissa tekniker. Handel eller import med embryon som skall underkastas tekniker som innebär att zona pellucida genombryts, och med sådana som är resultatet av befruktning in vitro får ske under förutsättning att de uppfyller kraven i direktiv 89/556/EEG samt vissa kompletterande skyddsåtgärder.
De åtgärder som föreskrivs i det här direktivet är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagorna till direktiv 89/556/EEG skall ändras enligt vad som framgår av bilagan till detta beslut.
Artikel 2
Detta beslut skall tillämpas från och med den 1 mars 1994.
Beslutet skall inte tillämpas på embryon som samlas, hanteras och förvaras före den 1 mars 1994.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 23 februari 1994 om inrättande av en rådgivande samordningskommitté för förebyggande av bedrägerier (94/140/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, och
med beaktande av följande: En sund förvaltning av gemenskapens finanser förutsätter att bedrägerier som skadar gemenskapens budget motarbetas effektivt.
Det är i första hand medlemsstaterna som har ansvaret för riktade åtgärder för bekämpning av bedrägeribrott. Detta kräver ett nära samarbete mellan medlemsstaterna och kommissionen.
Enligt vad som avses i artikel 209a i fördraget skall medlemsstaterna vidta samma åtgärder för att motarbeta bedrägerier som riktar sig mot gemenskapens finansiella intressen som de vidtar för att motarbeta bedrägerier som riktar sig mot deras egna finansiella intressen. Därför måste de med kommissionens hjälp samordna sina insatser för att skydda gemenskapens finansiella intressen och motarbeta bedrägerier.
Kommissionen har även ett stort ansvar som ett led i sin generella uppgift att se till att gemenskapens budget tillämpas korrekt och att fördragets bestämmelser genomförs.
Kommissionen bör därför kunna rådfråga en kommitté bestående av företrädare för medlemsstaterna, vilken kan rådfrågas om alla frågor som rör förebyggande verksamhet, samarbete mellan medlemsstaterna och kommissionen, bekämpning av bedrägeribrott samt alla andra frågor med anknytning till det rättsliga skyddet för gemenskapens finansiella intressen.
De befintliga kommittéernas arbetsuppgifter är begränsade till särskilda områden. Dessa kommittéer ersätts inte. Det finns dock behov av att få en samlad överblick över problematiken när det gäller bedrägerier som riktar sig mot gemenskapens budget. Därför bör en kommitté inrättas som kan behandla hela bedrägeriproblematiken.
Eftersom kommittén kommer att behandla alla aspekter av bedrägeriproblematiken och alla medlemsstater har behov av en representation på rätt nivå som avspeglar strukturen i den egna förvaltningen, bör det läggas fast att kommittén skall bestå av två företrädare från varje medlemsstat.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
1. Kommittén skall bestå av två företrädare för varje medlemsstat, vilka får biträdas av två tjänstemän från de berörda myndigheterna.
2. Kommittén skall ha en företrädare för kommissionen som ordförande.
3. Arbetsgrupper kan inrättas för att underlätta kommitténs arbete.
2. Kommissionen kan när den begär ett yttrande från kommittén fastställa en tidsfrist för avgivande av yttrandet.
3. De synpunkter som lagts fram av företrädarna för medlemsstaterna skall föras till protokollet.
RÅDETS BESLUT av den 19 april 1994 om en av rådet enligt artikel J 3 i Fördraget om den Europeiska unionen beslutad gemensam åtgärd till stöd för fredsprocessen i Mellanöstern (94/276/GUSP)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om Europeiska unionen, särskilt artiklarna J 3 och J 11 i detta,
med beaktande av de allmänna riktlinjer som utfärdades av Europeiska rådet den 29 oktober 1993,
med beaktande av ramen för den gemensamma åtgärd som Europeiska rådet enades om den 10 och 11 december 1993, och
med beaktande av artikel C i Fördraget om Europeiska unionen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
a) I syfte att verka för att en heltäckande fred i Mellanöstern sluts på grundval av FN:s säkerhetsråds resolutioner skall Europeiska unionen
- delta i de internationella arrangemang som parterna kommer överens om för att säkerställa fred inom ramen för den process som startades i Madrid,
- använda sitt inflytande för att uppmuntra alla parter att ovillkorligt stödja fredsprocessen på grundval av inbjudningar till Madrid-konferensen och arbeta för att stärka demokratin och respekten för de mänskliga rättigheterna,
- bidra till utformningen av de framtida förbindelserna mellan regionens parter i arbetsgruppen för vapenkontroll och regional säkerhet.
b) Europeiska unionen skall
- utveckla sin roll i den särskilda sambandskommitté som ansvarar för samordningen av internationellt stöd till de ockuperade områdena,
- bevara sin ledande roll i arbetsgruppen för regional ekonomisk utveckling (REDWG) och utveckla sitt deltagande i andra multinationella grupper,
- överväga andra sätt att bidra till regionens utveckling.
c) Europeiska unionen skall
- fortsätta att driva frågan om de förtroendeskapande åtgärder som den har förelagt parterna,
- fortsätta att rikta demarscher till de arabiska staterna i syfte att få till stånd ett slut på bojkotten mot Israel,
- följa utvecklingen vad avser israeliska bosättningar inom samtliga ockuperade områden och fortsätta att rikta demarscher till Israel i denna fråga.
Artikel 2
Rådet skall i enlighet med relevanta gemenskapsförfaranden behandla de förslag som kommissionen lägger fram om
- ett snabbt genomförande av biståndsprogrammen för utveckling av de ockuperade områdena och en palestinsk driftsbudget, i nära samråd med palestinierna och en lika nära samverkan med andra biståndsgivare,
- lämnande av stöd enligt befintliga riktlinjer till de andra parterna i de bilateral förhandlingarna, allteftersom dessa gör betydande framsteg mot fred.
Artikel 3
För att aktivt och snabbt bidra till att en palestinsk polisstyrka upprättas skall
a) Europeiska unionen lämna bistånd,
b) presidiet i nära samverkan med kommissionen underlätta samordningen genom utbyte av information mellan medlemsstaterna om deras bilaterala bistånd,
c) ett belopp på högst 10 miljoner ecu från gemenskapens budget som en brådskande åtgärd ställas till förfogande som bistånd till upprättandet av en palestinsk polisstyrka.
Artikel 4
Europeiska unionen skall på begäran av parterna medverka till att det palestinska folket skyddas genom tillfällig internationell närvaro på de ockuperade områdena i överensstämmelse med säkerhetsrådets resolution 904 (1994).
De praktiska arrangemangen och den finansiering som följer av denna artikel skall behandlas i ett särskilt, separat beslut.
Artikel 5
På begäran av parterna skall Europeiska unionen genomföra ett samordnat program för bistånd till förberedelse och övervakning av de val på de ockuperade områdena som påbjöds i principdeklarationen av den 13 september 1993. De exakta praktiska arrangemangen och finansieringen skall fastställas i ett särskilt rådsbeslut när Israel och PLO har enats om hur valet skall arrangeras. Europaparlamentet kommer att inbjudas att delta i dessa arrangemang.
Artikel 6
Europeiska unionen bekräftar att den är villig att fatta ytterligare praktiska beslut inom ramen för denna gemensamma åtgärd allteftersom fredsprocessen utvecklas.
Artikel 7
Detta beslut skall ha verkan från och med denna dag.
Artikel 8
Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS BESLUT av den 25 maj 1994 om tillämpningsföreskrifter till rådets direktiv 90/425/EEG vad avser provtagningen i samband med veterinärkontroller på bestämmelseorten (94/338/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden(1), senast ändrat genom direktiv 92/118/EEG(2), särskilt artikel 5.3 i detta, och med beaktande av följande:
Den behöriga myndigheten i medlemsstaterna får, med användning av icke-diskriminerande veterinära stickprovskontroller på bestämmelseorterna för djur och produkter, kontrollera att de krav som fastställs i artikel 3 i direktiv 90/425/EEG är uppfyllda. Myndigheten får samtidigt utföra provtagning i enlighet med artikel 5.1 a.
För att säkerställa att kontrollerna på bestämmelseorten utförs effektivt, och för att förhindra att det senare uppstår svårigheter i handeln inom gemenskapen, bör det, samtidigt som de berörda parternas intressen skyddas, fastställas vissa närmare bestämmelser om provtagningen.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
RÅDETS BESLUT av den 24 oktober 1994 om utsträckning av det rättsliga skyddet för kretsmönster i halvledarprodukter till personer från Canada (94/700/EG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 87/54/EEG av den 16 december 1986 om rättsligt skydd för kretsmönster i halvledarprodukter(1), särskilt artikel 3.7 i detta,
med beaktande av kommissionens förslag, och
med beaktande av följande: Rätten till rättsligt skydd för kretsmönster i halvledarprodukter i gemenskapen gäller för personer som har rätt till skydd i enlighet med artikel 3.1-3.5 i direktiv 87/54/EEG.
Rätten till skydd kan genom ett rådsbeslut utsträckas till personer som inte åtnjuter skydd genom de nämnda bestämmelserna.
Beslut om utsträckning av skyddet bör i största möjliga omfattning fattas av gemenskapen som helhet.
Detta skydd har tidigare, baserat på ömsesidighet, beviljats personer från vissa länder och territorier utanför gemenskapen, i vissa fall permanent, genom beslut 90/510/EEG(2), i andra interimistiskt, genom beslut 93/16/EEG(3).
Canada har bestämmelser som ger lämpligt skydd till kretsmönsterskapare och landet har tillkännagett att man planerar att uträcka tillämpningen av dessa bestämmelser från och med den 1 november 1994 till att omfatta gemenskapsmedborgare och fysiska och juridiska personer som bedriver verklig och stadigvarande verksamhet i gemenskapen i syfte att skapa kretsmönster eller tillverka integrerade kretsar.
I avtalet om handelsrelaterade aspekter på immateriella rättigheter, som är ett av förhandlingsresultaten i de multilaterala handelsförhandlingarna under Uruguay-rundan och ingår i Marrakesh-slutakten av den 15 april 1994, krävs det att medlemmarna skall ge skydd åt mönster i integrerade kretsar enligt bestämmelserna i det avtalet och bestämmelserna i konventionen om skydd av immateriella rättigheter beträffande integrerade kretsar, till vilket avtalet hänvisar.
Detta avtal och avtalet om inrättandet av Världshandelsorganisationen kommer att träda i kraft den 1 januari 1995 eller snarast möjligt efter den dagen. De industrialiserade länder som är parter i avtalet om inrättandet av Världshandelsorganisationen kommer att ha en frist av ett år efter det avtalets ikraftträdande för att genomföra bestämmelserna i avtalet om handelsrelaterade aspekter på immateriella rättigheter.
Med tanke på de kanadensiska myndigheternas åtaganden bör rätten till skydd enligt direktiv 87/54/EEG utsträckas, från och med den 1 november 1994 till dess bestämmelserna i avtalet om handelsrelaterade aspekter på immateriella rättigheter har genomförts, till att omfatta fysiska personer, bolag och andra juridiska personer från Canada.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Medlemsstaterna skall utsträcka det skydd som avses i direktiv 87/54/EEG enligt följande:
a) Fysiska personer som är medborgare i Canada eller som har sin vanliga vistelseort inom Canadas territorium skall behandlas som om de vore medborgare i en medlemsstat.
b) Bolag eller andra juridiska personer från Canada som bedriver verklig och stadigvarande industriell eller affärsmässig verksamhet i Canada skall behandlas som om de bedrev verklig och stadigvarande industriell eller affärsmässig verksamhet inom en medlemsstats territorium.
Artikel 2
Detta beslut skall tillämpas från och med den 1 november 1994.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 30 november 1994 om särskilda villkor för import av levande tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar med ursprung i Turkiet (Text av betydelse för EES) (94/777/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/492/EEG av den 15 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av levande tvåskaliga blötdjur(1), särskilt artikel 9 i detta, och
med beaktande av följande: En expertgrupp från kommissionen har gjort ett inspektionsbesök i Turkiet för att undersöka under vilka förhållanden levande tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar produceras och släpps ut på marknaden.
Enligt turkisk lagstiftning ansvarar Ministry of Agriculture and Rural Affairs för hälsokontrollen av levande tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar samt för övervakningen av de hygieniska och sanitära förhållandena vid produktionen. Enligt samma lagstiftning är Ministry of Agriculture and Rural Affairs bemyndigad att tillåta eller förbjuda upptagning av tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar i vissa områden.
Ministry of Agriculture and Rural Affairs och dess laboratorier kan effektivt kontrollera tillämpningen av gällande lagar i Turkiet.
De behöriga turkiska myndigheterna har åtagit sig att regelbundet och snabbt till kommissionen överlämna uppgifter om förekomsten av plankton som innehåller toxiner i upptagningsområdena.
De behöriga myndigheterna i Turkiet har officiellt garanterat att de krav som anges i kapitel V i bilagan till direktiv 91/492/EEG och att krav som motsvarar de som föreskrivs i det direktivet vad avser klassificering av upptagnings- och återutläggningsområden, godkännande av leveransanläggningar, hygienkontroll och övervakning av produktionen uppfylls. Kommissionen skall framför allt underrättas om alla eventuella ändringar av upptagningsområdena.
Turkiet kan tas upp i den förteckning över tredje länder som uppfyller de bestämmelser om likvärdighet som anges i artikel 9.3 a i direktiv 91/492/EEG.
I enlighet med artikel 9.3 c i direktiv 91/492/EEG bör en förteckning upprättas över de anläggningar från vilka import av tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar är tillåten. Anläggningar får tas upp i förteckningen endast om de är officiellt godkända av de behöriga myndigheterna i Turkiet. Det åligger de behöriga turkiska myndigheterna att se till att bestämmelserna i artikel 9.3 c i direktiv 91/492/EEG följs.
De särskilda importvillkoren påverkar inte tillämpningen av de beslut som fattas enligt rådets direktiv 91/67/EEG av den 28 januari 1991 om djurhälsovillkor för utsläppande på marknaden av djur och produkter från vattenbruk(2).
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
3. De skall vara förpackade i förseglade förpackningar av en godkänd leveransanläggning som är upptagen i förteckningen i bilaga C.
4. Varje förpackning skall ha en beständig hälsomärkning som innehåller minst följande uppgifter:
- Avsändande land: TURKIET.
- Art (gängse och vetenskapligt namn).
- Uppgift om upptagningsområdets och leveransanläggningens godkännandenummer.
- Förpackningsdatum med angivande av minst dag och månad.
Artikel 3
1. Intygen enligt artikel 2.1 skall vara utfärdade på minst ett officiellt språk i den medlemsstat där kontrollerna görs.
2. Intygen skall innehålla namn, tjänsteställning och underskrift av den veterinär som representerar Ministry of Agriculture and Rural Affairs och dettas officiella stämpel i en annan färg än den som använts för övriga noteringar.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 16 december 1994 om särskilda villkor för godkännandet av de förpackningsanläggningar som avses i rådets direktiv 77/99/EEG och om bestämmelser om saluhållandet av produkter därifrån (94/837/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De hygienvillkor som skall gälla för sådan verksamhet bör fastställas.
Bestämmelserna om kontrollmärkning av produkter från sådana förpackningsanläggningar bör fastställas.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Förpackningsanläggningar som endast plockar samman produkter utan att ta bort innerförpackningen skall uppfylla tillämpliga villkor enligt bilaga B, kapitel VII punkt 1 till direktiv 77/99/EEG.
2. Förpackningsanläggningar som tar bort innerförpackningen och förser produkterna med ny innerförpackning skall uppfylla gällande villkor enligt bilaga A, kapitlen I och II till direktiv 77/99/EEG och de relevanta villkoren enligt bilaga B, kapitel I punkterna 1 a, 1 b, 1 d, 1 e och 1 f samt 2 a, 2 c, 2 i och 2 j till ovannämnda direktiv.
Artikel 2
1. Produkter från de förpackningsanläggningar som avses i artikel 1.1 skall bibehålla kontrollmärket från det ursprungliga produktionsföretaget.
Produkter från de förpackningsanläggningar som avses i artikel 1.2 skall märkas med ett kontrollmärke i enlighet med de bestämmelser som fastställs i bilaga B, kapitel VI till direktiv 77/99/EEG. Den behöriga myndigheten skall tilldela förpackningsanläggningarna ett kontrollmärke.
Om produkter från olika produktionsföretag plockas samman skall förpackningsanläggningens kontrollmärke åsättas det yttersta emballaget som produkterna paketeras i på förpackningsanläggningen.
2. Förpackningsanläggningar skall upprätta ett särskilt registreringssystem som gör det möjligt för den behöriga myndigheten att spåra en ompaketerad produkt till ursprungsföretaget.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 28 december 1994 om godkännande av Finlands operativa program för bekämpning av salmonella hos vissa levande djur och i animaliska produkter (94/968/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 64/432/EEG av den 26 juni 1964 om djurhälsoproblem som påverkar handeln inom gemenskapen med nötkreatur och svin(1), ändrat genom del 1 kapitel 2 avsnitt A punkt 1. h i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 10a andra stycket i detta,
med beaktande av rådets direktiv 90/539/EEG av den 15 oktober 1990 om djurhälsoproblem för handeln inom gemenskapen med och import av fjäderfä och kläckningsägg från tredje land(2), ändrat genom del 1 kapitel 2 avsnitt A punkt 4. b och 4. c i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 9a, 9b och 10b i detta,
med beaktande av rådets direktiv 64/433/EEG av den 26 juni 1964 om hälsoproblem som påverkar handeln med färskt kött inom gemenskapen(3), ändrat genom del 1 kapitel 3 punkt 1. d i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 5.4 i detta,
med beaktande av rådets direktiv 71/118/EEG av den 15 februari 1971 om hälsoproblem som påverkar handeln med färskt fjäderfäkött(4), ändrat genom del 1 kapitel 3 punkt 3. b i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 5.4 i detta,
med beaktande av rådets direktiv 92/118/EEG av den 17 december 1992 om djurhälso- och hygienkrav för handel inom gemenskapen med produkter som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A. I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG, samt för import till gemenskapen av sådana produkter(5), ändrat genom del 1 kapitel 4 punkt 4. c i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt kapitel 2 första strecksatsen i bilaga 2 till denna, och med beaktande av följande:
Den 10 oktober och den 13 december 1994 förelade Finland kommissionen sitt operativa program för bekämpning av salmonella i enlighet med artikel 10a.2 i direktiv 64/432/EEG, artiklarna 9a, 9b och 10b i direktiv 90/539/EEG, artikel 5 i direktiv 64/433/EEG, artikel 5 i direktiv 71/118/EEG och första strecksatsen i kapitel 2 i bilaga 2 till direktiv 92/118/EEG.
Detta operativa program omfattar alla de åtgärder som Finland från och med dagen för ikraftträdandet av anslutningsfördraget har åtagit sig att vidta för att bekämpa salmonella hos nötkreatur och svin för avel, produktion och slakt, avelsfjäderfä, daggamla kycklingar som skall ingå i flockar av avelsfjäderfä eller flockar av produktionsfjäderfä, värphöns (produktionsfjäderfä som föds upp för att producera konsumtionsägg), slaktfjäderfä, nötkött och griskött, fjäderfäkött och ägg till direkt konsumtion som livsmedel.
Mot bakgrund av detta bör endast ett kommissionsbeslut antas om godkännande av det operativa programmet.
De salmonellagarantier som gäller för Finland, redan fastställda eller som kommer att fastställas i framtiden, skall specificeras för varje kategori av levande djur och animaliska produkter. Tillämpningen av nämnda garantier är beroende av att de åtgärder som Finland skall vidta inom varje sektor godkänns.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Det finska programmets åtgärder avseende nötkreatur och svin för avel, produktion och slakt godkänns.
Artikel 2
Det finska programmets åtgärder avseende avelsfjäderfä och dagsgamla kycklingar som skall ingå i flockar av avelshöns eller flockar av produktionsfjäderfä godkänns.
Artikel 3
Det finska programmets åtgärder avseende värphöns (produktionsfjäderfä som föds upp för att producera konsumtionsägg) godkänns.
Artikel 4
Det finska programmets åtgärder avseende slaktfjäderfä godkänns.
Artikel 5
Det finska programmets åtgärder avseende nötkött och svinkött godkänns.
Artikel 6
Det finska programmets åtgärder avseende fjäderfäkött godkänns.
Artikel 7
Det finska programmets åtgärder avseende ägg för direkt konsumtion som livsmedel godkänns.
Artikel 8
Finland skall på dagen för ikraftträdandet av anslutningsfördraget sätta i kraft de lagar och andra författningar som är nödvändiga för att vidta de åtgärder som avses i artiklarna 1, 2, 3, 4, 5, 6 och 7.
Artikel 9
Detta beslut träder i kraft om och på samma dag som anslutningsfördraget för Norge, Österrike, Finland och Sverige träder i kraft.
Artikel 10
Detta beslut riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EEG) nr 163/94 av den 24 januari 1994 om ändring av förordning (EEG) nr 386/90 om kontroll i samband med export av jordbruksprodukter som berättigar till exportbidrag eller andra belopp
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2), och
med beaktande av följande: Enligt rådets förordning (EEG) nr 386/90 av den 12 februari 1990 om kontroll i samband med export av jordbruksprodukter som berättigar till exportbidrag eller andra belopp(3), måste kommissionen för rådet framlägga en rapport om framstegen i tillämpningen av förordningen.
Det framgår klart av denna rapport och av tilläggsrapporten att den bristande smidigheten hos vissa regler kan motverka förbättringar av effektiviteten i kontrollerna; riskanalyser kan komma till bättre användning om kontrollorganen har större frihet att själva bestämma på vilka områden det särskilt skall genomföras kontroller.
Förpliktelsen att uppfylla en procentsats på 5 % per sektor och per tullkontor gör det svårare att koncentrera personella resurser på export med hög risk.
Generellt sett bör kontrollsatsen ligga kvar på 5 %, men ordningen kan göras smidigare, så att kontrollorganen kan koncentrera sina insatser på känsligare produkter.
För att minska risken för utbyte av produkter, särskilt när det gäller exportdeklarationer som framläggs och godkänns inne i medlemsstaten eller i exportörens lokaler måste det fastställas en lägsta procentsats av representativa fysiska stickprovskontroller som skall genomföras vid utförseltullkontoret.
Med tanke på nödvändigheten av att bestämmelserna om kontroll av exportbidrag tillämpas effektivt överallt i gemenskapen och mot bakgrund av de ekonomiska riskerna för gemenskapens tillgångar, måste regler antas på gemenskapsnivå.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 386/90 ändras på följande sätt:
- per tullkontor,
- per kalenderår, och,
- per produktsektor.
Procentsatsen på 5 % per produktsektor kan dock ersättas med en procentsats på 5 % för samtliga sektorer, förutsatt att medlemsstaten tillämpar ett urvalssystem baserat på riskanalys vilken utförs enligt kriterier som närmare skall fastställas i enlighet med det förfarande som anges i artikel 6. I så fall är en lägsta procentsats på 2 % per produktsektor obligatorisk."
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1966/94 av den 28 juli 1994 om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom kommissionens förordning (EG) nr 1737/94(2), särskilt artikel 9 i denna, och med beaktande av följande:
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovanstående förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
Om inte annat följer av de åtgärder som är i kraft i gemenskapen beträffande system med dubbelkontroll och med övervakning i för- och efterhand av import av textilprodukter till gemenskapen, är det lämpligt att de bindande klassificeringsbesked som getts ut av medlemsstaternas tullmyndigheter rörande klassificeringen av varor i Kombinerade nomenklaturen och som inte överensstämmer med denna förordning, fortsatt får åberopas av mottagaren under en tid av 60 dagar, enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3).
Beträffande produkterna nr 3, 5, 6 och 7 i bifogade tabell har Tullkodexkommitténs sektion för tulltaxe- och statistiknomenklatur inte avgivit något yttrande inom den tid som dess ordförande bestämt.
Beträffande produkterna nr 1, 2 och 4 i bifogade tabell är de åtgärder som föreskrivs i denna förordning förenliga med yttrandet från Tullkodexkommitténs sektion för tulltaxe- och statistiknomenklatur.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Om inte annat följer av de åtgärder som gäller i gemenskapen beträffande system med dubbelkontroll och med övervakning i för- och efterhand av import av textilprodukter till gemenskapen, får de bindande klassificeringsbesked som getts ut av medlemsstaternas tullmyndigheter rörande klassificeringen av varor i Kombinerade nomenklaturen och som inte överensstämmer med denna förordning, fortsatt åberopas av mottagaren enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en tid av 60 dagar.
Artikel 3
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2701/94 av den 7 november 1994 om ändring av bilagorna 1, 2, 3 och 4 till rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), senast ändrad genom kommissionens förordning (EG) nr 1430/94(2), särskilt artikel 6-8 i denna, och
med beaktande av följande: Sedan förordningen antogs har bilagorna ändrats ett antal gånger. På grund av ändringarnas antal, komplexitet och det faktum att de är spridda i olika nummer av Europeiska gemenskapernas officiella tidning är texterna svåra att använda och saknar den klarhet som bör vara utmärkande för all lagstiftning. De bör därför kodifieras. Samtidigt bör namnen på eller de kemiska beteckningarna för vissa föreningar rättas till eller preciseras och några sakfel korrigeras.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för anpassning till tekniska framsteg av direktiven om avskaffande av tekniska handelshinder inom sektorn veterinärmedicinska läkemedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagorna 1, 2, 3 och 4 till förordning (EEG) nr 2377/90 ändras på det sätt som anges i bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den sextionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 3129/94 av den 20 december 1994 om ändring av förordning (EEG) nr 2273/93 om fastställande av interventionsorter för spannmål till följd av Österrikes, Finlands och Sveriges anslutning
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Anslutningsakten för Norge, Österrike, Finland och Sverige(1), särskilt artikel 169.2 i denna, och
med beaktande av följande: Kommissionens förordning (EEG) nr 2273/93(2), ändrad genom förordning (EG) nr 2202/94(3), som gäller från och med den 1 januari 1995, skall ändras så att den överensstämmer med bestämmelserna i anslutningsakten.
Enligt artikel 2.3 i anslutningsfördraget(4) kan Europeiska unionens institutioner före anslutningen fatta de beslut som avses i artikel 169 i anslutningsakten, varvid dessa beslut träder i kraft om och när detta fördrag träder i kraft.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 2273/93 skall ändras på följande sätt: De interventionsorter med tillhörande upplysningar som anges i bilagan till denna förordning skall läggas till i bilagan till förordning (EEG) nr 2273/93.
Artikel 2
Denna förordning träder i kraft om och när Anslutningsfördraget för Norge, Österrike, Finland och Sverige träder i kraft.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS BESLUT av den 10 februari 1995 om fastställande av särskilda villkor för import av fiskeri- och vattenbruksprodukter från Marocko (Text av betydelse för EES) (95/30/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av fiskeriprodukter (1), särskilt artikel 11.1 i detta, och med beaktande av följande:
En grupp sakkunniga från kommissionen har företagit en resa till Marocko för att försäkra sig om villkoren för produktion, lagerhållning och sändning av fiskeriprodukter avsedda för gemenskapen.
De rättsliga bestämmelser som gäller i Marocko för hälsobesiktning och -kontroll av fiskeriprodukter kan anses vara likvärdiga med dem som fastställs i direktiv 91/493/EEG.
Direction de l'élevage, ministère de l'agriculture (DEMA) i Marocko är i stånd att på ett effektivt sätt kontrollera tillämpningen av den gällande lagstiftningen.
De villkor som gäller det intyg som avses i artikel 11.4 a i direktiv 91/493/EEG omfattar fastställandet av en förlaga till ett intyg, valet av det eller de språk som intyget skall vara avfattat på samt firmatecknarens tjänsteställning.
I enlighet med artikel 11.4 b i direktiv 91/493/EEG är det viktigt att på fiskeriprodukternas förpackningar fästa ett märke som anger namnet på det tredje land som avses och ursprungsanläggningens godkännandenummer.
I enlighet med artikel 11.4 c i direktiv 91/493/EEG är det viktigt att fastställa en förteckning över godkända anläggningar. Denna förteckning bör fastställas på grundval av ett meddelande till kommissionen från DEMA. Det åligger således DEMA att förvissa sig om att de villkor som fastställs för detta ändamål i artikel 11.4 i direktiv 91/493/EEG uppfylls.
DEMA har lämnat en officiell försäkran att de bestämmelser som anges i kapitel V i bilagan till direktiv 91/493/EEG och de krav som är likvärdiga med dem som fastställs i det direktivet för godkännande av anläggningar är uppfyllda.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Det intyg som avses i artikel 2.1 bör vara upprättat på minst ett av de officiella språken i den medlemsstat där kontrollen utförs.
2. Intyget bör vara försett med DEMA-ombudets namn, dennes tjänsteställning och underskrift samt med DEMA:s officiella stämpel och allt bör vara i en färg som avviker från de övriga uppgifter som finns på intyget.
Artikel 4
Detta beslut tillämpas från och med den 1 mars 1995.
Artikel 5
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EG) nr 1368/95 av den 16 juni 1995 om ändring av förordning (EEG) nr 2921/90 om beviljande av stöd för framställningen av kasein och kaseinater av skummjölk
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter (1), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94 (2), särskilt artikel 11.3 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 2921/90 ändras på följande sätt:
1. Artikel 2.1 skall ersättas med följande:
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1442/95 av den 26 juni 1995 med ändring av bilagorna I, II, III och IV i rådets förordning (EEG) nr 2377/90 som upprättar ett gemenskapsförfarande för fastställande av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 som upprättar ett gemenskapsförfarande för fastställande av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (1), vilket tidigare omformulerats genom kommissionens förordning (EEG) nr 1441/95 (2), särskilt artikel 6, 7 och 8 i denna, och
med beaktande av följande: I överensstämmelse med förordning (EEG) nr 2377/90 måste gränsvärden fortlöpande fastställas för högsta tillåtna restmängder för alla i gemenskapen använda farmakologiskt verkande substanser i veterinärmedicinska läkemedel avsedda att tillföras livsmedelsproducerande djur.
Gränsvärden för högsta tillåtna restmängder bör endast fastställas sedan prövningar gjorts av Kommittén för veterinärmedicinska läkemedel av all relevant information om den berörda substansens restmängder vad beträffar säkerheten för konsumenten av livsmedel med animaliskt ursprung samt restmängdernas inverkan på industriell förädling av livsmedel:
Det vid fastställandet av gränsvärden för högsta tillåtna restmängder vad gäller restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung är det nödvändigt att klargöra i vilken djurart restmängder förefinnes, såväl den befintliga mängden i samtliga berörda köttvävnader härrörande från det behandlade djuret (målvävnad), som vilken sorts restmängd, vilket är av betydelse vid kontrollen av restmängder (restmängd markör).
För kontrollen av restmängder bör vanligtvis gränsvärden för högsta tillåtna restmängder för målvävnaderna lever eller njure fastställas, för vilket är ombesörjt i tillämplig gemenskapslagstiftning; och med hänsyn till att levern och njuren emellertid ofta avlägsnas från djurkroppen vid transport inom internationell handel, bör gränsvärden för högsta tillåtna restmängder alltid fastställas även för muskel- eller fettvävnad.
Vad gäller veterinärmedicinska läkemedel avsedda för värpfåglar, mjölkdjur och honungsbin, måste gränsvärden för högsta tillåtna restmängder även för ägg, mjölk och honung fastställas.
Carazolol, diazinon och spiramycin (gäller nöt och kyckling) skulle tillföras bilaga I till förordning (EEG) nr 2377/90.
Lecirelin, natrium dikloroisocyanurat, dinoprost trometamin, saltsyra, äpplesyra, l-vinsyra och dess en- och tvåbasiska salter av natrium, kalium och kalcium, bensylalkohol, etanol, n-butanol bör bilaga II tillföras till förordning (EEG) nr 2377/90.
För att möjliggöra komplettering av vetenskapliga studier danofloxacin och erytromycin bör bilaga III föras till förordning (EEG) nr 2377/90.
För att möjliggöra komplettering av vetenskapliga studier, bör giltighetstiden för temporär MRL, tidigare definierad i bilaga III i förordning (EEG) nr 2377/90, förlängas för tylosin och spiramycin (gäller svin).
Då det förefaller som om resthalter av MRL, vid vilken nivå som helst, i livsmedel av animaliskt ursprung utgör hälsorisk för konsumenten, bör furazolidon därför föras till bilaga IV i förordning (EEG) nr 2377/90,
Denna förordning bör träda i kraft efter en period på 60 dagar, för att möjliggöra för medlemsländerna att föra de justeringar av tillstånden som kan komma att bli nödvändiga, samt för att få ut de berörda veterinärmedicinska läkemedlen på marknaden, vilket beviljats i överensstämmelse med rådets direktiv 81/851/EEG (3), senast ändrat genom direktiv 93/40/EEG (4), vilket tar hänsyn till denna förordnings bestämmelser.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för anpassning till tekniska framsteg av direktiven för avskaffande av tekniska handelshinder inom sektorn veterinärmedicinska läkemedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I, II, III och IV i förordning (EEG) nr 2377/90 skall ändras enligt denna förordning.
Artikel 2
Denna förordning träder i kraft den sextionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1662/95 av den 7 juli 1995 om fastställande av vissa närmare föreskrifter för genomförandet av gemenskapens beslutförande för att godkänna utsläppandet på marknaden av humanläkemedel och veterinärmedicinska läkemedel
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2309/93 av den 22 juli 1993 om gemenskapsförfaranden för godkännande för försäljning av och tillsyn över humanläkemedel och veterinärmedicinska läkemedel samt om inrättande av en europeisk läkemedelsmyndighet (1), särskilt artiklarna 10.3 och 32.3 i denna och, med beaktande av följande:
Med stöd av förordning (EEG) nr 2309/93, skall kommissionen anta de bestämmelser som krävs för det skriftliga förfarandet som avses i artiklarna 10.3 och 32.3 i den förordningen.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för humanläkemedel och yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Inom ramen för de beslut som rör tillstånden för utsläppande på marknaden av läkemedel fastställs i denna förordning vissa närmare föreskrifter för hur Ständiga kommittén för humanläkemedel och Ständiga kommittén för veterinärmedicinska läkemedel (nedan kallade "kommittén") skall genomföra det förfarande som föreskrivs i artikel 73 i förordning (EEG) nr 2309/93, i artikel 37b i rådets direktiv 75/319/EEG (2) eller i artikel 42k i rådets direktiv 81/851/EEG (3).
Artikel 2
Ordföranden skall hänskjuta ärenden till kommittén med stöd tillämpliga bestämmelser i förordning (EEG) nr 2309/93, direktiv 75/319/EEG eller direktiv 81/851/EEG.
Utom i undantagsfall, då det förslag till beslut som utarbetats av kommissionen inte är förenligt med yttrandet från Europeiska läkemedelsmyndigheten, skall ett skriftligt förfarande enligt bestämmelserna i artikel 3 tillämpas.
Artikel 3
Inom trettio dagar efter överlämnandet av förslaget till beslut skall medlemsstaterna meddela ordföranden sitt beslut att godkänna förslaget, underkänna det eller avstå från att yttra sig Medlemsstaterna kan komplettera sina beslut med skriftliga anmärkningar. En medlemsstat som inte har meddelat sina invändningar eller sitt beslut att avstå från att yttra sig inom de trettio dagarna anses ha givit förslaget sitt godkännande.
Om en medlemsstat inom tidsfristen på trettio dagar inkommer med en skriftlig begäran, vederbörligen motiverad, om att förslaget till beslut skall behandlas vid ett sammanträde med kommittén skall emellertid det skriftliga förfarandet avslutas, och ordföranden skall snarast möjligt sammankalla kommittén.
Artikel 4
Om kommissionen finner att de skriftliga anmärkningar som lämnats av en medlemsstat inom ramen för förfarandet i artikel 3 väcker betydelsefulla nya frågor av vetenskaplig eller teknisk natur vilka inte har behandlats i Europeiska läkemedelsmyndighetens yttrande, skall ordföranden avbryta förfarandet och kommissionen hänskjuta förslaget till myndigheten för vidare behandling. Ordföranden skall underrätta kommitténs medlemmar om detta.
Ett nytt förfarande skall öppnas inom trettio dagar efter det att kommissionen har mottagit myndighetens svar.
Artikel 5
När en medlemsstat har tillämpat det förfarande som föreskrivs i artikel 18.4 eller 40.4 i förordning (EEG) nr 2309/93 om brådskande tillfälligt förbud mot användning av ett läkemedel inom sitt territorium, skall den tidsfrist som anges i artikel 3 förkortas till femton dagar.
Artikel 6
Om förslaget till beslut skall behandlas vid ett sammanträde med kommittén skall kallelsen, dagordningen och, i fall enligt artikel 2 andra stycket, det förslag till beslut över vilket kommitténs yttrande begärs, av ordföranden överlämnas till medlemmarna i kommittén i enlighet med bestämmelserna i artikel 7.
Dessa handlingar måste nå adressaterna senast tio dagar före sammanträdesdagen eller, i fall enligt artikel 2 andra stycket, en månad före denna dag.
Artikel 7
Korrespondens till medlemmarna i kommittén skall, då kommittén sammanträder enligt det förfarande som avses i artikel 1, sändas genom skriftlig telekommunikation till de behöriga nationella organ som varje medlemsstat utsett för detta ändamål. En kopia skall sändas till den berörda medlemsstatens ständiga representation.
Artikel 8
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100c.3 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande, och
med beaktande av följande: Enligt artikel 100c.3 i Romfördraget skall rådet besluta om åtgärder som syftar till en enhetlig utformning av visumhandlingar före den 1 januari 1996.
Införandet av enhetliga visumhandlingar är ett viktigt steg mot harmoniseringen av viseringspolitiken. Artikel 7a i fördraget fastställer att den inre marknaden skall omfatta ett område utan inre gränser, där fri rörlighet för personer säkerställs i enlighet med bestämmelserna i fördraget. Åtgärden i fråga skall även ses som sammanhängande med de åtgärder som skall antas för tillämpningen av avdelning VI i Fördraget om Europeiska unionen.
Det är väsentligt att den enhetliga modellen för visumhandlingar innehåller alla nödvändiga uppgifter och svarar mot mycket högt ställda tekniska krav, bl.a i fråga om garantier mot efterbildningar och förfalskningar. Den enhetliga modellen måste även vara utformad så att den kan användas i samtliga medlemsstater och innefatta säkerhetsanordningar som är allmänt igenkännliga och kan uppfattas med blotta ögat.
Denna förordning fastställer endast de specifikationer som inte är av konfidentiell art. Dessa specifikationer skall kompletteras med andra som skall förbli hemliga för att förebygga risken för efterbildningar och förfalskningar och som inte får innefatta personliga uppgifter eller hänvisning till sådana. Behörigheten att fastställa andra specifikationer bör tillkomma kommissionen.
För att undvika att uppgifterna i fråga sprids till flera personer än nödvändigt är det också viktigt att endast ett organ i varje medlemsstat utses för tryckningen av den enhetliga visumhandlingen, dock utan hinder av att kunna ersättas av ett annat organ om så behövs. Av säkerhetsskäl skall varje medlemsstat underrätta kommissionen och de övriga medlemsstaterna om det behöriga organets namn.
För att uppnå sitt syfte skall denna förordning vara tillämplig på alla typer av visumhandlingar enligt artikel 5. Medlemsstaterna bör ha möjligheten att använda samma modell för att utfärda visumhandlingar för andra ändamål än de som anges i artikel 5, förutsatt att dessa, på grund av ändringar som kan uppfattas med blotta ögat, inte kan förväxlas med den enhetliga visumhandlingen.
När det gäller de personuppgifter som skall förekomma på den enhetliga visumhandlingen enligt bilagan till denna förordning, skall hänsyn tas till medlemsstaternas bestämmelser om skydd av personuppgifter och till gemenskapslagstiftningen på området.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De visum som beviljas av medlemsstaterna i enlighet med artikel 5 utformas enligt en modell (klistermärke). De skall uppfylla specifikationerna enligt bilagan.
Artikel 2
Kompletterande tekniska specifikationer för att förhindra efterbildningar eller förfalskningar av visumhandlingen skall fastställas i enlighet med förfarandet i artikel 6.
Artikel 3
1. De specifikationer som avses i artikel 2 är hemliga och skall inte offentliggöras. De meddelas enbart till de organ som utses av medlemsstaterna för tryckning och till personer som vederbörligen auktoriserats av en medlemsstat eller av kommissionen.
2. Varje medlemsstat skall utse endast ett organ som ansvarar för tryckningen av visumhandlingar. Namnet på detta organ meddelas till kommissionen och till de övriga medlemsstaterna. Två eller flera medlemsstater får utse samma organ för detta ändamål. Varje medlemsstat får byta detta organ. I så fall skall kommissionen och de andra medlemsstaterna underrättas.
Artikel 4
1. Utan att det påverkar tillämpningen av mer långtgående bestämmelser om skydd av uppgifter har de personer som beviljats ett visum rätt att kontrollera de personuppgifter som finns på visumhandlingen och i förekommande fall att få dessa rättade eller borttagna.
2. Modellen för visumhandlingen innehåller inga andra maskinellt läsbara upplysningar än de som också finns i de rutor som beskrivs i punkterna 6 till 12 i bilagan eller på motsvarande resehandling.
Artikel 5
I denna förordning avses med "visumhandling" ett tillstånd eller beslut av en medlemsstat, som krävs för inresa på dess territorium för
- en vistelse i denna medlemsstat eller i flera medlemsstater för en period som totalt inte överstiger tre månader,
- en resa genom territoriet eller transitzonen på en flygplats i denna medlemsstat eller flera medlemsstater.
Artikel 6
1. När hänvisning sker till förfarandet enligt denna artikel, gäller följande bestämmelser:
2. Kommissionen skall biträdas av en kommitté bestående av företrädare för medlemsstaterna med en företrädare för kommissionen som ordförande.
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över detta förslag inom den tidsfrist som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall anta sitt yttrande med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Vid omröstning inom kommittén skall medlemsstaternas företrädares röster vägas enligt samma artikel. Ordföranden skall inte delta i omröstningen.
3. a) Kommissionen skall anta förslaget om åtgärder om det är förenligt med kommitténs yttrande.
b) Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte har fattat något beslut inom två månader, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas, såvida inte rådet med enkel majoritet har uttalat sig emot förslaget.
Artikel 7
Om medlemsstaterna använder modellen för visumhandling för andra ändamål än dem som omfattas av artikel 5 skall de åtgärder vidtas som behövs för att undvika all förväxling med den visumhandling som beskrivs i artikel 5.
Artikel 8
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS FÖRORDNING (EG) nr 1935/95 av den 22 juni 1995 om ändring i förordning (EEG) nr 2092/91 om ekologisk produktion av jordbruksprodukter och uppgifter därom på jordbruksprodukter och livsmedel
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
med beaktande av följande: Kommissionen har inom ramen för förordning (EEG) nr 2092/91 (4), fått ett särskilt uppdrag att före den 1 juli 1994 göra en förnyad granskning av vissa bestämmelser i nämnda förordning samt att lägga fram lämpliga förslag med tanke på dess eventuella revidering.
Det har visat sig att bestämmelserna om märkning av jordbruksprodukter och livsmedel som innehåller en ingrediens med jordbruksursprung, producerad av odlare eller uppfödare som genomför omläggning av produktionen till ekologiskt jordbruk, som upphör att gälla den 1 juli 1995, bör förlängas för att denna produktion trots sina merkostnader, genom en lämplig märkning av produkterna, skall kunna göras lönande för producenterna.
Den av rådet begärda förnyade granskningen av artiklarna 5, 10 och 11 inför den 1 juli 1994 har visat nödvändigheten av att göra vissa tekniska och redaktionella ändringar i dessa artiklar samt i vissa andra bestämmelser för att kunna garantera en effektiv administrering och tillämpning av förordningen. Utarbetandet av dessa förändrade regler har följaktligen prioriterats och utformningen av regler för animalisk produktion måste därför skjutas upp under en begränsad tid.
Den förnyade granskningen har visat att bestämmelserna om märkning av livsmedel som endast till viss del beretts med hjälp av ingredienser med jordbruksursprung som producerats med ekologiska metoder bör förbättras för att åstadkomma bättre möjligheter att framhäva den ekologiskt producerade beståndsdelen i sådana livsmedel.
Det har också framkommit att den upplysning som anges i bilaga V bör förbli frivillig men att den, för att förhindra missbruk, också bör begränsas till försäljning av färdigförpackade livsmedel eller till direktförsäljning från producent eller beredare till slutkonsumenter med villkor att produktens sammansättning kan identifieras.
Det har dessutom framkommit, att förökningsmaterial bör härröra från ekologiskt odlade växter men att undantagsbestämmelser är nödvändiga för att under en övergångsperiod ge odlarna möjlighet att använda förökningsmaterial som erhållits på konventionellt sätt i fall då det inte finns tillgång till lämpligt material som erhållits enligt ekologiska odlingsmetoder.
Konventionellt erhållna plantor avsedda för växtproduktion bör av samma anledning kunna få användas under en övergångsperiod.
Det har framkommit att vissa av de produkter som användes i enlighet med vedertagna regler för ekologisk odling inom gemenskapen, innan förordning (EEG) nr 2092/91 antogs, inte har inkluderats i bilaga II till nämnda förordning. Användningen av dessa produkter bör tillåtas i den utsträckning som den också är tillåten i det konventionella jordbruket.
Artikel 1
Förordning (EEG) nr 2092/91 ändras på följande sätt:
1. I artikel 1.2 ersätts datumet "den 1 juli 1992" med datumet "den 30 juni 1995."
2. Artikel 4.2 ersätts med följande text:
"2. `produktion`: verksamheter på gården med avseende på framställning, förpackning och ursprunglig märkning som ekologiskt producerade produkter av jordbruksprodukter som produceras på den gården."
3. Artikel 4.3 ersätts med följande text:
"3. `beredning`: åtgärder för konservering och/eller bearbetning av jordbruksprodukter samt förpackning och/eller ändringar av presentationen av det ekologiska produktionsförfarandet som används vid märkningen av de färska konserverade och/eller bearbetade produkterna."
4. Artikel 6.4 ersätts med följande text:
"6. `ingredienser`: ämnen (inbegripet tillsatsämnen) som används vid beredningen av de produkter som avses i artikel 1.1 b såsom de definieras i artikel 6.4 i direktiv 78/112/EEG om tillnärmning av medlemsstaternas lagstiftning om märkning, presentation och reklam i fråga om livsmedel."
5. Följande punkter läggs till i artikel 4:
"9. `färdigförpackat livsmedel`: saluförd enhet såsom den definieras i artikel 1.3 b i direktiv 79/112/EEG,
10. `ingrediensförteckning`: en sådan ingrediensförteckning som avses i artikel 6 i direktiv 79/112/EEG."
6. I artikel 2, artikel 5.1 b, artikel 9.9 a, artikel 11.1 b, artikel 11.2 a och artikel 11.6 a ersätts orden "artikel 6 och 7" med orden "artikel 6".
7. Följande punkt läggs till artikel 5.1:
"d) för produkter som beretts efter den 1 januari 1997, skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som producenten är underställd. Valet av om namn eller kodnummer skall användas vid märkning åligger medlemsstaten som skall meddela sitt beslut till kommissionen."
8. Artikel 5.2 utgår.
9. Artikel 5.3 med följande text:
"3. Vid märkning av och reklam för en produkt som åsyftas i artikel 1.1 b får beskrivningen av den saluförda varan endast innehålla uppgifter som hänvisar till ekologisk produktion om följande villkor är uppfyllda:
a) minst 95 % av produktens ingredienser av jordbruksursprung är produkter eller är framställda ur produkter som har erhållits i enlighet med de regler som fastställs i artikel 6 eller som har importerats från tredje land inom ramen för den ordning som anges i artikel 11,
b) alla andra ingredienser av jordbruksursprung omfattas av bilaga VI punkt C eller har godkänts provisoriskt av ett medlemsland i enlighet med någon av de vidtagna genomförandeåtgärderna, vilken, i förekommande fall, antagits i enlighet med punkt 7,
c) produkten innehåller enbart ämnen som finns förtecknade i bilaga VI punkt a i deras egenskap av ingredienser som inte är av jordbruksursprung,
d) produkten eller dess ingredienser av jordbruksursprung som anges i punkt a har inte behandlats med andra ämnen än de som anges i bilaga VI punkt b,
e) produkten eller dess ingredienser har inte behandlats med joniserande strålning,
f) produkten har beretts eller importerats av en leverantör som är underkastad den kontroll som anges i artiklarna 8 och 9,
g) för produkter som beretts efter den 1 januari 1997 skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som den leverantör som har utfört den sista beredningsåtgärden är underställd. Valet av om namn eller kodnummer skall användas åligger medlemsstaten som skall meddela sitt beslut till kommissionen.
Uppgifter som hänvisar till ekologisk produktion skall klart visa att de gäller en produktionsmetod inom jordbruket och skall åtföljas av en hänvisning till de åsyftade ingredienserna av jordbruksursprung om detta inte klart framgår av ingrediensförteckningen."
10. Artikel 5.4 ersätts med följande text:
"4. Ingredienser av jordbruksursprung får ej förekomma i bilaga VI punkt C annat än när det visas att dessa ingredienser är av jordbruksursprung, att de inte produceras i tillräcklig mängd inom gemenskapen enligt reglerna i artikel 6 eller att de inte kan importeras från tredje land enligt reglerna i artikel 11."
11. Artikel 5.5 ersätts med följande text:
"5. Produkter som är föremål för märkning och reklam i enlighet med styckena 1 och 3 kan vara försedda med uppgifter som hänvisar till omställningen till ekologiskt jordbruk under förutsättning att:
a) de krav som anges i punkt 1 respektive 3 är helt uppfyllda utom vad gäller längden på den övergångsperiod som avses i punkt 1 i bilaga I,
b) en omställningsperiod om minst 12 månader före skörd har iakttagits,
c) uppgifterna inte vilseleder konsumenterna beträffande skillnader i förhållande till produkter som uppfyller alla krav i styckena 1 eller 3. Efter den 1 januari 1996 skall nämnda uppgifter bestå av orden `producerad under omställning till ekologiskt jordbruk` och presenteras i en färg, ett format och i en typstil som inte får vara mer framträdande än beskrivningen av den saluförda varan. Orden `ekologiskt jordbruk` får inte vara mer framträdande än orden `produkt under omställning till`,
d) produkten innehåller en enda ingrediens av jordbruksursprung,
e) för produkter som beretts efter den 1 januari 1997 skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som den leverantör som har utfört den sista beredningsåtgärden är underställd. Valet av om namn eller kodnummer skall användas åligger medlemsstaten som skall meddela sitt beslut till kommissionen."
12. Följande punkt skall införas efter artikel 5.5:
"5a. Utan det påverkar tillämpningen av punkt 3 får sådan märkning av och reklam för en produkt som anges i artikel 1.1 b inte vara försedd med uppgifter som hänvisar till den ekologiska produktionsmetoden annat än om följande villkor är uppfyllda:
a) minst 70 % av produktens ingredienser av jordbruksursprung är produkter eller härrör från produkter som erhållits i enlighet med de regler som anges i artikel 6 eller är importerade från tredje land inom ramen för den ordning som anges i artikel 11,
b) produktens alla andra ingredienser av jordbruksursprung omfattas av bilaga VI punkt C eller har godkänts provisoriskt av en medlemsstat i enlighet med vidtagna genomförandeåtgärder, i förekommande fall i enlighet med punkt 7,
c) uppgifter som hänvisar till ekologisk produktion nämns i ingrediensförteckningen och hänför sig uppenbarligen endast till de ingredienser som erhållits i enlighet med reglerna i artikel 6 eller som importerats från tredje land inom ramen för den ordning som anges i artikel 11. De skall presenteras i en färg, ett format och en typstil som helt överensstämmer med vad som används för övriga uppgifter som finns på ingrediensförteckningen. Dessa uppgifter skall också nämnas separat inom samma synfält som beskrivningen av den saluförda varan och skall innehålla upplysning om den procentuella andel av ingredienserna som är av jordbruksursprung eller som härrör från ingredienser som är av jordbruksursprung och som har erhållits i enlighet med reglerna i artikel 6 eller som importerats från tredje land inom ramen för den ordning som anges i artikel 11. Det nämnda får inte göras i en färg, ett format eller en typstil som gör den mer framträdande än beskrivningen av den saluförda varan. Omnämnandet skall ges följande utformning: `X % av ingredienserna av jordbruksursprung har erhållits i enlighet med reglerna för ekologisk produktion`,
d) produkten innehåller enbart ämnen som finns förtecknade i bilaga VI, punkt A i egenskap av ingredienser som inte är av jordbruksursprung,
e) produkten eller dess ingredienser av jordbruksursprung som anges i punkt a har inte behandlats med andra ämnen än de som finns i bilaga VI punkt B,
f) produkten eller dess ingredienser har inte behandlats med joniserande strålning,
g) produkten har beretts eller importerats av en leverantör som är underkastad den kontroll som anges i artiklarna 8 och 9,
h) för produkter som beretts efter den 1 januari 1997, skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som den leverantör som utfört den sista beredningsåtgärden är underställd. Valet av om namn eller kodnummer skall användas åligger medlemsstaten som skall meddela sitt beslut till kommissionen."
13. Artikel 5.6 ersätts med följande:
"6. Under en övergångsperiod som går ut den 31 december 1997, får märkning av och reklam för en produkt som anges i artikel 1.1 b och som delvis erhållits från ingredienser som inte uppfyller kraven i punkt 3 a hänvisa till ekologisk produktion om följande villkor är uppfyllda:
a) minst 50 % av produktens ingredienser av jordbruksursprung uppfyller kraven i punkt 3 a,
b) produkten uppfyller kraven i punkt 3 c, d, e och f,
c) de uppgifter som hänvisar till ekologisk produktion:
- förekommer uteslutande i ingrediensförteckningen i enlighet med direktiv 79/112/EEG, senast ändrat genom direktiv 89/395/EEG,
- hänför sig uppenbarligen endast till de ingredienser som erhållits i enlighet med de regler som avses i artikel 6, eller som har importerats inom ramen för den ordning som anges i artikel 11,
d) ingredienserna och deras andelar anges i fallande storleksordning efter vikt i ingrediensförteckningen,
e) uppgifterna i ingrediensförteckningen presenteras i samma färg, format och typstil."
14. Inledningen till 5.8 ersätts med följande text:
"8. Sådana begränsande förteckningar över de ämnen och produkter som avses i punkt 3 b, c och d, samt i punkt 5 a, b, d och e skall upprättas i enlighet med det förfarande som fastställs i artikel 14 och omfattas av punkterna A, B och C i bilaga VI."
15. Artikel 5.9 ersätts med följande text och punkterna 10 och 11 läggs till:
"9. Beräkningen av de i punkterna 3 och 6 angivna procentandelarna utförs med tillämpning av reglerna i artiklarna 6 och 7 i direktiv 79/112/EEG.
10. En produkt som anges i artikel 1.1 får inte innehålla både en ingrediens som har erhållits i enlighet med reglerna i artikel 6 och samma ingrediens som har erhållits enligt andra regler.
11. Kommissionen skall före den 1 juli 1999 göra en förnyad granskning av bestämmelserna i denna artikel och artikel 10 och presentera lämpliga förslag för deras eventuella ändring."
16. Artikel 6 ersätts med följande text:
"Artikel 6
1. Ekologisk produktion innebär vid framställning av de produkter som anges i artikel 1.1 a med undantag för utsäde och vegetativt förökningsmaterial följande
a) åtminstone de bestämmelser som anges i bilaga I och, i förekommande fall, de tillämpningsförfaranden som hör till dessa skall vara uppfyllda,
b) endast produkter som består av ämnen som finns förtecknade i bilagorna I och II får användas som växtskyddsmedel, tvätt- och rengöringsmedel, gödningsmedel eller markberedningsmedel eller för varje annat ändamål som med avseende på vissa ämnen anges i bilaga II. De får endast användas på de särskilda villkor som anges i bilagorna I och II i den mån deras motsvarande användning är tillåten i vanligt jordbruk i de berörda medlemsländerna i enlighet med tillämpningen av gemenskapsbestämmelser eller enligt nationella bestämmelser som överensstämmer med gemenskapslagstiftningen,
c) endast utsäde och vegetativt förökningsmaterial som har producerats med den ekologiska produktionsmetod som anges i stycke 2 får användas.
2. För utsäde och vegetativt förökningsmaterial innebär den ekologiska produktionsmetoden att både moderplantan - såvitt avser utsäde - och föräldragenerationens planta/plantor - såvitt avser reproduktionsmaterial - har producerats i överensstämmelse med bestämmelserna i punkt 1 a och b under minst en generation eller, när det gäller perenna odlingar, minst två säsonger.
3. a) Trots vad som sägs i punkt 1 c får utsäde och vegetativt förökningsmaterial som inte har erhållits i enlighet med den ekologiska produktionsmetoden användas under en övergångsperiod fram till den 31 december 2000 med godkännande från den behöriga myndigheten i medlemsstaten under förutsättning att användarna av sådant förökningsmaterial på ett för medlemsstatens kontrollmyndighet eller kontrollorgan tillfredsställande sätt kan visa att de på gemenskapsmarknaden inte har kunnat erhålla ett förökningsmaterial för en lämplig sort av ifrågavarande art som uppfyller kraven i stycke 2. I detta fall skall ett förökningsmaterial som inte har behandlats med andra produkter än de som anges i bilaga II punkt B användas, under förutsättning att sådant material finns på gemenskapsmarknaden. Medlemsstaterna skall anmäla godkännanden som lämnats enligt detta stycke till de andra medlemsstaterna och till kommissionen,
b) förfarandet i artikel 14 kan användas för att fatta beslut om:
- införande, före den 31 december 2000, av begränsningar gällande den provisoriska åtgärd som anges i a i fråga om vissa arter och/eller typer av förökningsmaterial och/eller avsaknad av kemisk behandling,
- bibehållande, efter den 31 december 2000, av det i a angivna undantaget i fråga om vissa arter och/eller typer av förökningsmaterial för hela eller delar av gemenskapens område,
- införande av procedurregler och kriterier rörande det i a angivna undantaget och information om detta till berörda yrkesorganisationer, andra medlemsstater samt kommissionen.
4. Före den 31 december 1999, skall kommissionen göra en förnyad granskning av bestämmelserna i denna artikel, särskilt punkt 1 c samt punkt 2 och i förekommande fall presentera lämpliga förslag till ändring av dem."
17. Följande artikel införs efter artikel 6:
"Artikel 6a
1. I denna artikel anses med `plantor` hela plantor, avsedda för plantering för produktion av växter.
2. Den ekologiska produktionsmetoden innebär att plantor som används för produktion också skall ha producerats i enlighet med bestämmelserna i artikel 6.
3. Trots vad som sägs i punkt 2, får plantor som inte erhållits i överensstämmelse med den ekologiska produktionsmetoden användas under en övergångsperiod fram till den 31 december 1997 förutsatt att följande villkor är uppfyllda:
a) medlemsstatens behöriga myndighet har godkänt användning under förutsättning att användaren eller användarna av sådant material på ett tillfredsställande sätt kunnat visa medlemsstatens kontrollmyndighet eller kontrollorgan att de inte kunnat erhålla lämplig sort av ifrågavarande art på gemenskapsmarknaden,
b) plantorna har efter sådden inte behandlats med andra produkter än de som räknas upp i bilaga II, delarna A och B,
c) plantorna härstammar från en producent som har accepterat ett kontrollsystem som är likvärdigt med det system som avses i artikel 9 och som har accepterat att tillämpa förbehållet i punkt b. Denna bestämmelse träder i kraft den 1 januari 1996,
d) efter plantering skall plantorna ha odlats i enlighet med bestämmelserna i artikel 6.1 a och b under en period av minst sex veckor före skörden,
e) märkningen av produkter som innehåller ingredienser som härrör från sådana plantor får inte innehålla den uppgift som anges i artikel 10,
f) utan att detta påverkar någon inskränkning som följer av det i punkt 4 angivna förfarandet skall alla godkännanden som lämnats i enlighet med denna punkt återkallas när bristsituationen avhjälpts och de skall löpa ut senast den 31 december 1997.
4. a) När godkännanden som avses i punkt 3 har lämnats skall medlemsstaten omedelbart lämna följande upplysningar till övriga medlemsstater och kommissionen:
- datum för godkännandet,
- benämning för berörd sort och art,
- nödvändiga mängder samt skälen för detta,
- trolig varaktighet för bristsituationen,
- övriga upplysningar som begärts av kommissionen eller medlemsstaterna.
4. b) Om upplysningar, som av en medlemsstat lämnats till kommissionen och den medlemsstat som har lämnat godkännande, visar att en lämplig sort finns tillgänglig under den tid brist råder, får medlemsstaten återkalla ett godkännande eller förkorta dess giltighetstid. Medlemsstaten skall i sådant fall meddela kommissionen och de andra medlemsstaterna om de åtgärder den vidtagit senast inom tio dagar efter det att den mottagit upplysningarna.
4. c) På begäran av en medlemsstat eller på kommissionens initiativ, skall ärendet föreläggas den kommitté som avses i artikel 14. I enlighet med det förfarande som avses i artikel 14 kan beslut fattas om att återkalla eller förkorta godkännandets giltighetstid."
18. I artikel 7 skall följande stycke läggas till efter punkt 1:
"1a. De villkor som anges i punkt 1 gäller inte för produkter, som före antagandet av denna förordning allmänt användes i enlighet med vedertagna regler för ekologisk odling inom gemenskapen".
19. I artikel 9.1 skall orden "leverantörerna av produkter av det slag som anges i artikel 1" ersättas med orden "leverantörer som producerar, bereder eller från tredje land importerar produkter av det slag som anges i artikel 1."
20. I artikel 9.5 b ersätts ordet "avvikelser" med orden "avvikelser och/eller överträdelser".
21. I artikel 9.6 c ersätts ordet "överträdelser" med orden "avvikelser och/eller överträdelser".
22. I artikel 9.6 d ersätts orden "punkt 7-9" med orden "punkterna 7, 8, 9 och 11".
23. I artikel 9 införs följande punkt efter punkt 6:
"6a. Medlemsstaterna skall före den 1 januari 1996 tilldela varje kontrollorgan eller kontrollmyndighet som godkänts eller utsetts i enlighet med bestämmelserna i denna förordning ett kodnummer. De skall meddela övriga medlemsstater och kommissionen om detta och kommissionen skall offentliggöra kodnummer i den förteckning som anges i sista stycket i artikel 15."
24. Följande stycke skall införas i artikel 9:
"11. Utan att det påverkar tillämpningen av punkterna 5 och 6 skall de behöriga kontrollorganen från och med den 1 januari 1998 uppfylla kraven i EN 45011 av den 26 juni 1989."
25. Artikel 10.1 ersätts med följande text:
"1. Uppgift och/eller logotyp utvisande att produkterna omfattas av ett särskilt kontrollsystem som visas i bilaga V, får uteslutande ingå i märkningen av produkter av det slag som avses i artikel 1 när sådana produkter
a) överensstämmer med artikel 5.1 eller 5.3,
b) har varit underkastad den kontroll som avses i artikel 9 under hela produktions- och beredningsprocessen,
c) säljs direkt i slutna förpackningar av producent eller beredare till slutlig konsument, eller släpps ut på marknaden som färdigförpackade livsmedel. Vid direktförsäljning av producent eller beredare till slutlig konsument är slutna förpackningar inte nödvändiga när det av märkningen klart och tydligt framgår vilken produkt det är fråga om,
d) i märkningen är försedda med tillverkarens, beredarens eller säljarens namn på och/eller firma samt namn på eller kodnummer för kontrollmyndigheten eller kontrollorganet och övriga uppgifter som krävs i enlighet med reglerna för märkning av livsmedel som gäller i enlighet med gemenskapens lagstiftning."
26. I artikel 10.3 a ersätts orden "artikel 5-7" med orden "artiklarna 5 och 6".
27. Artikel 10.5, 10.6 och 10.7 ersätts med följande text:
"Allmänna åtgärder för verkställighet
Artikel 10a
1. När en medlemsstat med avseende på en produkt som härrör från en annan medlemsstat och som är försedd med de uppgifter som anges i artikel 2 och/eller bilaga V konstaterar avvikelser eller överträdelser rörande tillämpningen av denna förordning, skall den informera den medlemsstat som har utsett kontrollmyndigheten eller godkänt kontrollorganet och kommissionen om detta.
2. Medlemsstaterna skall vidta nödvändiga åtgärder för att undvika bedräglig användning av de uppgifter som anges i artikel 2 och/eller bilaga V."
28. I artikel 11.3 a ersätts orden "kontrollmyndigheterna" med orden "kontrollorgan och/eller kontrollmyndighet".
29. I artikel 11.6 a ersätts datumet den 31 juli 1995 med datumet den 31 december 2002.
30. I artikel 11.6 a ersätts den sista meningen med följande text:
"Den upphör från och med den tidpunkt då beslut att föra in ett tredje land i förteckningen som anges i punkt 1 a fattas, förutsatt att den inte rör en produkt som härrör från ett område som inte närmare preciseras i det beslut som anges i punkt 1 a och att den inte har granskats inom ramen för det tredje landets ansökan. Det tredje landet skall vara införstått med den fortsatta tillämpningsregeln av det förfarande för godkännande som anges i denna punkt."
31. I artikel 11 läggs följande punkt till:
"7. Kommissionen får på begäran av en medlemsstat i enlighet med det i artikel 14 angivna förfarandet godkänna ett tredje lands kontrollorgan, som den berörda medlemsstaten på förhand har utvärderat, och föra upp den på den förteckning som anges i punkt 1 a. Kommissionen skall underrätta det tredje landet om detta."
32. I artikel 13 införs följande strecksats före första strecksatsen:
"- tillämpningsföreskrifter för denna förordning."
33. I artikel 13 ersätts sista strecksatsen med följande strecksats:
"- de ändringar som skall göras i bilaga V för att fastlägga en logotyp för gemenskapen som kan användas tillsammans med eller i stället för uppgiften om att produkterna omfattas av ett särskilt kontrollsystem."
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter dess offentliggörande i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2694/95 av den 21 november 1995 om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 2588/95 (2), särskilt artikel 9 i denna, och med beaktande av följande:
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt motsvarande KN-nummer som anges i kolumn 2 med de motiveringar som ges i kolumn 3.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2802/95 av den 4 december 1995 om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 2588/95 (2), särskilt artikel 9 i denna, och med beaktande av följande:
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapens officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2805/95 av den 5 december 1995 om fastställande av exportbidrag inom vinsektorn och upphävande av förordning (EEG) nr 2137/93
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 822/87 av den 16 mars 1987 om den gemensamma organisationen av marknaden för vin (1), senast ändrad genom förordning (EG) nr 1544/95 (2), särskilt artikel 55.8 i denna, och
Förhållandena i den internationella handeln eller vissa marknaders särskilda krav kan göra det nödvändigt att differentiera bidraget med hänsyn till en bestämd produkts användning eller destination.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. De exportbidrag som avses i artikel 55 i förordning (EEG) nr 822/87 fastställs i bilagan till den här förordningen.
2. Förordning (EEG) nr 2137/93 skall upphöra att gälla.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2916/95 av den 18 december 1995 om ändring av vissa förordningar om den gemensamma organisationen av marknaderna för fjäderfäkött och ägg och om det gemensamma handelssystemet för äggalbumin och mjölkalbumin
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 234/79 av den 5 februari 1979 om förfarandet vid anpassning av Gemensamma tulltaxans nomenklatur för jordbruksprodukter (1), ändrad genom förordning (EEG) nr 3209/89 (2), särskilt artikel 2.1 i denna,
med beaktande av rådets förordning (EEG) nr 2771/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för ägg (3), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94 (4), särskilt artiklarna 3.2, 5.4, 6.4 och 18.13 i denna,
med beaktande av rådets förordning (EEG) nr 2777/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för fjäderfäkött (5), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94, särskilt artiklarna 5.4 och 8.12 i denna,
med beaktande av rådets förordning (EEG) nr 2783/75 av den 29 oktober 1975 om det gemensamma handelssystemet för äggalbumin och mjölkalbumin (6), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94, särskilt artiklarna 2.2, 3.4 och 4.4 i denna,
med beaktande av rådets förordning (EEG) nr 715/90 av den 5 mars 1990 om de bestämmelser som gäller för jordbruksprodukter och vissa varor som framställts genom förädling av jordbruksprodukter som har sitt ursprung i AVS-staterna eller i de utomeuropeiska länderna och territorierna (ULT) (7), senast ändrad genom förordning (EG) nr 2484/94 (8), särskilt artikel 27.2 i denna,
med beaktande av rådets förordning (EG) nr 3491/93 av den 13 december 1993 om vissa förfaranden vid tillämpning av Europaavtalen om upprättandet av en associering mellan Europeiska gemenskaperna och dess medlemsstater å ena sidan och Ungern, å andra sidan (9), senast ändrad genom förordning (EG) nr 3379/94 (10), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 3492/93 av den 13 december 1993 om vissa förfaranden för tillämpningen av Europaavtalet om upprättandet av en associering mellan Europeiska gemenskaperna och deras medlemsstater å ena sidan och Polen, å den andra sidan (11), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 3296/94 av den 19 december 1994 om vissa förfaranden för tillämpning av Europaavtalet om associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Tjeckien, å andra sidan (12), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 3297/94 av den 19 december 1994 om vissa förfaranden för tillämpning av Europaavtalet om associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Slovakien, å andra sidan (13), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EEG) nr 1601/92 av den 15 juni 1992 om särskilda åtgärder för Kanarieöarna rörande vissa jordbruksprodukter (14), senast ändrad genom kommissionens förordning (EG) nr 2537/95 (15), särskilt artikel 3.4 i denna,
med beaktande av rådets förordning (EG) nr 774/94 av den 29 mars 1994 om öppnande och förvaltning av vissa gemenskapstullkvoter för nötkött av hög kvalitet, griskött, fjäderfäkött, vete och blandsäd av vete och råg samt kli och andra restprodukter (16), senast ändrad genom kommissionens förordning (EG) nr 2198/95 (17), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 3641/93 av den 20 december 1993 om vissa förfaranden vid tillämpning av interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Bulgarien, å andra sidan (18), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 3642/93 av den 20 december 1993 om vissa förfaranden vid tillämpning av interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Rumänien, å andra sidan (19), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 1275/95 av den 29 maj 1995 om vissa förfaranden för tillämpningen av avtalet om frihandel och vissa handelsrelaterade frågor mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Estland, å andra sidan (20), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 1276/95 av den 29 maj 1995 om vissa förfaranden för tillämpningen av avtalet om frihandel och vissa handelsrelaterade frågor mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Lettland, å andra sidan (21), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 1277/95 av den 29 maj 1995 om vissa förfaranden för tillämpningen av avtalet om frihandel och vissa handelsrelaterade frågor mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Litauen, å andra sidan (22), särskilt artikel 1 i denna, och med beaktande av följande:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. KN-nummer 0207 31 skall ersättas med KN-nummer 0207 34. KN-nummer 0207 39 90 och 0207 50 skall ersättas med numren 0207 13 91, 0207 14 91, 0207 26 91, 0207 27 91, 0207 35 91, 0207 36 81, 0207 36 85 och 0207 36 89. Nummer 1602 32 skall införas efter nummer 1602 31
- i artikel 1.1 i förordning (EEG) nr 2777/75,
- i artikel 1 i kommissionens förordning (EEG) nr 109/80 (24).
2. KN-nummer 0105 12 skall införas före KN-nummer 0105 19
3. KN-nummer 1602 32 skall införas före KN-nummer 1602 39
- i artikel 6.2 i rådets förordning (EEG) nr 715/90,
- i artiklarna 1 och 3.1 b i kommissionens förordning (EEG) nr 903/90 (26).
4. KN-nummer 0207 23 skall ersättas med KN-nummer 0207 33 i bilaga I till kommissionens förordning (EEG) nr 1729/92 (27).
- kommissionens förordning (EEG) nr 2699/93 (28),
- kommissionens förordning (EG) nr 1431/94 (29),
- kommissionens förordning (EG) nr 1559/94 (30),
- kommissionens förordning (EG) nr 1474/95 (31),
- kommissionens förordning (EG) nr 1484/95 (32),
- kommissionens förordning (EG) nr 1866/95 (33).
6. Artikel 1 i rådets förordning (EEG) nr 2783/75 skall ersättas med följande:
"Artikel 1 Om inte annat föreskrivs i denna förordning skall Gemensamma tulltaxans tullsatser tillämpas för följande produkter:
>Plats för tabell>
Artikel 2
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 84.2 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
i enlighet med det i artikel 189c i fördraget angivna förfarandet (3), och
med beaktande av följande: Gemenskapen är allvarligt oroad över fartygsolyckor där människoliv går till spillo.
Internationella säkerhetsorganisationskoden för säker drift av fartyg och för förhindrande av förorening (hädanefter kallad "ISM-koden") antogs av Internationella sjöfartsorganisationen (IMO) genom församlingens resolution A.741(18) av den 4 november 1993 i medlemsstaternas närvaro och kommer, genom att den införlivas med 1974 års internationella konvention om säkerheten för människoliv till sjöss, att från och med den 1 juli 1998 tillämpas på ro-ro-passagerarfartyg.
Detta utgör en av en serie åtgärder för att förbättra säkerheten till sjöss. ISM-koden har ännu inte tvingande utan endast rekommenderande karaktär.
Människors säkerhet till sjöss kan förbättras avsevärt om ISM-koden tillämpas strikt och tvingande.
Den mest brådskande angelägenheten för gemenskapen utgörs av säkerhetsorganisationen på ro-ro-passagerarfartyg. Ett enhetligt och sammanhängande genomförande av ISM-koden i alla medlemsstater kan utgöra ett steg i riktning mot en säkerhetsorganisation för ro-ro-passagerarfartyg.
I sin resolution av den 22 december 1994 om säkerheten på ro-ro-passagerarfartyg (4) uppmanade rådet kommissionen att lägga fram ett förslag om ett påskyndat tvingande genomförande av ISM-koden för alla ro-ro-passagerarfartyg som bedriver reguljär trafik till eller från europeiska hamnar, i överensstämmelse med internationell rätt.
En strikt och tvingande tillämpning av ISM-koden är nödvändig för att säkerställa att säkerhetsorganisationssystem inrättas och bibehålls på vederbörligt sätt på både företags- och fartygsnivå av företag som bedriver havsgående trafik med ro-ro-passagerarfartyg.
Åtgärder på gemenskapsnivå är det bästa sättet att säkerställa ett påskyndat, tvingande genomförande av bestämmelserna i ISM-koden och en effektiv kontroll av tillämpningen av denna, samtidigt som en snedvridning av konkurrensen mellan olika gemenskapshamnar och ro-ro-passagerarfartyg undviks. Endast en förordning som är direkt tillämplig kan säkerställa ett sådant genomförande. För ett påskyndat genomförande krävs att förordningen tillämpas från och med den 1 juli 1996.
För det tvingande och påskyndade genomförandet av ISM-koden för alla ro-ro-passagerarfartyg, oavsett deras flagg, beaktas även anmodan enligt punkt 2 i IMO:s resolution A.741(18), vilken är en kraftfull uppmaning till regeringarna att införa ISM-koden snarast möjligt, i första hand för passagerarfartyg.
Fartygssäkerheten är flaggstaternas huvudansvar, och medlemsstaterna kan säkerställa att adekvata bestämmelser om säkerhetsorganisation följs av de fartyg som för deras flagg och de företag som bedriver trafik med dessa. Det enda sättet att garantera säkerheten på alla ro-ro-passagerarfartyg, oberoende av flagg, som bedriver eller önskar bedriva reguljär trafik från medlemsstaternas hamnar är att medlemsstaterna, som villkor för att bedriva reguljär trafik från deras hamnar, kräver att säkerhetsbestämmelserna verkligen följs.
Företag som endast bedriver trafik med ro-ro-passagerarfartyg i skyddade vatten mellan hamnar i samma medlemsstat utgör en mera begränsad risk och kommer att behöva utföra en proportionellt sett större mängd administrativt arbete än andra företag och bör därför beviljas ett temporärt undantag.
Det är nödvändigt att ange de krav som uppställs för att säkerställa genomförandet av ISM-koden och att definiera villkoren för utfärdande och kontroll av dokumentet om godkänd säkerhetsorganisation och av certifikatet om godkänd säkerhetsorganisation.
Medlemsstaterna kan komma att anse det nödvändigt att delegera eller att förlita sig på specialiserade organ för att uppfylla sina förpliktelser enligt denna förordning. Det lämpliga sättet att säkerställa en enhetlig och tillräcklig kontrollnivå är att kräva att dessa organ endast får vara sådana som uppfyller kraven i rådets direktiv 94/57/EG av den 22 november 1994 om gemensamma regler och standarder för organisationer som utför inspektioner och utövar tillsyn av fartyg och för sjöfartsadministrationernas verksamhet i förbindelse därmed (5).
En medlemsstat måste under förutsättning av att ett för medlemsstaterna bindande beslut fattas inom ramen för en föreskrivande kommitté ha rätt att tillfälligt dra in rätten att bedriva trafik med vissa ro-ro-passagerarfartyg från dess hamnar när den anser att det föreligger risk för allvarlig fara för säkerheten för liv eller egendom eller för miljön.
Ett förenklat förfarande som omfattar en kommitté med föreskrivande uppgifter är nödvändigt för att ändra denna förordning under beaktande av utvecklingen på internationell nivå.
Ett snabbt införande av dessa säkerhetsregler medför särskilda tekniska och administrativa problem för Grekland på grund av det mycket stora antal företag som är etablerade i Grekland och bedriver färjetrafik under grekisk flagg och uteslutande mellan grekiska hamnar. Ett undantag under begränsad tid för att hantera denna situation bör därför beviljas under beaktande även av att reguljär passagerar- och färjetrafik mellan grekiska hamnar fram till och med den 1 januari 2004 undantagits från tillämpningen av rådets förordning (EEG) nr 3577/92 av den 7 december 1992 om tillämpning av principen om frihet att tillhandahålla tjänster på sjötransportområdet inom medlemsstaterna (cabotage) (6).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syftet med denna förordning är att öka säkerheten vid ledning och drift av ro-ro-passagerarfartyg samt att förhindra förorening som orsakas av sådana fartyg i reguljär trafik till eller från hamnar i medlemsstater inom Europeiska gemenskapen, genom att säkerställa att företag som bedriver trafik med ro-ro-passagerarfartyg följer bestämmelserna i ISM-koden genom
- att företagen inrättar och på lämpligt vis upprätthåller ombordbaserade och landbaserade säkerhetsorganisationssystem, och
- att administrationerna i flagg- och hamnstaterna kontrollerar dessa.
Artikel 2
I denna förordning och för genomförandet av ISM-koden avses med
a) ro-ro-passagerarfartyg: ett havsgående passagerarfartyg som är utrustat med anordningar som gör det möjligt för väg- eller järnvägsfordon att rulla på och av fartyget, och som medför fler än 12 passagerare,
b) reguljär trafik: en serie av resor med ett ro-ro-passagerarfartyg som upprätthåller trafik mellan två eller flera platser, antingen
1. enligt en offentliggjord tidtabell, eller
2. med resor som företas så regelbundet eller så ofta att de utgör en uppenbar, systematisk serie.
c) företag: ro-ro-passagerarfartygets ägare eller någon annan organisation eller person, t.ex. redaren eller den som hyr fartyget utan besättning, som har övertagit fartygsägarens ansvar för ro-ro-passagerarfartygets drift.
d) erkänd organisation: ett organ som erkänts i enlighet med bestämmelserna i direktiv 94/57/EG.
e) ISM-koden: de internationella organisationsreglerna för säker drift av fartyg och för förhindrande av förorening, som antogs av IMO genom församlingens resolution A.741(18) av den 4 november 1993 och som utgör en bilaga till denna förordning,
f) administration: regeringen i den stat vars flagg ro-ro-passagerarfartyget har rätt att föra,
g) dokument om godkänd säkerhetsorganisation: det dokument som i enlighet med punkt 13.2 i ISM-koden utfärdas till företag,
h) certifikat om godkänd säkerhetsorganisation: det certifikat som i enlighet med punkt 13.4 i ISM-koden utfärdas till ro-ro-passagerarfartyg,
i) skyddade vatten: områden där sannolikheten per år för att det bildas vågor med en signifikant våghöjd över 1,5 m är mindre än 10 % och inom vilka ett ro-ro-passagerarfartyg aldrig befinner sig på större avstånd än 6 nautiska mil från en plats där fartyg kan söka skydd och där nödställda kan ta sig iland.
Artikel 3
Denna förordning skall tillämpas på alla företag som bedriver reguljär trafik med minst ett ro-ro-passagerarfartyg till eller från en hamn i en medlemsstat inom den Europeiska gemenskapen, oavsett fartygets flagg.
Artikel 4
1. Alla företag skall följa samtliga bestämmelser i punkterna 1.2 13.1 och 13.3 i ISM-koden, som om dessa bestämmelser vore tvingande, som ett villkor för att deras fartyg skall få bedriva reguljär trafik till eller från en hamn i en medlemsstat inom den Europeiska gemenskapen.
2. Utan hinder av bestämmelserna i punkt 1 får företag som bedriver reguljär trafik med ett eller flera ro-ro-passagerarfartyg enbart i skyddade vatten mellan hamnar som är belägna i en och samma medlemsstat uppskjuta efterlevnaden av bestämmelserna i denna förordning till den 1 juli 1997.
Artikel 5
1. Medlemsstaterna skall, med avseende på företag och ro-ro-passagerarfartyg, följa bestämmelserna i punkterna 13.2, 13.4 och 13.5 i ISM-koden som om dessa bestämmelser vore tvingande.
2. För tillämpningen av punkt 1 får medlemsstaterna endast godkänna, eller helt eller delvis förlita sig på, en erkänd organisation.
För tillämpningen av punkt 13.2 i ISM-koden får en medlemsstat endast utfärda dokument om godkänd säkerhetsorganisation för ett företag som har sin huvudsakliga verksamhetsort på dess eget territorium. Före ett sådant utfärdande skall medlemsstaterna samråda med administrationen i de stater vars flagg ifrågavarande företags ro-ro-passagerarfartyg har rätt att föra, om denna administration inte är den utfärdande medlemsstatens.
3. Dokumentet om godkänd säkerhetsorganisation skall endast gälla i fem år från dagen för dess utfärdande, under förutsättning att en kontroll görs en gång om året, för att bekräfta att säkerhetsorganisationssystemet fungerar väl, och att eventuella ändringar som gjorts sedan den senaste kontrollen uppfyller ISM-kodens bestämmelser.
4. Certifikatet om godkänd säkerhetsorganisation skall endast gälla i fem år från dagen för dess utfärdande, under förutsättning att en mellanliggande kontroll görs åtminstone var trettionde månad eller oftare för att bekräfta att säkerhetsorganisationssystemet fungerar väl och att eventuella ändringar som gjorts sedan den senaste kontrollen överensstämmer med ISM-kodens bestämmelser.
5. För tillämpningen av denna förordning och särskilt artikel 6 skall varje medlemsstat godkänna ett dokument om godkänd säkerhetsorganisation eller ett certifikat om godkänd säkerhetsorganisation som utfärdats av administrationen i någon annan medlemsstat eller av en erkänd organisation som handlar på dess vägnar.
6. En medlemsstat skall erkänna dokument om godkänd säkerhetsorganisation och certifikat om godkänd säkerhetsorganisation som utfärdats av administrationerna i tredje land, eller för dessas räkning, om det kan visas att de följer bestämmelserna i denna förordning.
Dokument om godkänd säkerhetsorganisation och certifikat om godkänd säkerhetsorganisation som utfärdats för administrationer i tredje land får endast erkännas om de har utfärdats av en erkänd organisation.
Artikel 6
Medlemsstaterna skall förvissa sig om att bestämmelserna i denna förordning följs av alla företag som bedriver reguljär färjetrafik med ro-ro-passagerarfartyg till eller från deras hamnar.
Artikel 7
Om en medlemsstat anser att ett företag, trots att det har ett dokument om godkänd säkerhetsorganisation, inte kan bedriva reguljär trafik med ett ro-ro-passagerarfartyg till eller från dess hamnar på grund av risk för allvarlig fara för säkerheten för liv eller egendom eller för miljön får rätten att bedriva denna trafik dras in tills faran har undanröjts.
Under ovannämnda förhållanden skall följande förfarande tillämpas:
Artikel 8
För att kunna beakta ISM-kodens allmänna begrepp skall kommissionen tre år efter denna förordnings ikraftträdande se över genomförandet av förordningen och föreslå lämpliga åtgärder.
Artikel 9
För att ta hänsyn till utvecklingen på det internationella planet och särskilt inom IMO får följande ändras, särskilt för att i bilagan införa riktlinjer för administrationer för genomförande av ISM-koden, i enlighet med förfarandet i artikel 10.2:
a) Definitionen av ISM-koden i artikel 2.
b) Giltighetstiden för dokumentet om godkänd säkerhetsorganisation och/eller certifikatet om godkänd säkerhetsorganisation och intervallen mellan kontrollerna av dem i artikel 5.3 och 5.4.
c) Bilagan.
Artikel 10
1. Kommissionen skall biträdas av den kommitté som inrättas enligt artikel 12.1 i rådets direktiv 93/75/EEG (7).
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag från kommissionen. Medlemsstaternas röster skall vägas enligt bestämmelserna i samma artikel. Ordföranden får inte rösta.
3. a) Kommissionen skall själv anta förslaget om det är förenligt med kommitténs yttrande.
b) Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
c) Om rådet inte har fattat något beslut vid utgången av en period på 40 dagar från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 11
Utan att det påverkar första stycket skall denna förordning inte tillämpas före den 31 december 1997 på företag som lyder under grekisk lag, har sin huvudsakliga verksamhetsort i Grekland och bedriver färjetrafik med ro-ro-passagerarfartyg som är registrerade i Grekland, för grekisk flagg och bedriver reguljär trafik endast mellan hamnar som är belägna i Grekland.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS BESLUT av den 25 juni 1996 om förbättring av gemenskapens jordbruksstatistik (96/411/EG)
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av rådets beslut 93/464/EEG av den 22 juli 1993 om ramprogram för prioriterade åtgärder för statistik information 1993 1997 (3), särskilt artikel 4 a i detta, och med beaktande av följande:
I ramprogrammet 1993 1997 som avses i beslut 93/464/EEG fastställs bland annat behovet av att bättre utnyttja de resurser som ägnas åt jordbruksstatistik genom genomförandet av resultaten av den "övervakningsverksamhet" som utfördes under det föregående statistiska programmet, som avses i rådets resolution av den 19 juni 1989 om genomförandet av en plan för prioriterade åtgärder för statistik: Europeiska gemenskapernas statistiska program (1989 1992) (4).
Genom denna övervakningsverksamhet har de viktigaste aspekterna på de förändringar av gemenskapens jordbruksstatistik som krävs fastställts.
Bland dessa förändringar återfinns de huvudområden där det är möjligt att göra besparingar och där det finns nya eller växande behov. Förändringarna bör vara i överensstämmelse med de överenskomna allmänna principerna.
Anpassningar på det nationella planet måste samordnas på gemenskapsnivå för att säkerställa att
a) uppgifterna fortsätter att vara tillräckligt tillförlitliga för varje medlemsstat och jämförbara medlemsstaterna emellan,
b) eventuella nödvändiga ändringar i rådets lagstiftning i god tid kan identifieras, förberedas och föreslås av kommissionen samt dessutom att kommissionen kan anta genomförandebestämmelser till rådets lagstiftning i god tid,
c) olika medlemsstaters metodologiska undersökningar om effektiva sätt att möta de nya informationsbehoven är lämpliga.
d) planeringen av nationella åtgärder tar tillbörlig hänsyn till det kollektiva gemenskapsintresset,
e) gemenskapens ekonomiska resurser till stöd för detta program utnyttjas så effektivt som möjligt som ett komplement till andra nationella resurser.
Denna samordning uppnås bäst genom att fastställa en formell struktur som gör det möjligt att gemensamt studera tekniska begränsningar och preferenser samt att fatta beslut som tar hänsyn både till gemenskapsintressen och nationella intressen.
Ett finansiellt bidrag till medlemsstaterna, i förhållande till deras objektiva behov, krävs för att underlätta nödvändiga anpassningar.
För att uppnå önskade besparingar kan det bli nödvändigt med anpassningar av det tekniska genomförandet av vissa undersökningar. Innan dessa anpassningar beviljas bör de undergå lämpliga säkerhetskontroller.
Nödvändiga åtgärder bör vidtas för en eventuell förlängning av detta beslut inom ramen för nästa ramprogram för prioriterade åtgärder för statistik avseende åren efter 1997.
Fördelningen av uppgifter mellan kommissionen och medlemsstaterna är helt i överensstämmelse med subsidiaritetsprincipen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte
För att jordbruksstatistiken bättre skall tillfredsställa det informationsbehov som reformen av den gemensamma jordbrukspolitiken leder till, skall medlemsstaterna, inom ramen för tillgängliga resurser, vidta lämpliga åtgärder för att anpassa sina nationella system för jordbruksstatistik. Medlemsstaterna skall härvidlag beakta de arbetsområden som anges i bilagorna I och II till detta beslut samt de mål, variabler och kriterier som anges i bilaga III.
Artikel 2
Kommissionens uppgift
Kommissionen skall i samråd med medlemsstaterna
a) fastställa en gemensam plan för samordning av arbetet och en allmän ram för nödvändiga metodologiska beskrivningar,
b) kontrollera uppgifternas kvalitet och jämförbarhet, samt
c) fastställa och genomföra åtgärder på gemenskapsnivå som är betydelsefulla för syftet med detta beslut.
Artikel 3
Tidsplan och förfarande
Den anpassningsprocess för gemenskapens jordbruksstatistik som avses i artikel 1 skall samordnas av kommissionen med hjälp av tekniska handlingsplaner i enlighet med vad som anges i artikel 4. Efter denna period kan rådet besluta om en förlängning i enlighet med kommissionens förslag i artikel 11.
Artikel 4
Tekniska handlingsplaner för jordbruksstatistiken
1. Kommissionen skall varje år fastställa en teknisk handlingsplan för jordbruksstatistiken i enlighet med förfarandet i artikel 10. Dessa planer skall omfatta de åtgärder som medlemsstaterna skall genomföra i enlighet med artikel 1. Disponibla resurser skall användas på ett sådant sätt att största möjliga förbättring av den gemensamma jordbruksstatistikens kostnadseffektivitet sker när kraven från gemenskapslagstiftningen, de informella avtalen och de nya informationsbehoven skall uppfyllas.
2. Varje årlig teknisk handlingsplan skall innehålla en detaljerad verksamhetsplan för det kommande året och en preliminär tidsplan för de två följande åren. Vid utarbetandet av denna tidsplan skall hänsyn tas till följande:
a) Befintliga åtaganden för åren i fråga, t.ex. en förteckning över de gemenskapsundersökningar som medlemsstaterna skall genomföra och frekvensen av dessa, samt andra uppgifter som skall lämnas till kommissionen.
b) Skriftlig information som medlemsstaterna skall lämna enligt artikel 5 b och 5 c.
c) Nödvändiga och tillgängliga resurser för alla planerade åtgärder.
Artikel 5
Medlemsstaternas rapporter
Medlemsstaterna skall senast den 31 mars varje år (år n) överlämna
a) en kort rapport om genomförandet av de åtgärder som beslutades för det föregående året (år ng 1),
b) en kortfattad beskrivning av de åtgärder som anges i planen för det kommande året (år n + 1),
c) information om viktiga, större åtgärder som planeras för eller avses genomföras under de två följande åren (åren n + 2 och n + 3) och som är av betydelse för syftet med detta beslut.
Beskrivningen skall omfatta de ändringar som anges avseende metodologin för genomförandet, arbeten som skall utföras, förutsedda svårigheter och förslag till lösningar på dem, konsekvenser för nationella och gemensamma resurser samt förslag till förbättringar på gemenskapsnivå. De åtgärder för vilka ekonomiskt gemenskapsstöd kommer att begäras skall anges.
I enlighet med det förfarande som anges i artikel 10 kommer kommissionen att utarbeta förenklade modeller för att underlätta utarbetandet av dessa rapporter.
Artikel 6
Finansiella bestämmelser
1. Kommissionen skall bidra till medlemsstaternas kostnader för att anpassa sina nationella system för jordbruksstatistik eller till kostnaderna för de förberedande arbeten som hänger samman med nya eller växande behov och som utgör en del av en teknisk handlingsplan.
2. Kommissionen skall varje år i samband med den tekniska handlingsplanen och i enlighet med förfarandet i artikel 10 fastställa beloppet för gemenskapsbidraget till varje medlemsstat.
3. Bidraget skall ges till medlemsstaterna årsvis efter det att de överlämnat den årliga rapporten om genomförandet av planerade åtgärder under det föregående året och den blivit godkänd av kommissionen. Kommissionen kan i samarbete med behöriga myndigheter i medlemsstaterna utföra alla kontrollåtgärder på plats som den anser nödvändiga.
Artikel 7
Flexibilitet
Då det med hänsyn till syftet med detta beslut är nödvändigt, kan kommissionen för en period som motsvarar en teknisk handlingsplan, i enlighet med förfarandet i artikel 10, godkänna en medlemsstats begäran om att anpassa en eller flera av följande undersökningskarakteristika i bilaga IV: undersökta regioner, territoriella underindelningar, definitioner, undersökningsmetodik, undersökningstidpunkt, variabellista och klassernas storlek.
Artikel 8
Anpassning till nya omständigheter
Kommissionen kan göra ändringar i bilaga I (statistiska områden där möjliga besparingar har fastställts) och i bilaga II (statistiska områden där det finns nya eller växande behov) i enlighet med förfarandet i artikel 10. Den skall informera Europaparlamentet och rådet om de ändringar som gjorts.
Artikel 9
Ständiga kommittén för jordbruksstatistik
Ständiga kommittén för jordbruksstatistik, som inrättades genom rådets beslut 77/279/EEG (5) skall sammanträda minst en gång om året för att diskutera följande:
a) Medlemsstaternas rapporter om genomförandet av åtgärderna under det föregående året.
b) De åtgärder som medlemsstaterna föreslår för det kommande året och utsikterna för de följande två åren.
c) Den tekniska handlingsplanen för det kommande året.
d) Gemenskapens finansiella bidrag enligt artikel 6.
e) Eventuella ändringar i bilagorna I och II.
Artikel 10
Nödvändiga åtgärder för tillämpningen
Kommissionen skall vidta de åtgärder som är nödvändiga för tillämpningen av detta beslut. Den skall biträdas av Ständiga kommittén för jordbruksstatistik, nedan kallad "kommittén".
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittéen skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen, varvid medlemsstaternas röster skall vägas enligt samma artikel. Ordföranden får inte rösta.
Kommissionen skall själv anta de föreslagna åtgärderna om de är förenliga med kommitténs yttrande.
Om de föreslagna åtgärderna inte är förenliga med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall besluta med kvalificerad majoritet.
Om rådet inte har beslutat inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 11
Rapport
Senast den 1 november 1997 och efter samråd med Ständiga kommittén för jordbruksstatistik skall kommissionen till Europaparlamentet och rådet överlämna en rapport om genomförandet av detta beslut, vid behov åtföljd av förslag till dess förlängning.
Artikel 12
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 20 maj 1996 om utsläppande på marknaden av en genetiskt modifierad hansteril cikoria med partiell tolerans mot herbiciden glufosinatammonium (Cichorium intybus L.) enligt rådets direktiv 90/220/EEG (Text av betydelse för EES) (96/424/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/220/EEG av den 23 april 1990 om avsiktlig utsättning av genetiskt modifierade organismer i miljön (1), ändrat genom kommissionens direktiv 94/15/EG (2), särskilt artikel 13 i detta, och med beaktande av följande:
I artikel 10 till 18 i direktiv 90/220/EEG fastställs ett gemenskapsförfarande som bemyndigar en medlemsstats behöriga myndighet att medge utsläppande på marknaden av levande produkter som består av genetiskt modifierade organismer.
En anmälan om utsläppande på marknaden av en sådan produkt har inlämnats till den behöriga myndigheten i en medlemsstat (Nederländerna).
Nederländernas behöriga myndighet har överlämnat handlingarna i ärendet till kommissionen med tillstyrkan. De behöriga myndigheterna i andra medlemsstater har rest invändningar mot handlingarna.
Enligt artikel 13.3 skall kommissionen därför besluta enligt förfarandet i artikel 21 i direktiv 90/220/EEG.
Efter att ha granskat de handlingar som inlämnats enligt direktiv 90/220/EEG och beaktat all den information som överlämnats av medlemsstaterna har kommissionen kommit fram till följande slutsatser:
- Det finns ingen anledning att tro att det skulle uppstå negativa inverkningar genom en överföring av bar-genen till vilda cikoriapopulationer; eftersom en sådan överföring endast skulle utgöra en konkurrensmässig eller selektiv fördel gentemot vilda populationer om herbiciden glufosinatammonium vore den enda faktorn som begränsade dessa populationer, vilket inte är fallet.
- Tillstånd till utsläppande på marknaden av denna produkt bör inte omfatta dess användning som livsmedel eller djurfoder, eftersom den anmälan som ingått omfattar dessa aspekter.
- Det föreligger inga säkerhetsskäl för att på etiketten ange att produkten erhållits genom genetisk förändring.
- Eftersom 50 % av det hybrida utsädet är tolerant mot herbiciden i fråga, bör etiketten ange att produkten kan vara tolerant mot herbiciden glufosinatammonium, så att odlarna är medvetna om att det eventuellt inte är möjligt att kontrollera oönskade groddar av produkter med glufosinatammonium.
Tillstånd för användning av kemiska herbicider på växter, samt utvärderingen av deras inverkan på människors hälsa och på miljön är underkastade rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande på marknaden av växtskyddsprodukter (3), senast ändrat genom kommissionens direktiv 96/12/EG (4), och faller därför inte under tillämpningsområdet för direktiv 90/220/EEG.
Artiklarna 11.6 och 16.1 i direktivet ger ytterligare skydd om ny kunskap om risker förknippade med produkten blir tillgänglig.
Detta beslut är förenligt med yttrandet från den kommitté bestående av företrädare för medlemsstaterna som inrättas enligt artikel 21 i direktiv 90/220/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Utan att det påverkar gemenskapslagstiftningen, och i överensstämmelse med de villkor som fastställs i styckena 2, 3 och 4, skall tillstånd för utsläppande på marknaden ges av de nederländska myndigheterna för följande produkt anmäld av Bejo-Zaden BV (ref. C/NL/94/25) i enlighet med artikel 13 i direktiv 90/220/EEG.
Produkten består av frön och plantor från cikorialinjerna Cichorium intybus L. subspecies radicchio rosso (RM3-3, RM3-4 och RM3-6) som framställts med hjälp av Agrobacterium tumefaciens-modifierad Ti-plasmid och som innehåller följande inom T-DNA-gränserna:
i) Barnase-genen från Bacillus amyloliquefaciens (ribonukleas) med promotorn PTA29 från Nicotiana tabaccum och terminatorn från nopalinsyntasgenen från Agrobacterium tumefaciens.
ii) Bar-genen från Streptomyces hygroscopicus (fosfinotricinacetyltransferas) med promotorn PSsuAra-tp från Arabidopsis thaliana och TL-DNA-gen-7-promotorn från Agrobacterium tumefaciens.
iii) Neo-genen från Escherichia coli (neomycinfosfotransferas II) med promotorn från nopalinsyntasgenen från Agrobacterium tumefaciens och octopinsyntasgenterminatorn från Agrobacterium tumefaciens.
2. Medgivandet avser utsäde av alla hybrider mellan denna produkt och icke genetiskt modifierad cikoria.
3. Medgivandet avser användning av produkten för odlingsverksamhet.
4. Utan att det påverkar bestämmelserna om etikettering och märkning i övrig gemenskapslagstiftning skall det på etiketten till varje utsädesförpackning anges att produkten
- skall användas för odlingsverksamhet.
- och kan vara tolerant mot herbiciden glufosinatammonium.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 28 juni 1996 om särskilda importvillkor för fiskeri- och vattenbruksprodukter med ursprung i Mauretanien (Text av betydelse för EES) (96/425/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av fiskeriprodukter (1), senast ändrat genom direktiv 95/71/EG (2) uppfylls, särskilt artikel 11 i detta, och med beaktande av följande:
En expertdelegation utsänd av kommissionen har kommit tillbaka från Mauretanien efter att ha förvissat sig om villkoren för produktion, lagring och transport av fiskeriprodukter med gemenskapen som destination.
Föreskrifterna i den mauretanska lagstiftningen i fråga om inspektion om hygienkontroll av fiskeriprodukter kan betraktas som likvärdiga med dem som fastställs genom direktiv 91/493/EEG.
"Ministère des Pêches et de l'Économie Maritime - Centre National de Recherches Océanographiques et des Pêches - Département Valorisation et Inspection Sanitaire (MPEM - CNROP - DVIS)" kan på ett effektivt sätt granska tillämpningen av den gällande lagstiftningen.
Villkoren för det intyg som avses i artikel 11.4 a i direktiv 91/493/EEG omfattar fastställande av en mall för intyget, vilket eller vilka språk intyget skall vara avfattat på och vilken ställning den som undertecknar intyget skall ha.
Det är lämpligt att i enlighet med artikel 11.4 b i direktiv 91/493/EEG anbringa ett märke med uppgifter om det tredje landets namn och ursprungsanläggningens eller frysfartygets godkännandenummer på förpackningen för fiskeriprodukterna.
I enlighet med artikel 11.4 c i direktiv 91/493/EEG är det viktigt att fastställa en förteckning över godkända anläggningar eller frysfartyg. Denna förteckning bör fastställas på grundval av ett meddelande från MPEM - CNROP - DVIS till kommissionen. Det åligger alltså MPEM - CNROP - DVIS att försäkra sig om att de åtgärder som föreskrivs i detta syfte i artikel 11.4 i direktiv 91/493/EEG efterlevs.
MPEM - CNROP - DVIS har officiellt gett försäkringar i fråga om efterlevnaden av de regler som anges i kapitel V i bilagan till direktiv 91/493/EEG och i fråga om krav som är likvärdiga med dem som föreskrivs i det direktivet för godkännande av anläggningar och frysfartyg.
De åtgärder om föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Det intyg som avses i artikel 2.1 skall utfärdas på minst ett av de officiella språken i den medlemsstat där kontrollen äger rum.
2. I intyget skall finnas namn och tjänstebeteckning på representanten för "Ministère des Pêches et de l'Économie Maritime - Centre National de Recherches Océanographiques et des Pêches - Département Valorisation et Inspection Sanitaire (MPEM - CNROP - DVIS)", dennes namnteckning samt den officiella stämpeln för MPEM - CNROP - DVIS; allt detta skall vara i en annan färg än övriga uppgifter i intyget.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 14 oktober 1996 om särskilda importvillkor för fiskeri- och vattenbruksprodukter med ursprung i Elfenbenskusten (Text av betydelse för EES) (96/609/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av fiskeriprodukter (1), senast ändrat genom direktiv 95/71/EG (2), särskilt artikel 11 i detta, och med beaktande av följande:
En expertdelegation utsänd av kommissionen har kommit tillbaka från Elfenbenskusten efter att ha förvissat sig om villkoren för produktion, lagring och transport av fiskeriprodukter med gemenskapen som destination.
Föreskrifterna i Elfenbenskustens lagstiftning i fråga om inspektion och hygienkontroll av fiskeriprodukter kan betraktas som likvärdiga med dem som fastställs genom direktiv 91/493/EEG.
"Ministère de l'agriculture et des ressources animales - Direction générale des ressources animales (MARA-DGRA)" kan på ett effektivt sätt granska tillämpningen av den gällande lagstiftningen.
Villkoren för det intyg som avses i artikel 11.4 a i direktiv 91/493/EEG omfattar fastställande av en mall för intyget, vilket eller vilka språk intyget skall vara avfattat på och vilken ställning den som undertecknar intyget skall ha.
Det är lämpligt att i enlighet med artikel 11.4 b i direktiv 91/493/EEG anbringa ett märke med uppgifter om det tredje landets namn och ursprungsanläggningens godkännandenummer på förpackningen för fiskeriprodukterna.
I enlighet med artikel 11.4 c i direktiv 91/493/EEG är det viktigt att fastställa en förteckning över godkända anläggningar. Denna förteckning bör fastställas på grundval av ett meddelande från Ministère de l'agriculture et des ressources animales - Direction générale des ressources animales (MARA-DGRA) till kommissionen. Det åligger alltså MARA-DGRA att försäkra sig om att de åtgärder som föreskrivs i detta syfte i artikel 11.4 i direktiv 91/493/EEG efterlevs.
MARA-DGRA har officiellt gett försäkringar i fråga om efterlevnaden av de regler som anges i kapitel V i bilagan till direktiv 91/493/EEG och i fråga om krav som är likvärdiga med dem som föreskrivs i det direktivet för godkännande av anläggningar.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Det intyg som avses i artikel 2.1 skall utfärdas på minst ett av de officiella språken i den medlemsstat där kontrollen äger rum.
2. I intyget skall finnas namn och tjänstebeteckning på representanten för MARA-DGRA, dennes namnteckning samt den officiella stämpeln för MARA-DGRA; allt detta skall vara i en annan färg än övriga uppgifter i intyget.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
RÅDETS DIREKTIV 96/22/EG av den 29 april 1996 om förbud mot användning av vissa ämnen med hormonell och tyreostatisk verkan samt av â-agonister vid animalieproduktion och om upphävande av direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande Ekonomiska och sociala kommitténs yttrande (3), och
med beaktande av följande: 1. Genom rådets direktiv 81/602/EEG (4) förbjöds vissa ämnen med hormonell eller tyreostatisk verkan och genom direktiv 88/146/EEG (5) förbjöds användningen av vissa ämnen med hormonell verkan i animalieproduktion men tilläts samtidigt vissa undantag.
2. I rådets direktiv 88/299/EEG (6) fastställs villkor för undantag från förbudet att handla med vissa djurkategorier som anges i artikel 7 i direktiv 88/146/EEG, samt kött från dessa.
3. Vissa substanser med tyreostatisk, östrogen, androgen eller gestagen verkan kan, p.g.a. de restsubstanser de ger i kött och andra livsmedel av animaliskt ursprung, vara farliga för konsumenterna och de kan även påverka kvalitén i livsmedel av animaliskt ursprung.
4. Nya ämnen med anabol verkan såsom â-agonister används illegalt vid uppfödning i syfte att stimulera djurens tillväxt och produktivitet.
5. Resultaten från den undersökning som genomfördes av kommissionen 1990 till 1992 i medlemsstaterna visar på stor tillgång av â-agonister i animalieproduktionen vilket gynnar illegal användning.
6. Olämplig användning av â-agonister kan innebära allvarlig fara för människors hälsa. För konsumenternas skull bör innehav av â-agonister liksom tillförsel till alla slags djur samt avyttring för detta syfte förbjudas. Innehav av stilbener och tyreostatiska medel liksom tillförsel till alla slags djur och avyttring bör också förbjudas. Användningen av andra ämnen bör regleras.
7. Tillförsel av läkemedel baserade på â-agonister kan emellertid tillåtas i noggrant definierade terapeutiska syften för vissa kategorier nötkreatur, hästdjur och sällskapsdjur.
8. Det är dessutom nödvändigt att garantera alla konsumenter samma villkor vid anskaffande av kött och livsmedel från kött, samt att erbjuda dem en produkt som motsvarar deras förväntningar. Med tanke på konsumenternas mottaglighet kan möjligheterna att få avsättning för produkterna i fråga härigenom enbart öka.
9. Det är lämpligt att behålla förbudet mot hormonella ämnen i tillväxtbefrämjande syfte. Om tillförsel av vissa ämnen kan tillåtas i terapeutiskt eller zootekniskt syfte skall den noggrant kontrolleras för att undvika varje form av felaktig användning.
10. Bristande harmonisering på gemenskapsnivå beträffande karenstid och de stora skillnader som föreligger mellan medlemsstater, särskilt beträffande godkända veterinärmedicinska läkemedel som innehåller hormonella substanser eller â-agonister, gör att maximala karenstider för dessa läkemedel i harmoniseringssyfte bör bestämmas.
11. Levande djur som behandlas på detta sätt i terapeutiskt eller zootekniskt syfte och kött från dessa djur kan i princip inte bli föremål för handel med tanke på den inverkan det skulle ha på en effektiv kontroll av systemet. Undantag från detta förbud kan emellertid göras under vissa villkor beträffande handel inom gemenskapen och import från tredje land av djur avsedda för avel samt av uttjänta avelsdjur.
12. Undantag kan tillåtas om tillräckliga garantier ges för att förebygga obalans i handeln. Dessa garantier bör gälla produkter som kan användas, villkor för deras användning och kontroll av dessa villkor, särskilt när det gäller att respektera den nödvändiga karenstiden.
13. Effektiv kontroll av tillämpningen av bestämmelserna i detta direktiv bör säkerställas.
14. Direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG bör upphävas.
15. För att illegal användning av tillväxtbefrämjande och produktivitetshöjande medel i animalieproduktion skall kunna bekämpas effektivt i alla medlemsstater bör de åtgärder som skall vidtas organiseras på gemenskapsnivå.
16. Den 18 januari 1996 uppmanades kommissionen och rådet av Europaparlamentet att fortsätta att motsätta sig import av hormonbehandlat kött till gemenskapen; parlamentet önskade att totalförbudet mot användning av tillväxtbefrämjande medel i uppfödningen skulle kvarstå och uppmanade i detta syfte rådet att snarast anta kommissionens förslag om vilket parlamentet yttrat sig den 19 april 1994.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. I detta direktiv tillämpas de definitioner för kött och köttprodukter som återfinns i direktiv 64/433/EEG (7), 71/118/EEG (8), 77/99/EEG (9), 91/495/EEG (10) för vattenbruksprodukter som återfinns i direktiv 91/493/EEG (11), samt de definitioner för veterinärmedicinska läkemedel som återfinns i direktiv 81/851/EEG (12) och 81/852/EEG (13).
2. Dessutom avses med
a) husdjur: tama djur av arterna nötkreatur, svin, får getter, hovdjur, fjäderfä och kaniner, samt vilda djur av dessa arter och vilda idisslare, uppfödda i hägn,
b) terapeutisk behandling: tillförsel av godkända ämnen genom tillämpning av artikel 4 i det här direktivet, till ett enstaka husdjur i syfte att, efter undersökning av en veterinär, behandla fertilitetsstörningar inklusive avbrytande av oönskad dräktighet och när det gäller â-agonister, för att motverka livmoderkontraktioner hos kor vid kalvning samt behandla andningssvårigheter och motverka livmoderkontraktioner hos hästdjur som uppfötts av andra skäl än för köttproduktion,
c) zooteknisk behandling:
i) tillförsel till enstaka husdjur av ett av de ämnen som tillåts enligt artikel 5 i detta direktiv, i syfte att synkronisera östrus och förbereda donatorer och recipienter vid implantation av embryon, efter det att djuret undersökts av veterinär eller enligt artikel 5, stycke 2, på dennes ansvar,
ii) till vattenbruksdjur, till en avelsgrupp i syfte att erhålla inverterat kön, efter förskrivning av veterinär och på dennes ansvar,
d) illegal behandling: användning av icke godkända ämnen eller produkter eller användning av enligt gemenskapslagstiftningen godkända ämnen eller produkter för andra ändamål eller på andra villkor än vad som föreskrivs i gemenskapslagstiftningen eller - i förekommande fall - i de olika nationella lagstiftningarna.
Artikel 3
Medlemsstaterna skall säkerställa att följande förbjuds:
a) Tillförsel av ämnen med tyreostatisk, östrogen, androgen eller gestagen verkan, samt â-agonister till ett husdjur eller vattenbruksdjur, oavsett på vilket sätt det sker.
b) Innehav av djur som avses i a i ett jordbruksföretag, utom under officiell kontroll samt avyttring eller slakt, som livsmedel, av husdjur eller vattenbruksdjur som innehåller ämnen som avses i a eller i vilka förekomsten av sådana ämnen har konstaterats, utom i det fall det kan bevisas att dessa djur har behandlats enligt artikel 4 eller 5.
c) Avyttring av vattenbruksdjur, som livsmedel, om djuren tillförts ämnen som avses i a, samt bearbetade produkter av dessa djur.
d) Avyttring av kött från djur som avses i b.
e) Bearbetning av kött som avses i d.
Artikel 4
Trots artikel 2 och 3, får medlemsstaterna tillåta följande:
1. Tillförsel till husdjur i terapeutiskt syfte av östradiol 17 â, testosteron, progesteron eller derivat som efter resorption på platsen för applicering vid hydrolys bildar den ursprungliga komponenten. Veterinärmedicinska läkemedel som används för terapeutisk behandling skall uppfylla föreskrifterna för avyttring enligt direktiv 81/851/EEG och kan tillföras endast av veterinär på husdjur som noggrant identifierats och i form av injektion eller för behandling av äggstocksrubbningar i form av vaginalspiral, men inte i form av implantat. Behandling av identifierade djur skall registreras av den ansvarige veterinären. Denne skall i ett register, som kan vara det som föreskrivs i direktiv 81/851/EEG, anteckna minst följande upplysningar:
- slag av behandling,
- slag av godkända produkter,
- behandlingsdatum,
- behandlade djurs identititet.
Detta register skall på begäran ställas till behörig myndighets förfogande.
2. Tillförsel i terapeutiskt syfte av registrerat veterinärmedicinskt läkemedel som innehåller
i) trenbolon allyl som skall intas oralt eller â-agonister till hästdjur eller sällskapsdjur under förutsättning att de används enligt tillverkarens specifikationer,
ii) â-agonister i form av injektion för att motverka livmoderkontraktioner hos kor i samband med kalvning.
Tillförseln skall utföras av veterinär eller, vad beträffar veterinärmedicinska läkemedel enligt i, på dennes direkta ansvar; behandlingen skall registreras av den ansvarige veterinären, och minst de upplysningar som anges i punkt 1 skall anges.
Innehav av veterinärmedicinska läkemedel som innehåller â-agonister vilka kan användas för att motverka livmoderkontraktioner är förbjuden.
Utan att det påverkar tillämpningen av första stycket i punkt 2 ii är emellertid terapeutisk behandling förbjuden för produktionsdjur, inklusive uttjänta avelsdjur.
Artikel 5
Trots artikel 3 a och utan att det påverkar tillämpningen av artikel 2, kan medlemsstaterna i zootekniskt syfte tillåta tillförsel till husdjur av veterinärmedicinska läkemedel med östrogen, androgen eller gestagen verkan, godkända enligt direktiv 81/851/EEG och 81/852/EEG. Tillförseln skall utföras av en veterinär till noggrant identifierade djur och behandlingen skall registreras av den ansvarige veterinären enligt artikel 4.1.
Medlemsstaterna kan emellertid tillåta att synkronisering av östrus samt förberedelser av donatorer och recipienter för implantation av embryon inte utförs av veterinär utan endast på dennes ansvar.
När det gäller vattenbruksdjur kan fiskyngel behandlas med veterinärmedicinska läkemedel med androgen verkan under de tre första månaderna för att erhålla inverterat kön; medicinerna skall vara godkända enligt direktiv 81/851/EEG och 81/852/EEG.
I de fall som avses i denna artikel, skall veterinären utfärda ett recept som inte kan förnyas, i vilket den aktuella behandlingen skall specificeras och nödvändig mängd av produkten anges, och veterinären skall också registrera förskrivna produkter.
Behandling i zootekniskt syfte är emellertid förbjuden på produktionsdjur, inklusive under gödningsperiod för uttjänta avelsdjur.
Artikel 6
1. Hormonprodukter och â-agonister vars tillförsel till husdjur enligt artikel 4 och 5 är tillåten, skall motsvara kraven i direktiv 81/851/EEG och 81/852/EEG.
2. Följande kan emellertid inte tillåtas enligt punkt 1:
a) Nedanstående hormonprodukter:
i) Produkter med depåeffekt.
ii) Produkter där karenstiden är längre än 15 dygn efter behandling.
iii) Produkter
- som är godkända enligt de bestämmelser som var i kraft före ändringen genom förordning (EEG) nr 2309/93 (14),
- med okända användningsvillkor,
- för vilka det inte finns någon reagens eller utrustning som krävs till analysmetoder för att upptäcka förekomst av restsubstanser som överstiger de tillåtna gränserna.
b) Veterinärmedicinska läkemedel som innehåller â-agonister med en karenstid som överstiger 28 dygn efter avslutad behandling.
Artikel 7
1. I handelssyfte kan medlemsstaterna tillåta avyttring av djur avsedda för avel, eller uttjänta avelsdjur, som under sin aktiva period varit föremål för någon av behandlingarna enligt artikel 4 och 5, samt tillåta anbringande av gemenskapens kontrollmärke på kött från sådana djur, om villkoren i artikel 4 och 5 och om minimal karenstid enligt artikel 6.2 a ii eller b eller karenstiden som avses i avyttringstillståndet respekterats.
Handel med hästar med högt värde, särskilt kapplöpningshästar, tävlingshästar, cirkushästar eller hästar avsedda för betäckning eller utställning, inklusive registrerade hästdjur som tillförts veterinärmedicinska läkemedel innehållande trenbolon allyl eller â-agonister i de syften som anges i artikel 4, kan emellertid äga rum innan karenstiden är över, under förutsättning att villkoren för tillförsel har uppfyllts och att slag av behandling samt datum för behandling anges på det intyg eller pass som följer med dessa djur.
2. Kött eller produkter från djur som tillförts ämnen med östrogen, androgen eller gestagen verkan eller â-agonister kan enligt reglerna om undantag från detta direktiv avyttras för konsumtion endast om djuren i fråga har behandlats med veterinärmedicinska läkemedel som uppfyller kraven i artikel 6, och under förutsättning att den föreskrivna karenstiden har iakttagits innan djuren slaktas.
Artikel 8
Medlemsstaterna skall säkerställa följande:
1) Att innehav av ämnen som avses i artikel 2 och artikel 3 a begränsas till personer som har tillstånd enligt nationell lagstiftning i enlighet med artikel 1 i direktiv 90/676/EEG (15), vid import, tillverkning, lagring, distribution, försäljning eller användning.
2) Att utöver de kontroller som föreskrivs i direktiv om avyttring av olika produkter i fråga, de officiella kontrollerna enligt artikel 11 i direktiv 96/23/EG (16) genomförs av behöriga nationella myndigheter utan förvarning i syfte att konstatera
a) om förbjudna ämnen eller produkter som är avsedda för tillförsel till djur i tillväxtbefrämjande syfte enligt artikel 2 innehas eller förekommer,
b) om djur behandlas illegalt,
c) om karenstider enligt artikel 6 respekteras,
d) om restriktionerna i artikel 4 och 5 för användning av vissa substanser eller produkter respekteras.
3) Att sökande efter
a) förekomst av ämnen som avses under punkt 1 i djur eller djurens dricksvatten, samt på samtliga platser där djuruppfödning eller djurhållning äger rum,
4) Att när kontrollerna enligt punkt 2 och 3
a) visar på förekomst av ämnen eller produkter där användning eller innehav är förbjudet eller förekomsten av restsubstanser från ämnen vars tillförsel inneburit illegal behandling, skall dessa ämnen eller produkter beslagtas medan djur som eventuellt behandlats, eller deras kött, placeras under officiell kontroll till dess att nödvändiga påföljder genomförts,
b) visar att kraven under punkt 2 b och 2 c inte iakttagits, skall den behöriga myndigheten vidta lämpliga åtgärder, i proportion till överträdelsens omfattning.
Artikel 9
Utan att det påverkar tillämpningen av direktiv 81/851/EEG skall företag som köper eller tillverkar ämnen med tyreostatisk, östrogen, androgen eller gestagen verkan eller â-agonister och de företag som har något slag av tillstånd för att utöva handel med nämnda substanser, samt de företag som köper eller producerar farmaceutiska produkter och veterinärmedicinska läkemedel utifrån dessa ämnen, upprätta ett register i kronologisk ordning över tillverkade eller införskaffade produkter och dem som överlåtits eller används för tillverkning av läkemedelspreparat och veterinärmedicinska läkemedel och till vem dessa har överlåtits eller sålts.
Upplysningarna som avses i första stycket skall på begäran ställas till behörig myndighets förfogande, och om de föreligger i elektronisk form, även som papperskopia.
Artikel 10
När resultaten av de kontroller som utförts i en medlemsstat visar att kraven i detta direktiv inte iakttagits i djurens eller produkternas ursprungsland, skall den behöriga myndigheten i den medlemsstaten tillämpa reglerna i rådets direktiv 89/608/EEG av den 21 november 1989 beträffande ömsesidigt stöd mellan medlemsstaternas administrativa myndigheter, samt samarbetet mellan dessa och kommissionen, i syfte att garantera att lagstiftningen på det veterinära och zootekniska området tillämpas korrekt (17).
Artikel 11
1. Tredje länder vilkas lagstiftning tillåter avyttring och tillförsel av stilbener, stilbenderivat, deras salter eller estrar samt tyreostatiska medel i syfte att tillföra dem till alla djurarter, får inte finnas på någon lista som enligt gemenskapslagstiftningen reglerar från vilka länder medlemsländerna har tillstånd att importera husdjur eller vattenbruksdjur eller kött eller produkter från sådana djur.
2. Medlemsstaterna skall dessutom säkerställa att import från tredje land som förekommer på en av de listor som avses i punkt 1 förbjuds
a) av husdjur eller vattenbruksdjur
i) som på något sätt tillförts produkter eller ämnen som avses i artikel 2 a,
ii) som tillförts de ämnen eller produkter som avses i artikel 3 a, utom om tillförseln sker enligt bestämmelser och krav i artikel 4, 5 och 7 i detta direktiv och om den karenstid som tillåts i de internationella rekommendationerna iakttagits,
b) av kött eller produkter från djur som enligt punkt a ej får importeras.
3. Djur avsedda för avel, uttjänta avelsdjur, eller deras kött, vilka härrör från tredje land, får emellertid importeras under förutsättning att de uppfyller garantier som minst motsvarar dem som anges i detta direktiv och som inrättats enligt förfarandet i artikel 33 i rådets direktiv 96/23/EG, och med tillämpning av kapitel V i det direktivet.
4. Kontroller beträffande import från tredje land skall utföras enligt föreskrifterna i artikel 4.2 c i rådets direktiv 91/496/EEG av den 15 juli 1991 om fastställande av regler för hur veterinärkontroller skall organiseras för djur som importeras till gemenskapen från tredje land (18) och som enligt artikel 8.2 i rådets direktiv 90/675/EEG av den 10 december 1990 om principerna för organisering av veterinärkontroller av produkter som förs in i gemenskapen (19) från tredje land.
Artikel 12
Rådet får, på förslag av kommissionen och med kvalificerad majoritet, anta nödvändiga övergångsåtgärder innan den ordning som föreskrivs i detta direktiv trätt i kraft.
Artikel 13
1. Direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG skall upphöra att gälla den 1 juli 1997.
2. Hänvisningar till de upphävda direktiven skall läsas som hänvisningar till detta direktiv och skall läsas enligt jämförelsetabellen i bilagan.
Artikel 14
1. Medlemsstaterna skall anta de lagar och andra författningar, i förekommande fall med påföljder, som är nödvändiga för att följa detta direktiv den 1 juli 1997 och vad beträffar â-agonister, senast den 1 juli 1997. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter för hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
3. Innan bestämmelserna i detta direktiv avseende â-agonister genomförs, skall de nationella reglerna på området vara tillämpliga, varvid allmänna bestämmelser i fördraget skall iakttas.
Artikel 15
KOMMISSIONENS DIREKTIV 96/28/EG av den 10 maj 1996 om anpassning till teknisk utveckling av rådets direktiv 76/116/EEG om tillnärmning av medlemsstaternas lagstiftning om gödselmedel (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av rådets direktiv 76/116/EEG av den 18 december 1975 om tillnärmning av medlemsstaternas lagstiftning om gödselmedel (1), senast ändrat genom direktiv 89/530/EEG (2), särskilt artikel 9.1 i detta, och
med beaktande av följande: I artikel 7a i fördraget föreskrivs ett område utan inre gränser med fri rörlighet för varor, personer, tjänster och kapital.
I direktiv 76/116/EEG fastställs bestämmelser för saluföring av gödselmedel på den inre marknaden.
För att nya gödselmedel skall kunna dra fördel av den "EEG-märkning" som avses i bilaga II i direktiv 76/116/EEG måste de läggas till bilaga I till det direktivet.
I meddelande 94/C 138/04 (3) fastställs det förfarande som bör följas av dem (tillverkare eller dennes ombud) som vill att ett gödselmedel skall få betecknas som "EEG-gödselmedel" enligt bilaga II i direktiv 76/116/EEG, genom att lämna i sina tekniska uppgifter till medlemsstatens myndighet. Myndigheten fungerar som rapportör i Europeiska kommissionens arbetsgrupp för gödselmedel.
Åtgärderna i detta direktiv är förenliga med yttrandet från Kommittén för anpassning till teknisk utveckling av direktiven om avskaffandet av tekniska hinder för handel med gödselmedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till direktiv 76/116/EEG ändras på följande sätt:
1. Det gödselmedel som anges i bilaga I till detta direktiv skall läggas till del A punkt 1 "Kvävegödselmedel".
Följande produkt och tolerans läggs till under A.1 i bilaga III till direktiv 76/116/EEG:
>Plats för tabell>
Artikel 3
1. Medlemsstaterna skall anta de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 maj 1997. De skall genast underrätta kommissionen om detta.
2. Medlemsstaterna skall underrätta kommissionen om de nationella bestämmelser de antar inom det område som omfattas av detta direktiv.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV 96/42/EG av den 25 juni 1996 om ändring av direktiv 77/388/EEG om ett gemensamt system för mervärdeskatt
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
med beaktande av följande: I artikel 12.3 d i direktiv 77/388/EEG (3), anges att de regler som gäller beskattningen av andra jordbruksprodukter än dem som tillhör kategori 1 i bilaga H enhälligt skall antas av rådet på kommissionens förslag senast den 31 december 1994. Till och med denna dag tilläts de medlemsstater som redan tillämpade en reducerad skattesats behålla denna medan de som tillämpade normalskattesatsen inte fick använda en reducerad skattesats. Denna bestämmelse tillät en senareläggning av tillämpningen av normalskattesatsen med två år.
Erfarenheten visar att det har förekommit fall av bedräglig verksamhet på grund av den strukturella obalansen mellan de mervärdeskattesatser som medlemsstaterna tillämpar för jordbruksprodukter från blomster- och trädgårdsodling. Eftersom den strukturella obalansen direkt kan hänföras till tillämpningen av artikel 12.3 d bör detta ändras.
Den bästa lösningen består i att tillåta alla medlemsstater att provisoriskt tillämpa en reducerad skattesats för tillhandahållande av jordbruksprodukter från blomster- och trädgårdsodling samt av vedbränsle.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 77/388/EEG ändras på följande sätt:
1. I artikel 12.3 skall punkt d utgå.
2. Följande punkt skall införas i artikel 28.2:
"i) medlemsstaterna får tillämpa en reducerad skattesats för tillhandahållande av levande växter och andra produkter från blomsterodling (inklusive lökar, rötter och liknande produkter, snittblommor och prydnadsbladväxter) liksom för tillhandahållande av vedbränsle."
Artikel 2
Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 3
Detta direktiv gäller från och med den 1 januari 1995.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 96/57/EG av den 3 september 1996 om energieffektivitetskrav för elektriska kylskåp och frysar (även i kombination) för hushållsbruk
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
i enlighet med det i artikel 189b i fördraget angivna förfarandet (3), och
med beaktande av följande: 1. Det är viktig att främja åtgärder som syftar till att den inre marknaden fungerar väl.
2. I sin resolution av den 15 januari 1985 om förbättring av energibesparingsprogrammen i medlemsstaterna (4) uppmanade rådet medlemsstaterna att fortsätta och i förekommande fall öka sina ansträngningar att främja en mer rationell användning av energi genom att utveckla en samordnad politik i fråga om energibesparingsåtgärder.
3. Den elektricitet som förbrukas av kylskåp och frysar för hushållsbruk utgör en icke obetydlig del av hushållens elförbrukning och därigenom av gemenskapens totala elförbrukning. Elförbrukningen, dvs. energieffektiviteten, varierar kraftigt mellan de olika modeller av kylskåp och frysar med samma volym och egenskaper som erbjuds på gemenskapsmarknaden.
4. Några medlemsstater står i begrepp att anta bestämmelser om energieffektiviteten hos kylskåp och frysar för hushållsbruk, vilka bestämmelser är av sådant slag att de kan medföra handelshinder för dessa produkter inom gemenskapen.
5. Det är nödvändigt att utgå från en hög skyddsnivå när det gäller förslagen om tillnärmning av bestämmelser i medlemsstaternas lagar och andra författningar rörande hälsa, säkerhet, miljöskydd och konsumentskydd. Detta direktiv garanterar en hög skyddsnivå för miljön och konsumenterna samtidigt som det syftar till en betydande förbättring av kylskåps och frysars energieffektivitet.
6. Vidtagandet av sådana åtgärder omfattas av gemenskapens befogenheter. Kraven i detta direktiv går inte utöver vad som är nödvändigt för att uppnå direktivets mål och direktivet överensstämmer således med bestämmelserna i artikel 3b i fördraget.
7. I artikel 130r i fördraget föreskrivs dessutom att gemenskapens miljöpolitik skall bidra till bland annat målen att skydda och förbättra miljön samt att utnyttja naturresurserna varsamt och rationellt. Produktion och förbrukning av elektricitet bidrar till ungefär 30 % av koldioxidutsläpp (CO2) förorsakade av människor och motsvarar ungefär 35 % av gemenskapens bruttoenergiförbrukning och denna andel ökar.
8. Rådets beslut 89/364/EEG av den 5 juni 1989 om ett åtgärdsprogram för gemenskapen för förbättrad effektivitet i elutnyttjandet (5) har den dubbla målsättningen att uppmuntra konsumenterna att välja apparater och utrustning som är mest energieffektiva samt att förbättra apparaternas och utrustningens energieffektivitet.
9. I sina slutsatser av den 29 oktober 1990 fastställde rådet målet att till år 2000 stabilisera koldioxidutsläppen (CO2) i gemenskapen på 1990 års nivå. För att nå detta mål krävs kraftigare åtgärder för att stabilisera gemenskapens koldioxidutsläpp.
10. Genom rådets beslut 91/565/EEG (6) upprättades ett program för att främja effektiv energianvänding i gemenskapen (Save-programmet).
11. De åtgärder för en förbättrad energieffektivitet som genomförts på de senaste modellerna av kylskåp och frysar som finns på marknaden ökar inte påtagligt deras tillverkningskostnader och kan uppvägas inom några få år, eller till och med ännu snabbare, av de elektricitetsbesparingar de innebär. Denna beräkning tar inte hänsyn till den ytterligare fördel det innebär att externa kostnader i samband med elproduktionen försvinner, såsom exempelvis koldioxidutsläpp (CO2) och andra föroreningar.
12. Den energieffektivitetsvinst som automatiskt uppstår till följd av påtryckningar från marknaden och förbättringar av tillverkningsmetoderna och som uppskattas till ungefär 2 % per år, kommer att bidra till ansträngningarna att få till stånd strängare normer för energiförbrukning.
13. Direktiv 92/75/EEG (7) (ramdirektivet) och kommissionens direktiv 94/2/EG (8) (om genomförandet av direktiv 92/75/EEG) som föreskriver obligatorisk märkning av apparater och andra former av upplysningar om energiförbrukning kommer att öka konsumenternas medvetenhet om energieffektivitet hos kylskåp och frysar för hushållsbruk. Denna åtgärd kommer följaktligen även att leda till att de konkurrerande tillverkarna erbjuder apparater med högre energieffektivitet än vad som föreskrivs i direktivets normer. I konsumentupplysningarna bör normerna ändå anges för att de ska bli så effektiva som möjligt och leda till en verklig förbättring av de sålda apparaternas genomsnittliga samlade effektivitet.
14. Detta direktiv som syftar till att avlägsna tekniska hinder för en förbättrad energieffektivitet hos kylskåp och frysar för hushållsbruk skall följa den "nya metoden" som fastställs i rådets resolution av den 7 maj 1985 om en ny metod för teknisk harmonisering och standardisering (9) i vilken det uttryckligen bestäms att rättslig harmonisering begränsas till att genom direktiv anta de grundläggande krav vilka skall uppfyllas av varor som släpps ut på marknaden.
15. Det är viktigt att upprätta ett effektivt verktyg för att säkerställa ett felfritt genomförande av direktivet, rättvisa konkurrensvillkor för tillverkarna och skydd för konsumenternas rättigheter.
16. Hänsyn bör tas till beslut 93/465/EEG av den 22 juli 1993 om moduler för olika stadier i förfaranden vid bedömning av överensstämmelse samt regler inför anbringande och användning av CE-märkning om överensstämmelse, avsedda att användas i tekniska harmoniseringsdirektiv (10).
17. Med hänsyn till den internationella handeln bör internationell standard användas. Elförbrukningen för kylskåp och frysar definieras av Europeiska standardiseringsorganisationens standard EN 153 från juli 1995, på grundval av en internationell standard.
18. Kylskåp och frysar för hushållsbruk som överensstämmer med de energieffektivitetskrav som fastställs i detta direktiv skall förses med EG-märkning och tillhörande upplysningar för att möjliggöra deras fria rörlighet.
19. Detta direktiv omfattar inte kylskåp och frysar som tillverkats enligt särskilda specifikationer utan endast nätanslutna kylskåp och frysar för hushållsbruk, avsedda för livsmedel. Kyl- och frysanläggningar för kommersiellt bruk är avsevärt mer varierade och kan därför inte omfattas av detta direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Detta direktiv skall tillämpas på nya nätanslutna kylskåp, frysfack och frysar, även i kombination, för hushållsbruk, enligt bilaga I, nedan kallade "kyl- och frysapparater". Apparater som även kan utnyttja andra energikällor, t.ex. batterier, samt kyl- och frysapparater för hushållsbruk som bygger på absorptionsprincipen och apparater som tillverkats enligt särskilda specifikationer omfattas inte av direktivet.
Artikel 2
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att se till att de kyl- och frysapparater som omfattas av detta direktiv endast får släppas ut på marknaden i gemenskapen om deras elförbrukning är mindre än eller lika med den högsta tillåtna elförbrukningen för denna kategori apparater, vilken skall beräknas enligt de förfaranden som anges i bilaga I.
2. Tillverkaren av en kyl- och frysapparat som omfattas av detta direktiv, dennes i gemenskapen etablerade ombud eller den person som ansvarar för att apparaten släpps ut på marknaden inom gemenskapen åläggs att se till att varje apparat som släppts ut på marknaden uppfyller kravet som avses i punkt 1.
Artikel 3
1. Medlemsstaterna får inte inom sitt respektive territorium förbjuda, begränsa eller hindra att kyl- och frysapparater, försedda med den EG-märkning som intygar att de överensstämmer med samtliga bestämmelser i detta direktiv, släpps ut på marknaden.
2. Om det inte finns bevis om motsatsen skall medlemsstaterna utgå från att kyl- och frysapparater med EG-märkning enligt artikel 5 överensstämmer med samtliga bestämmelser i detta direktiv.
3. a) Om kyl- och frysapparater omfattas av andra direktiv i vilka andra frågor behandlas och i vilka EG-märkning också föreskrivs innebär denna märkning att sådana kyl- och frysapparater skall förutsättas överensstämma även med bestämmelserna i dessa direktiv om det inte finns bevis om motsatsen.
b) Om tillverkaren likväl under en övergångsperiod kan välja mellan att tillämpa olika bestämmelser i ett eller flera av dessa direktiv, anger EG-märkningen endast överensstämmelse med bestämmelserna i de direktiv som tillverkaren har tillämpat. I de handlingar, anvisningar och instruktioner som medföljer kyl- och frysapparaterna skall i så fall numren på dessa direktiv anges, enligt den text som offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 4
De förfaranden som skall tillämpas för bedömning av överensstämmelse och de skyldigheter som rör EG-märkning av kyl- och frysapparater anges i bilaga II.
Artikel 5
1. Apparaterna skall, då de släpps ut på marknaden, vara försedda med EG-märkning. Denna skall bestå av bokstäverna "CE". Den utformning som skall användas visas i bilaga III. EG-märkningen skall vara väl synlig, läsbar och outplånligt anbringad på kyl- och frysapparaterna samt vid behov på emballaget.
2. Det är förbjudet att på kyl- och frysapparaterna anbringa märkningar som skulle kunna vilseleda tredje man i fråga om EG-märkningens betydelse och grafiska utformning. Annan märkning får anbringas på apparaterna, emballaget, bruksanvisningen eller andra handlingar endast om EG-märkningen förblir synlig och läsbar.
Artikel 6
1. Om en medlemsstat konstaterar att EG-märkningen har använts på ett oriktigt sätt är tillverkaren eller dennes i gemenskapen etablerade ombud skyldig att anpassa produkten till bestämmelserna och upphöra med överträdelsen på de villkor som medlemsstaten föreskriver. Om varken tillverkaren eller dennes ombud är etablerade i gemenskapen åligger denna skyldighet den person som ansvarar för att kyl- och frysapparaten släpps ut på marknaden i gemenskapen.
2. Om överträdelsen fortgår skall medlemsstaten i enlighet med artikel 7 vidta alla nödvändiga åtgärder för att begränsa eller förbjuda att varan i fråga släpps ut på marknaden eller säkerställa att den tas ur försäljning.
Artikel 7
1. Alla beslut som fattas enligt detta direktiv och som innehåller inskränkningar av villkoren för att släppa ut kyl- och frysapparater på marknaden skall noga ange på vilka grunder beslutet är fattat. Den berörda parten skall omedelbart underrättas om beslutet och samtidigt få information om vilka möjligheter till överklagande som gäller i den berörda medlemsstaten och inom vilken tid detta skall äga rum.
2. Medlemsstaten skall utan dröjsmål underrätta kommissionen om och ange skälen för en sådan åtgärd. Kommissionen skall underrätta de övriga medlemsstaterna om detta.
Artikel 8
Senast fyra år efter det att detta direktiv har antagits skall kommissionen utvärdera de resultat som uppnåtts i förhållande till de förväntade resultaten. Med sikte på att gå vidare med nästa steg i förbättringen av energieffektiviteten skall kommissionen därefter i samråd med de berörda parterna undersöka om det finns behov av att upprätta ytterligare en rad lämpliga åtgärder för att på ett märkbart sätt förbättra energieffektiviteten för kyl- och frysapparater för hushållsbruk. Om så är fallet skall åtgärderna och tidpunkten för deras ikraftträdande grundas på energieffektivitetsnivåer som är ekonomiskt och tekniskt motiverade med hänsyn till de omständigheter som råder vid det tillfället. Andra åtgärder som har bedömts vara lämpliga för att förbättra effektiviteten för kyl- och frysapparater för hushållsbruk kommer också att beaktas.
Artikel 9
1. Medlemsstaterna skall anta och offentliggöra de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast inom ett år efter antagandet av detta direktiv. De skall omedelbart underrätta kommissionen om detta.
Medlemsstaterna skall tillämpa sådana bestämmelser tre år efter antagandet av detta direktiv.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser de antar inom det område som omfattas av detta direktiv.
3. Under en tid av tre år efter antagandet av detta direktiv skall medlemsstaterna tillåta att sådana kyl- och frysapparater släpps ut på marknaden som är godkända i respektive medlemsstat vid den tidpunkt detta direktiv antas.
Artikel 10
KOMMISSIONENS DIREKTIV 96/63/EG av den 30 september 1996 om ändring av rådets direktiv 76/432/EEG om bromsutrustning på jordbruks- eller skogsbrukstraktorer med hjul (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100 a i detta,
med beaktande av rådets direktiv 74/150/EEG av den 4 mars 1974 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av jordbruks- eller skogsbrukstraktorer med hjul (1), senast ändrat genom direktiv 88/297/EEG (2), särskilt artiklarna 12 och 13 i detta, och med beaktande av följande:
Bromsprovningstestet kan förbättras genom att medelretardationen ersätts med en formel som anger bromssträckan som en funktion av hastigheten. Denna ändring kommer att följas av ytterligare ändringar i syfte att öka säkerheten för traktorer och de element som berör deras användning.
Bestämmelserna i detta direktiv är förenliga med yttrandet från Kommittén för anpassning till tekniska framsteg, som upprättades i direktiv 74/150/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I och II som är bilagor till rådets direktiv 76/432/EEG (3) ändras i enlighet med bilagan till detta direktiv.
Artikel 2
1. Från och med den 1 oktober 1997 får medlemsstaterna inte
- vägra att bevilja EG-typgodkännande eller ett sådant dokument som avses i artikel 10.1 sista strecksatsen i direktiv 74/150/EEG eller nationellt typgodkännande för en traktortyp, eller
2. Från och med den 1 mars 1998 får medlemsstaterna
- inte längre bevilja EG-typgodkännande eller ett sådant dokument som avses i artikel 10.1 sista strecksatsen i direktiv 74/150/EEG, och
- får vägra att bevilja nationellt typgodkännande
för en traktortyp av skäl som hänför sig till bromsutrustningen, om kraven i direktiv 76/432/EEG, ändrat genom detta direktiv, inte är uppfyllda.
Artikel 3
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 1 oktober 1997. De skall genast underrätta kommissionen om detta.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
3. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 96/73/EG av den 16 december 1996 om vissa metoder för kvantitativ analys av binära textilfiberblandningar
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
i enlighet med det i artikel 189b i fördraget angivna fördraget (3), och
med beaktande av följande: Rådets direktiv 72/276/EEG av den 17 juli 1972 om tillnärmning av medlemsstaternas lagstiftning om vissa metoder för kvantitativ analys av binära textilfiberblandningar (4), har vid ett flertal tillfällen ändrats på väsentliga punkter. Av klarhets- och effektivitetsskäl bör direktivet kodifieras.
Europaparlamentets och rådets direktiv 96/74/EG av den 16 december 1996 om benämningar på textilier (5) föreskriver obligatorisk märkning för att ange vilka fibrer som ingår i textilvaror. Att märkningarna överensstämmer med innehållet i varorna kontrolleras genom analyser.
De metoder som används vid officiella provningar i medlemsstaterna för att bestämma fibersammansättningen för textilvaror bör vara enhetliga både vad beträffar förbehandlingen av provet och den kvantitativa analysen.
Direktivet 96/74/EG föreskriver att den provtagning och de analysmetoder som skall användas i medlemsstaterna för att bestämma fibersammansättningen i varor skall anges i särdirektiv. Följaktligen fastställs i bilaga II till detta direktiv femton enhetliga analysmetoder för de flesta på marknaden förekommande textilvaror som består av binära blandningar.
Den tekniska utvecklingen gör det nödvändigt att med täta mellanrum anpassa de tekniska specifikationer som definieras i särdirektiven om metoder för analys av textilier. För att underlätta genomförandet av de åtgärder som krävs för detta bör ett förfarande fastställas som upprättar ett nära samarbete mellan medlemsstaterna och kommissionen, i Kommittén för direktiv om benämningen och märkningen av textilier.
I fråga om binära blandningar för vilka det inte finns någon enhetlig analysmetod på gemenskapsnivå, får det laboratorium som ansvarar för provningen bestämma sammansättningen av sådana blandningar. De får därvid använda någon vedertagen metod och ange resultatet i analysrapporten samt hur tillförlitlig den använda metoden är, i den mån detta är känt.
Bestämmelserna i detta direktiv överensstämmer med det yttrande som avgivits av Kommittén för direktiv om benämningen och märkningen av textilier.
Detta direktiv skall inte påverka medlemsstaternas skyldigheter att överföra direktiven inom de tidsfrister som anges i bilaga III del B.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Detta direktiv gäller metoder för kvantitativ analys av vissa binära textilfiberblandningar, inklusive framtagning av analysprov och provexemplar.
Artikel 2
Analysprov avser ett med hänsyn till analysen lämpligt stort prov, som tas ut från laboratorieprovet, som i sin tur tagits ut från ett varuparti för analys.
Provexemplar avser den del av analysprovet som behövs för ett enskilt provningsresultat.
Artikel 3
Medlemsstaterna skall vidta alla nödvändiga åtgärder för att i enlighet med direktivet 96/74/EG säkerställa att bestämmelserna i bilaga I och II om metoder för den kvantitativa analysen av vissa binära blandningar, inklusive framtagningen av analysprov och provexemplar, tillämpas vid alla officiella provningar för att bestämma sammansättningen av de textilvaror som släpps ut på marknaden.
Artikel 4
Det laboratorium som ansvarar för provningen av binära blandningar för vilka det inte finns någon enhetlig analysmetod på gemenskapsnivå skall bestämma sammansättningen av sådana blandningar genom att använda en vedertagen metod och ange resultatet i analysrapporten och hur tillförlitlig den använda metoden är, i den mån detta är känt.
Artikel 5
1. Härmed inrättas en kommitté för direktiv om benämningen och märkningen av textilier (nedan kallad "kommittén"). Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
2. Kommittén skall själv fastställa sin arbetsordning.
3. Anpassning av metoderna för kvantitativ analys till den tekniska utvecklingen enligt bestämmelserna i bilaga II skall ske i enlighet med det förfarande som anges i artikel 6.
Artikel 6
1. När det förfarande skall tillämpas som anges i denna artikel skall ärendet hänskjutas till kommittén av ordföranden, antingen på hans eget initiativ eller på begäran av en företrädare för en medlemsstat.
2. Kommissionens företrädare skall till kommittén lämna ett förslag om åtgärder som skall beslutas. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande ärendet är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen, varvid medlemsstaternas röster skall vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
3. a) Kommissionen skall anta de föreslagna åtgärderna om det är förenligt med kommitténs yttrande.
b) Om förslaget inte är förenligt med kommitténs yttrande, eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas.
Rådet skall besluta med kvalificerad majoritet.
c) Om rådet inte har fattat något beslut inom tre månader från det att förslaget har mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 7
Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 8
Direktiven som nämns i bilaga III del A upphävs utan att detta påverkar medlemsstaternas skyldigheter vad gäller de tidsfrister för överförande som anges i bilaga III del B.
Hänvisningar till de upphävda direktiven skall uppfattas som hänvisningar till detta direktiv och läsas enligt jämförelsetabellen i bilaga IV.
Artikel 9
Detta direktiv riktar sig till medlemsstaterna.
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS DIREKTIV 96/75/EG av den 19 november 1996 om system för befraktning och prissättning inom området nationella och internationella transporter av varor på inre vattenvägar inom gemenskapen
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 75 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
i enlighet med det i artikel 189c i fördraget angivna röstningsförfarandet (3), och
med beaktande av följande: De tilltagande problem som rör överbelastning av vägtrafikleder och järnvägslinjer, transportsäkerheten, miljön, energisparande och medborgarnas livskvalitet kräver i allmänhetens intresse en längre driven utveckling och ett bättre utnyttjande av transportmöjligheterna på inre vattenvägar, genom bland annat förbättrad konkurrenskraft för dessa transporter.
Olikheterna i nationell lagstiftning i fråga om sätten att kommersiellt bedriva transport på inre vattenvägar gynnar inte den inre marknadens funktion inom denna sektor, och därför bör på gemenskapsnivå gemensamma bestämmelser införas för hela marknaden för transport på inre vattenvägar, i enlighet med rådets resolution av den 24 oktober 1994 om strukturella förbättringar av transport på inre vattenvägar (4).
För den inre marknadens funktion krävs det i fråga om varutransporter på inre vattenvägar att system med befraktning i turordning anpassas i riktning mot större kommersiell smidighet i syfte att skapa ett system med fri befraktning och fri prissättning för transporter.
För detta ändamål bör en övergångsperiod föreskrivas med en successiv begränsning av tillämpningsområdet för systemet med befraktning i turordning för att transportörerna skall kunna anpassa sig till den fria marknadens villkor och i förekommande fall genomföra former för kommersiella sammanslutningar som är bättre anpassade till avlastarnas logistiska behov.
Med hänsyn till subsidiaritetsprincipen är det både nödvändigt och tillräckligt att på gemenskapsnivå fastställa en enhetlig tidsplan för successiv liberalisering av marknaden, samtidigt som ansvaret för genomförandet av liberaliseringen överlåts på medlemsstaterna.
Det är viktigt att anta bestämmelser som gör det möjligt att ingripa på den aktuella transportmarknaden om en allvarlig störning skulle inträffa, och för detta ändamål bör kommissionen ges befogenhet att vidta lämpliga åtgärder i enlighet med förfarandet med rådgivande kommitté.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I detta direktiv avses med
a) system med befraktning i turordning: ett system som består i att transportförfrågningar från kundkretsen fördelas i en befraktningspool till fastställda priser och enligt offentliggjorda villkor, i den ordning som fartygen blir tillgängliga efter lossning. Transportörerna erbjuds, i den ordning de anmält sig till turordningen, att välja ut en transport bland dem som bjuds ut. De som inte väljer behåller likväl sin plats i turordningen,
b) transportör: den som äger eller bedriver transport med ett eller flera fartyg på inre vattenvägar,
c) behörig myndighet: myndighet som av medlemsstaten utsetts att förvalta och organisera systemet med befraktning i turordning,
d) allvarlig marknadsstörning: uppträdande på marknaden för varutransport på inre vattenvägar av specifika problem av ett slag som kan medföra ett allvarligt och eventuellt bestående överskott av utbud i förhållande till efterfrågan och som innebär ett allvarligt hot mot den ekonomiska stabiliteten och överlevnaden för ett betydande antal företag som transporterar varor på inre vattenvägar, under förutsättning att de kort- och medellångsiktiga prognoserna på den aktuella marknaden inte visar betydande och varaktiga förbättringar.
Artikel 2
Inom området nationella och internationella varutransporter på inre vattenvägar inom gemenskapen, skall avtal ingås fritt mellan berörda parter och priser förhandlas fritt.
Artikel 3
Med undantag från artikel 2 får medlemsstaterna under en övergångsperiod fram till den 1 januari 2000 upprätthålla ett system med obligatoriska minimitaxor och system med befraktning i turordning under förutsättning
- att de villkor som räknas upp i artikel 4, 5 och 6 efterlevs, och
- att systemen med befraktning i turordning och de fastställda priserna är fritt tillgängliga på samma villkor för alla transportörer i medlemsstaterna.
Artikel 4
Under den övergångsperiod som avses i artikel 3 skall följande undantas från tillämpningsområdet för befraktningssystem i turordning:
a) Transporter av olja och gas, flytande och torr last i bulk, specialtransporter av tungt och odelbart gods, containertransporter, transporter inom hamnområden, alla slags transporter för egen räkning samt alla slags transporter som redan utförs utanför systemet med befraktning i turordning.
b) Transporter som inte kan utföras effektivt av dessa system, bland annat
- transporter som kräver utrustning för godshantering,
- kombinerade transporter, det vill säga transporter med flera olika transportmedel där de huvudsakliga sträckorna utgörs av inre vattenvägar och där de inledande och/eller avslutande sträckorna, som skall vara så korta som möjligt, antingen utgör väg eller järnväg.
Artikel 5
Under den övergångsperiod som avses i artikel 3 skall medlemsstaterna vidta nödvändiga åtgärder för att så långt som möjligt göra systemen med befraktning i turordning mer flexibla, bland annat genom att
- föreskriva möjlighet för avlastarna att ingå avtal om flera transporter, det vill säga en serie på varandra följande transporter utförda av ett och samma fartyg,
- föreskriva att enstaka eller upprepade transporter, som erbjudits två gånger efter varandra inom systemet med befraktning i turordning utan att ha funnit någon användare, skall tas ur detta system och förhandlas fritt.
Artikel 6
Inom en frist på två år från och med ikraftträdandet av detta direktiv skall de medlemsstater som berörs av systemen med befraktning i turordning vidta nödvändiga åtgärder för att avlastarna fritt skall kunna välja mellan följande tre slag av avtal:
- Tidsavtal, inbegripet hyresavtal, enligt vilket transportören ställer ett eller flera fartyg med besättning till en kunds exklusiva förfogande för en fastställd tid för att transportera de varor den senare anförtror honom mot betalning av ett fastställt dagsbelopp. Avtalet skall ingås fritt mellan parterna.
- Tonnageavtal enligt vilket transportören förbinder sig att under en i avtalet fastlagd period transportera ett fastställt antal ton mot betalning av en fraktavgift per ton. Avtalet skall ingås fritt mellan parterna; det måste omfatta betydande godsmängder.
- Avtal om enstaka eller upprepade transporter.
Artikel 7
1. Vid allvarlig störning på marknaden får kommissionen, utan att det påverkar tillämpningen av rådets förordning (EEG) nr 1101/89 av den 27 april 1989 om strukturella förbättringar inom inlandssjöfarten (5), på en medlemsstats begäran vidta lämpliga åtgärder, bland annat åtgärder som syftar till att förhindra alla nya ökningar av den transportkapacitet som erbjuds på den ifrågavarande marknaden. Beslutet skall fattas i enlighet med förfarandet i artikel 8.2.
2. Om en medlemsstat begär lämpliga åtgärder, skall beslut fattas inom tre månader efter det att begäran har mottagits.
3. En medlemsstats begäran om att lämpliga åtgärder skall vidtas skall åtföljas av alla uppgifter som krävs för en bedömning av den ekonomiska situationen inom sektorn i fråga, bland annat
- uppgifter om genomsnittskostnader och priser för olika slags transporter,
- uppgift om i vilken grad lastutrymmet har utnyttjats,
- prognoser om utvecklingen av efterfrågan.
Upplysningarna får användas endast i statistiskt syfte. Det är förbjudet att använda dem för beskattningsändamål och att vidarebefordra dem till tredje man.
4. De beslut som fattas i enlighet med denna artikel, vilka inte får gälla längre än störningen på marknaden varar, skall medlemsstaterna utan dröjsmål underrättas om.
Artikel 8
1. Kommissionen skall biträdas av den kommitté som inrättats genom direktiv 91/672/EEG (6).
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är, i förekommande fall genom omröstning.
Yttrandet skall protokollföras, och dessutom har varje medlemsstat rätt att begära att få sin uppfattning tagen till protokollet.
Kommissionen skall ta största hänsyn till det yttrande som kommittén avgett. Den skall underrätta kommittén om det sätt på vilket dess yttrande har beaktats.
Artikel 9
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 1 januari 1997 och skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser, skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras, skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall genast till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 10
KOMMISSIONENS FÖRORDNING (EG) nr 242/96 av den 7 februari 1996 om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 3009/95 (2), särskilt artikel 9 i denna, och med beaktande av följande:
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
Det är lämpligt att bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning förfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen (3) ändrad genom Kommissionens förordning (EEG) nr 2454/93 (4), under en period av tre månader.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från sektionen för tulltaxe- och statistiknomenklatur inom tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan förfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapens officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 569/96 av den 29 mars 1996 om ändring av förordningarna (EEG) nr 1362/87 och (EEG) nr 1158/91 vad gäller interventionsuppköp och beviljande av stöd för privat lagring av skummjölkspulver och förordning (EEG) nr 1756/93 om avgörande faktorer för den jordbruksomräkningskurs som tillämpas för mjölk och mjölkprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter (1), senast ändrad genom kommissionens förordning (EG) nr 2931/95 (2), särskilt artiklarna 7.5 och 28 i denna,
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas inom den gemensamma jordbrukspolitiken (3), senast ändrad genom förordning (EG) nr 150/95 (4), särskilt artikel 6.2 i denna, och
med beaktande av följande: Rådets förordning (EEG) nr 1014/68 av den 20 juli 1968 om allmänna bestämmelser om offentlig lagring av skummjölkspulver (5), senast ändrad genom förordning (EEG) nr 3577/90 (6), upphörde att gälla från och med den 1 mars 1996 genom rådets förordning (EG) nr 1538/95 (7). Vissa bestämmelser i förordning (EEG) nr 1014/68 har införts i artikel 7 i förordning (EEG) nr 804/68 i dess ändrade lydelse genom förordning (EG) nr 1538/95. Kommissionens förordning (EEG) nr 625/78 av den 30 mars 1978 om tillämpningsföreskrifter för offentlig lagring av skummjölkspulver (8), senast ändrad genom förordning (EG) nr 1802/95 (9), omarbetades när den anpassades till följd av att förordning (EEG) nr 1014/68 upphävdes. Förordning (EEG) nr 625/78 har följaktligen likaså upphört att gälla från och med den 1 mars 1996 genom kommissionens förordning (EG) nr 322/96 av den 22 februari 1996 om tillämpningsföreskrifter för offentlig lagring av skummjölkspulver (10).
I kommissionens förordning (EEG) nr 1362/87 av den 18 maj 1987 om tillämpningsföreskrifter till rådets förordning (EEG) nr 777/87 med avseende på uppköp och beviljandet av stöd för privat lagring av skummjölkspulver (11), senast ändrad genom förordning (EG) nr 1137/94 (12), kommissionens förordning (EEG) nr 1158/91 av den 3 maj 1991 om interventionsorgans uppköp av skummjölkspulver genom anbud (13), senast ändrad genom förordning (EG) nr 1802/95, och kommissionens förordning (EEG) nr 1756/93 (14), senast ändrad genom förordning (EG) nr 315/96 (15), görs det hänvisningar till förordningarna (EEG) nr 1014/68 och (EEG) nr 625/78. I dessa förordningar bör det istället hänvisas till förordning (EG) nr 322/96. Dessutom bör förordning (EEG) nr 1158/91 ändras för att närmare fastställa sättet att beräkna uppköpspriset i förhållande till proteinhalten i skummjölkspulver.
Vad gäller stöd till privat lagring av skummjölkspulver föreskrivs det i artikel 5 i förordning (EEG) nr 1362/87 att kontraktsparten vid export av skummjölkspulver genom undantag från gällande bestämmelser kan sälja ut lager när en kontraktsperiod på 30 dagar har löpt ut. Denna undantagsbestämmelse används sällan och försvårar i onödan förvaltning av ordningen. Den bör därför upphävas.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 1362/87 ändras på följande sätt:
a) Punkt a skall ersättas med följande:
"a) har framställts av en produktionsenhet som förbundit sig att löpande föra de register som avses i artikel 2.1 b i förordning (EG) nr 322/96,".
b) Punkt e skall ersättas med följande:
3. Artikel 5 skall utgå.
Artikel 2
Förordning (EEG) nr 1158/91 ändras på följande sätt:
2. I artikel 3 skall punkt 1 ersättas med följande:
"1. Anbudsgivare får delta i anbudsförfaranden endast
- avseende skummjölkspulver som framställts under de 21 dagarna som omedelbart föregår den sista anbudsdagen; i det fall som avses i bilaga III e andra meningen i förordning (EG) nr 322/96 fastställs denna period till tre veckor,
- om de skriftligen åtar sig att följa artikel 4.6 i förordning (EG) nr 322/96."
3. I artikel 7.1 andra stycket skall punkt c ersättas med följande:
"c) Det lager dit det skall levereras. Artiklarna 5 och 6 i förordning (EG) nr 322/96 skall tillämpas."
4. Artikel 9 skall ersättas med följande:
"Artikel 9
Inom en period som börjar löpa den 120:e dagen efter övertagandet av skummjölkspulvret och som löper ut den 140:e dagen därefter, skall interventionsorganet betala anbudsgivare som tilldelats kontrakt det pris som anges i vederbörandes anbud. Betalning skall ske för varje övertagen kvantitet under förutsättning att kraven i artikel 1 andra stycket är uppfyllda.
Uppköpspriset skall beräknas på följande sätt:
- Om proteinhalten i den fettfria torrsubstansen är minst 35,6 % skall uppköpspriset vara det pris som anges i anbudet.
- Om proteinhalten i den fettfria torrsubstansen är lägre än 35,6 % men minst 31,4 % skall uppköpspriset vara det pris som anges i anbudet minskat med ett belopp "d" som räknas fram på följande sätt:
d = anbudspriset × [(0,356 - proteinhalten) × 1,75].
Proteinhalten fastställs enligt den metod som anges i bilaga I till förordning (EG) nr 322/96."
Bestämmelserna i artiklarna 2 och 3 i förordning (EG) nr 322/96 skall tillämpas."
Artikel 3
I bilagan till förordning (EEG) nr 1756/93 skall punkt 1 i avdelning C.I i del C och punkt 3 i del D ersättas med följande:
>Plats för tabell>
Artikel 4
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS FÖRORDNING (EG) nr 753/96 av den 22 april 1996 om ändring av förordning (EEG) nr 3906/89 i syfte att utvidga det ekonomiska stödet till att omfatta Bosnien-Hercegovina
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 235 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande (1), och
KOMMISSIONENS FÖRORDNING (EG) nr 779/96 av den 29 april 1996 om tillämpningsföreskrifter till rådets förordning (EEG) nr 1785/81 i fråga om informationslämnande inom sockersektorn
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1785/81 av den 30 juni 1981 om den gemensamma organisationen av marknaden för socker (1), senast ändrad genom förordning (EG) nr 1101/95 (2), särskilt artikel 39 i denna, och
med beaktande av följande: I artikel 39 i förordning (EEG) nr 1785/81 anges att medlemsstaterna och kommissionen skall lämna varandra de uppgifter som behövs för tillämpningen av förordningen. Således fastställdes tillämpningsbestämmelser i kommissionens förordning (EEG) nr 787/83 av den 29 mars 1983 om informationslämnande inom sockersektorn (3), senast ändrad genom förordning (EEG) nr 3819/85 (4). Med tanke på den utveckling som sedan skett av den gemensamma organisationen av marknaden för socker och särskilt gemenskapens åtaganden till följd av det jordbruksavtal som slöts efter Uruguayrundans multilaterala förhandlingar, finns det anledning att se över bestämmelserna i sin helhet och fastställa nya och att upphäva förordning (EEG) nr 787/83 inför regleringsåret 1996/97.
För att på ett korrekt sätt kunna bedöma situationen när det gäller socker som köpts eller sålts med stöd av de regler om interventionsåtgärder som fastställts i förordning (EEG) nr 1785/81 måste relevant information finnas, särskilt i fråga om de kvantiteter som hålls av interventionsorganen, samt om fördelningen av dessa kvantiteter på lager som godkänts i enlighet med artikel 1.2 i rådets förordning (EEG) nr 447/68 av den 9 april 1968 om allmänna bestämmelser för interventionsköp av socker (5), senast ändrad genom förordning (EEG) nr 1359/77 (6). För att kunna följa tillämpningen av interventionssystemet är det också viktigt att regelbundet få information om de kvantiteter socker som blivit otjänliga för konsumtion och de kvantiteter som har använts för att tillverka vissa kemiska produkter, varvid också måste anges de kvantiteter socker som antingen har denaturerats i enlighet med någon av de processer som beskrivs i bilagan till kommissionens förordning (EEG) nr 100/72 av den 14 januari 1972 om föreskrifter för denaturering av socker till foderändamål (7), senast ändrad genom förordning (EG) nr 260/96 (8), eller som använts vid tillverkning av de kemiska produkter som räknas upp i bilagan till rådets förordning (EEG) nr 1010/86 av den 25 mars 1986 om allmänna bestämmelser om produktionsbidrag för vissa sockerprodukter som används i den kemiska industrin (9), senast ändrad genom förordning (EG) nr 1101/95, samt de produkter som räknas upp i bilagan till kommissionens förordning (EEG) nr 1729/78 av den 24 juli 1978 om tillämpningsföreskrifter för produktionsbidrag för socker som används i den kemiska industrin (10), senast ändrad genom förordning (EG) nr 260/96.
För att noggrant kunna följa utvecklingen av handeln med tredje land behövs en nära och regelbunden övervakning med hänsyn till de intressekonflikter som kan uppkomma beroende på å ena sidan gemenskapens åtaganden inom ramen för ovan nämnda jordbruksavtal och åtgärder som kan behöva vidtas i samband med detta, särskilt i fråga om tillämpningen av artikel 23.4a i förordning (EEG) nr 1785/81, och å andra sidan gemenskapens åtaganden inom ramen för Internationella sockeravtalet. Det finns anledning för kommissionen att från början ha tillgång till relevant regelbunden information, inte bara vad gäller import och export av sådana produkter som omfattas av fastställda avgifter eller bidrag där licens utfärdas i enlighet med kommissionens förordning (EG) nr 1464/95 av den 27 juni 1995 om särskilda tillämpningsföreskrifter för systemet med import- och exportlicenser för socker (11), ändrad genom förordning (EG) nr 2136/95 (12), och när det gäller att iaktta de mera allmänna bestämmelserna i kommissionens förordning (EEG) nr 3719/88 (13), senast ändrad genom kommissionens förordningar (EG) nr 2137/95 (14) och (EEG) nr 3665/87 (15), senast ändrad genom förordning (EG) nr 1384/95 (16), utan även om import och export av sådana produkter som exporterats utan bidrag, med eller utan utfärdad licens, särskilt enligt bestämmelserna om aktiv förädling. Även importen av förmånssocker bör kunna följas för att ge möjlighet till effektiv tillämpning av bestämmelserna i kommissionens förordning (EEG) nr 2782/76 av den 17 november 1976 om fastställande av tillämpningsföreskrifter för import av förmånssocker (17), senast ändrad genom förordning (EEG) nr 1714/88 (18).
För att det kvoteringssystem som fastställts i avdelning III i förordning (EEG) nr 1785/81 skall fungera effektivt, är det nödvändigt att ha tillgång till all relevant information, särskilt med hänsyn till gemenskapens åtaganden inom ramen för nämnda jordbruksavtal. Detta berör tillämpningen av rådets förordning (EEG) nr 206/68 av den 20 februari 1968 om rambestämmelser för avtal och branschöverenskommelser rörande inköp av betor (19), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige, rådets förordning (EEG) nr 193/82 av den 26 januari 1982 om allmänna bestämmelser för överföring av kvoter inom sockersektorn (20), kommissionens förordning (EEG) nr 2670/81 av den 14 september 1981 om fastställande av tillämpningsföreskrifter för sockerproduktion utöver kvoten (21), senast ändrad genom förordning (EG) nr 158/96 (22), samt kommissionens förordning (EEG) nr 1443/82 av den 8 juni 1982 om tillämpningsföreskrifter för kvotsystemet på sockerområdet (23), senast ändrad genom förordning (EEG) nr 392/94 (24). Ovanstående gäller också för det system för kompensation för lagringskostnader som fastställts i artikel 8 i förordning (EEG) nr 1785/81. Därvid berörs tillämpningen av rådets förordning (EEG) nr 1358/77 av den 20 juni 1977 om allmänna bestämmelser för kompensation för lagringskostnader för socker, samt om upphävande av förordning (EEG) nr 750/68 (25), senast ändrad genom förordning (EEG) nr 3042/78 (26), liksom kommissionens förordning (EEG) nr 1998/78 av den 18 augusti 1978 om tillämpningsföreskrifter för kompensation för lagringskostnader för socker (27), senast ändrad genom förordning (EEG) nr 1758/93 (28).
De personer som berörs skall försäkras om att information som rör enskilda företag omfattas av tystnadsplikt.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för socker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Vad gäller interventionsåtgärder som vidtagits i enlighet med artiklarna 9.1 och 11.1 i förordning (EEG) nr 1785/81 skall varje medlemsstat varje vecka, med avseende på närmast föregående vecka, till kommissionen anmäla
a) de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som erbjudits men ännu inte tagits över av interventionsorganet,
b) de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som tagits över av interventionsorganet,
c) de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som sålts av interventionsorganet.
Artikel 2
På begäran av kommissionen skall varje medlemsstat överlämna en förteckning till kommissionen över de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som tagits över av interventionsorganet, samt över fördelningen av dessa kvantiteter på godkända lager.
Artikel 3
Vad gäller interventionsåtgärder som vidtagits i enlighet med artikel 9.2 i förordning (EEG) nr 1785/81 skall varje medlemsstat till kommissionen anmäla följande:
1. Varje vecka, med avseende på närmast föregående vecka, anmäla de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, för vilka en licens om denatureringsbidrag har utfärdats.
2. På begäran av kommissionen, med avseende på en bestämd period, anmäla de kvantiteter vitsocker och råsocker som har denaturerats och ange vilken av de metoder som anges i bilagan till förordning (EEG) nr 100/72, som har använts.
Artikel 4
Vad gäller interventionsåtgärder som vidtagits i enlighet med artikel 9.3 i förordning (EEG) nr 1785/81 skall varje medlemsstat till kommissionen anmäla följande:
1. Senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, anmäla de kvantiteter vitsocker, råsocker och sirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans för vilka:
a) en licens om produktionsbidrag har utfärdats,
b) ett produktionsbidrag har utbetalats.
2. Senast vid utgången av september månad varje år, med avseende på närmast föregående regleringsår, anmäla de kvantiteter vitsocker, råsocker och sirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans, fördelade på de produkter som räknas upp i bilagan till förordning (EEG) nr 1010/86, för vilka
a) en licens om produktionsbidrag har utfärdats,
b) ett produktionsbidrag har utbetalats.
3. Senast vid utgången av september månad varje år, med avseende på närmast föregående regleringsår, anmäla de kvantiteter basprodukter som avses i punkt 2 ovan vilka använts för framställning av sådana mellanprodukter som räknas upp i bilagan till förordning (EEG) nr 1729/78.
Artikel 5
Vad gäller export till tredje land skall varje medlemsstat till kommissionen anmäla följande:
1. Varje vecka, med avseende på närmast föregående vecka:
a) de kvantiteter för vilka licens har utfärdats med angivande av motsvarande exportbidrag fastställda i enlighet med artikel 17.5 andra stycket a i förordning (EEG) nr 1785/81, angivna var för sig enligt följande:
- vitsocker KN-nr 1701 91 00, 1701 99 10, 1701 99 90,
- råsocker angivet i icke omräknad vikt KN-nr 1701 11 90 och 1701 12 90,
- sackarossirap uttryckt som vitsocker KN-nr 1702 60 90, 1702 90 60, 1702 90 71, 1702 90 99 och 2106 90 59,
- isoglukos uttryckt som torrsubstans KN-nr 1702 40 10, 1702 60 10, 1702 90 30 och 2106 90 30,
- inulinsirap uttryckt som torrsubstans, socker/isoglukos ekvivalent, KN-nr ex 1702 60 90,
b) de kvantiteter vitsocker KN-nr 1701 99 10 för vilka licens har utfärdats med angivande av motsvarande exportbidrag fastställda i enlighet med artikel 17.5 andra stycket b i förordning (EEG) nr 1785/81,
c) de kvantiteter C-vitsocker, C-råsocker, C-isoglukos, C-inulinsirap, uttryckta som vitsocker, torrsubstans respektive som socker/isoglukos ekvivalent, för vilka exportlicens har utfärdats,
d) med angivande av exportbidrag fastställda i enlighet med artikel 17.5 andra stycket a i förordning (EEG) nr 1785/81 de kvantiteter vitsocker, råsocker och sackarossirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans, för vilka exportlicens har utfärdats för att exportera i form av produkter enligt artikel 1.1 b i rådets förordning (EEG) nr 426/86 (29).
2. Senast i slutet av varje kalendermånad, med avseende på närmast föregående kalendermånad, de kvantiteter vitsocker enligt punkt 1 b som exporterats i enlighet med artikel 8.4 och 8.5 i förordning (EEG) nr 3719/88.
3. För varje kalendermånad och senast vid utgången av den tredje månaden efter den kalendermånad som anmälan avser:
a) de kvantiteter - med angivande av exportbidrag för varje kvantitet - socker och sirap uttryckt som vitsocker, som avses i artikel 2 i förordning (EG) nr 1464/95, vilka exporterats i obearbetat skick utan exportlicens,
b) de kvantiteter socker ur kvoten som exporterats som vitsocker eller som bearbetad produkt uttryckt som vitsocker, för vilka exportlicens har utfärdats med anledning av livsmedelbistånd i gemenskapens eller nationell regi inom ramen för internationella överenskommelser eller andra kompletterande program eller till följd av andra åtgärder inom gemenskapen som avser kostnadsfri livsmedelstilldelning,
c) de kvantiteter socker och sackarossirap uttryckt som vitsocker, samt isoglukos uttryckt som torrsubstans, som exporterats obearbetat i enlighet med artikel 2a andra stycket i förordning (EEG) nr 3665/87 med angivande av motsvarande bidrag,
d) med angivande av exportbidrag fastställda i enlighet med artikel 17.5 andra stycket a i förordning (EEG) nr 1785/81 de kvantiteter vitsocker, råsocker och sackarossirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans, som exporterats i form av produkter enligt bilaga I i rådets förordning (EEG) nr 804/68 (30), samt produkter enligt bilagan till kommissionens förordning (EG) nr 1222/94 (31),
e) för export enligt 1 d och d i denna punkt de kvantiteter som exporterats utan bidrag.
De uppgifter som avses i d och e ovan skall lämnas var för sig till kommissionen i enlighet med de bestämmelser som gäller för respektive bearbetad produkt.
Artikel 6
Varje medlemsstat skall till kommissionen anmäla följande:
1. Varje vecka, med avseende på närmast föregående vecka, de kvantiteter vitsocker och råsocker angivna i icke omräknad vikt, förutom, förmånssocker, sirap, isoglukos och inulinsirap, för vilka importlicens har utfärdats.
2. För varje kvartal, senast vid utgången av den tredje kalendermånaden efter det kvartal anmälan avser, de kvantiteter socker, uttryckt som vitsocker, som
a) importerats från tredje land i form av bearbetade produkter enligt 5.1 d och 5.3 d,
b) importerats från eller exporterats till en annan medlemsstat i obearbetat skick eller i form av bearbetade produkter.
Artikel 7
Varje medlemsstat skall till kommissionen anmäla följande:
1. Varje vecka, med avseende på närmast föregående vecka, de kvantiteter vitsocker och råsocker angivna i icke omräknad vikt, för vilka import- eller exportlicens utfärdats i enlighet med artikel 10 i förordning (EG) nr 1464/95.
2. För varje kvartal, senast vid utgången av den andra kalendermånaden efter det kvartal anmälan avser, var för sig de kvantiteter socker som införts från tredje land och utförts i form av ersättningsprodukter inom ramen för förfarandet för aktiv förädling enligt definition i artikel 116 i förordning (EEG) nr 2913/92 (32).
Artikel 8
Vad gäller import av förmånssocker åligger följande varje medlemsstat:
1. Att senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, till kommissionen anmäla de kvantiteter socker, angivet i icke omräknad vikt, för vilka importlicenser har utfärdats i enlighet med förordning (EEG) nr 2782/76, med angivande av varje ursprungsland var för sig.
2. Att senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, till kommissionen vidarebefordra
a) kopior av relevanta varucertifikat EUR.1,
b) kopior av de dokument som avses i artikel 7.2 i förordning (EEG) nr 2782/76,
c) kopior, i förekommande fall, av den deklaration som avses i artikel 1.3 andra stycket i förordning (EEG) nr 2782/76.
De dokument som avses i a och b ovan skall förutom de uppgifter som anges i artiklarna 6 och 7 i förordning (EEG) nr 2782/76 innehålla uppgift, med en noggrannhet av sex decimaler, om graden av polarisering av varje importerad kvantitet.
3. Att senast vid utgången av oktober månad varje år till kommissionen överlämna en förteckning över intyg och attester som utfärdats i enlighet med artiklarna 6 och 7 i förordning (EEG) nr 2782/76 och ange
a) den totala kvantiteten vitsocker, angiven i ton,
b) den totala kvantiteten råsocker, angiven i ton i icke omräknad vikt,
c) den totala kvantiteten råsocker, angiven i ton i icke omräknad vikt, som är avsedd för direkt konsumtion,
som importerats i enlighet med förordning (EEG) nr 2782/76 till medlemsstaten under den leveransperiod som löper ut den 30 juni i frågavarande år.
Artikel 9
Varje medlemsstat skall till kommissionen anmäla följande:
1. Före den 1 mars varje år, med avseende på vart och ett av de sockerproducerande företagen och de företag som framställer inulinsirap, vilka är belägna på dess territorium, anmäla den beräknade socker- och inulinsirapproduktionen under det löpande regleringsåret fastställd i enlighet med artikel 3.1 i förordning (EEG) nr 1443/82. För de franska departementen Guadeloupe och Martinique samt för Spanien skall när det gäller rörsocker emellertid denna dag ersättas med den 1 juli.
2. Senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, anmäla produktionen av isoglukos, fastställd i enlighet med artikel 3.2 och punkt 2a i förordning (EEG) nr 1443/82, vid vart och ett av de isoglukosproducerande företagen på dess territorium. De kvantiteter isoglukos som varje månad producerats inom ramen för bestämmelserna om aktiv förädling skall redovisas separat.
3. Före den 15 september varje år för vart och ett av de sockerproducerande, isoglukosproducerande och inulinsirapproducerande företagen på dess territorium, anmäla den slutliga produktionen under det närmast föregående regleringsåret av socker, isoglukos och inulinsirap, fastställd i enlighet med artikel 3.3 i förordning (EEG) nr 1443/82.
Artikel 10
Varje medlemsstat skall varje kalendermånad, med avseende på den närmast föregående kalendermånaden, och allt efter vad som är lämpligt uttryckt som vitsocker, torrsubstans eller som socker/isoglukos ekvivalent, anmäla följande:
a) de kvantiteter socker, isoglukos och inulinsirap som avsatts på dess territorium för konsumtion,
b) de kvantiteter socker som har denaturerats,
Artikel 11
Utan att det påverkar tillämpningen av artikel 2.1 andra stycket i förordningen (EEG) nr 2670/81 skall varje medlemsstat före den 15 mars varje år, med avseende på närmast föregående regleringsår, till kommissionen anmäla de kvantiteter C-socker, C-isoglukos och C-inulinsirap som enligt artikel 1.1 i förordning (EEG) nr 2670/81 anses vara avsatt på gemenskapens inre marknad.
Artikel 12
Varje medlemsstat skall till kommissionen anmäla följande:
1. Före den femtonde dagen varje månad, med avseende på den närmast föregående kalendermånaden, anmäla de totala kvantiteter B-socker och C-socker som i förekommande fall har förts över enligt artikel 27 i förordning (EEG) nr 1785/81.
2. Före den 1 mars varje år, med avseende på det löpande regleringsåret och för vart och ett av de sockerproducerande företagen, anmäla de totala kvantiteter B-socker och C-socker som förts över till påföljande regleringsår.
Emellertid:
- vad gäller produktionen av betsocker i Spanien skall datumet den 1 mars ersättas med den 15 april,
Artikel 13
Varje medlemsstat skall till kommissionen anmäla följande:
1. De godkännanden som avses i artikel 2.1 c och d i förordning (EEG) nr 1358/77 samt i förekommande fall godkännanden som har dragits tillbaka med stöd av artikel 1 i förordning (EEG) nr 1998/78.
2. Före den femtonde dagen i varje månad, med avseende på den näst senaste kalendermånaden och på det sätt som framgår av exemplet i bilaga I anmäla
a) de kvantiteter som avses i artikel 4.2 i förordning (EEG) nr 1358/77,
b) de kvantiteter som har avsatts enligt artikel 12.1 i förordning (EEG) nr 1998/78.
Artikel 14
Varje medlemsstat skall till kommissionen anmäla följande:
1. Före den 1 september varje år, med avseende på närmast föregående regleringsår, och före den 1 januari varje år, med avseende på närmast föregående produktionsår, uppgifter rörande försörjningsbalanserna för socker, isoglukos och inulinsirap för ifrågavarande period enligt exemplet i bilaga II.
2. Före den 1 oktober efter varje regleringsår och med avseende på det regleringsåret uppgifter rörande försörjningsbalansen för melass enligt exemplet i bilaga III.
Artikel 15
Varje medlemsstat skall för varje kalendermånad och senast vid utgången av den tredje påföljande kalendermånaden till kommissionen lämna de statistiska uppgifter som rör gemenskapens åtaganden inom ramen för Internationella sockeravtalet i enlighet med exemplen i bilagorna IV och V.
Artikel 16
I denna förordning avses med
a) närmast föregående vecka: referensperioden från torsdag till onsdag,
b) närmast föregående kvartal: den tre månader långa referensperioden juli-september, oktober-december, januari-mars eller april-juni, allt efter vad som är aktuellt,
c) närmast föregående produktionsår: referensperioden från och med den 1 oktober ett kalenderår till och med den 30 september påföljande kalenderår.
Artikel 17
Kommissionen skall se till att den information som har överlämnats till den i enlighet med denna förordning blir tillgänglig för medlemsstaterna.
Om informationen innehåller upplysningar som rör ett enskilt företag, dess tekniska installationer eller arten och omfattningen av dess produktion, eller upplysningar som kunde göra det möjligt att rekonstruera sådana fakta, skall emellertid informationen endast lämnas till de personer som inom kommissionen är ansvariga för marknadsfrågor i sockersektorn. Sådan information får inte lämnas ut till tredje man.
Artikel 18
Artikel 19
Denna förordning träder i kraft den 1 juli 1996.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 2214/96 av den 20 november 1996 om harmoniserade konsumentprisindex: överföring och spridning av HIKP:s delindex (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2494/95 av den 23 oktober 1995 om harmoniserade konsumentprisindex (1), och
med beaktande av följande: Varje medlemsstat anmodas, enligt artikel 5,1 b i förordning (EG) nr 2494/95, att ta fram ett harmoniserat konsumentprisindex (HIKP) där ett första index skall gälla för januari 1997.
I artikel 9 i förordning (EG) nr 2494/95 krävs att medlemsstaterna behandlar insamlade data/uppgifter så att HIKP kan tas fram som omfattar kategorierna COICOP (Classification of individual consumption by purpose) och där dessa kategorier behöver anpassas.
I artikel 11 i förordning (EG) nr 2494/95 krävs att HIKP och motsvarande delindex skall publiceras av kommissionen (Eurostat). Dessa delindex behöver specifieras.
Det är nödvändigt att vidta åtgärder för att säkerställa att HIKP blir jämförbara enligt artikel 5.3 i förordning (EG) nr 2494/95.
De åtgärder som denna förordning föreskriver överensstämmer med yttrandet från Statistiska programkommittén (SPC), inrättad genom rådets beslut 89/382/EEG, Euratom (2).
Enligt artikel 5.3 i förordning (EG) nr 2494/95 har samråd skett med Europeiska monetära institutet som har avgett ett positivt yttrande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Mål
Målet för denna förordning är att fastställa delindexen till de harmoniserade konsumentprisindexen (HIKP) som varje månad skall beräknas och överlämnas till kommissionen (Eurostat) för vidare spridning.
Artikel 2
Definitioner
I denna förordning defineras ett "delindex till HIKP" som ett prisindex för en av de utgiftskategorier som anges i bilaga I och beskrivs i bilaga II till förordningen. De bygger på COICOP/HIKP-klassifikationen (Classification of individual consumption by purpose adopted to the needs of HICPs) (3). "Spridning" avser utlämnande av uppgifter i vilken form som helst.
Artikel 3
Framtagande och överföring av delindex
Medlemsstaterna skall varje månad beräkna och överlämna till kommissionen (Eurostat) alla delindex (bilaga I) som har en vikt som är större än en promille av de totala utgifterna som täcks av HIKP (4). Tillsammans med index för januari 1997 skall medlemsstaterna även till kommissionen (Eurostat) överföra motsvarande uppgifter om vikterna, och därefter vid varje tillfälle som vikterna ändras.
Artikel 4
Spridning av delindex
Kommissionen (Eurostat) skall låta sprida delindex av HIKP för de kategorier som anges i bilaga I till denna förordning där index för 1996=100.
Artikel 5
Kvalitetskontroll
Medlemsstaterna skall till kommissionen (Eurostat), på dess begäran, lämna information om fördelningen av varor och tjänster på de olika utgiftskategorierna i bilagorna I och II i tillräcklig omfattning för att kunna utvärdera att förordningen följs.
Artikel 6
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS BESLUT av den 28 januari 1997 om fastställandet av ett identifieringssystem för förpackningsmaterial i enlighet med Europaparlamentets och rådets direktiv 94/62/EG om förpackningar och förpackningsavfall (Text av betydelse för EES) (97/129/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets direktiv 94/62/EG av den 20 december 1994 om förpackningar och förpackningsavfall (1), särskilt artikel 8.2 i detta, och
med beaktande av följande: Identifieringssystemet skall vara frivilligt, åtminstone i ett inledande skede, men det skall genomgå en översyn för att fastställa om det skall införas på obligatorisk grund i ett senare skede.
Identifieringssystemet kommer regelbundet att ses över och kommer, vid behov, att ändras genom det förfarande som fastställts i artikel 21 i direktiv 94/62/EG.
De åtgärder som avses i detta beslut är förenliga med yttrandet från den kommitté som inrättas genom artikel 21 i direktiv 94/62/EG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Målet med detta beslut, vilket omfattar alla förpackningar enligt direktiv 94/62/EG, är att fastställa den numrering och de förkortningar som identifieringssystemet bygger på och ange vilket/vilka förpackningsmaterial som använts, samt specificera vilka material som bör omfattas av identifieringssystemet.
Artikel 2
I detta beslut skall följande gälla:
- De definitioner som anges i artikel 3 i direktiv 94/62/EG skall gälla om tillämpligt.
- Kompositmaterial betecknar förpackningar gjorda av olika material som inte kan separeras för hand och som inte i något fall överstiger en viss viktprocent som skall fastställas enligt det förfarande som anges i artikel 21 i direktiv 94/62/EG. Eventuella undantag för vissa material får fastställas genom samma förfarande.
Artikel 3
Numreringen och förkortningarna i identifieringssystemet skall vara de som anges i bilagorna.
Användningen av dessa skall vara frivillig när det gäller de plastmaterial som anges i bilaga I, papper och papp som anges i bilaga II, de metaller som anges i bilaga III, de trämaterial som anges i bilaga IV, de textilmaterial som anges i bilaga V, de glasmaterial som anges i bilaga VI och de kompositmaterial som anges i bilaga VII.
Beslut om att införa ett obligatoriskt identifieringssystem för något av materialen får antas enligt det förfarande som anges i artikel 21 i direktiv 94/62/EG.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 12 februari 1997 om precisering av principer för inkomst från institut för kollektiv investering, för tillämpning av rådets direktiv 89/130/EEG, Euratom om harmonisering av beräkningen av bruttonationalinkomst till marknadspris (Text av betydelse för EES) (97/157/EG, Euratom)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Fördraget om upprättandet av Europeiska atomenergigemenskapen,
med beaktande av rådets direktiv 89/130/EEG, Euratom av den 13 februari 1989 om harmonisering av beräkningen av bruttonationalinkomst till marknadspris (1), och
med beaktande av följande: För att kunna fastställa bruttonationalinkomsten till marknadspris (BNImp) i enlighet med artikel 1 i direktiv 89/130/EEG, Euratom, som enligt artikel 8.1 i rådets förordning (EG) nr 2223/96 av den 25 juni 1996 om det europeiska national- och regionalräkenskapssystemet i gemenskapen (2) skall fortsätta att tillämpas så länge som beslut 94/728/EG, Euratom (3) gäller, är det nödvändigt att klargöra principerna för inkomst från institut för kollektiv investering i enlighet med gällande upplaga av Europasystemet för integrerad ekonomisk redovisning (ENS).
I nuvarande upplaga av ENS beskrivs inte närmare hur inkomst från institut för kollektiv investering skall bokföras, och detta gäller i synnerhet för ej utdelad inkomst.
Det är därför nödvändigt att uttolka reglerna för nuvarande upplaga av ENS i enlighet med dessa grundprinciper, så att det kan fastställas hur denna inkomst skall bokföras.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som inrättas genom artikel 6 i direktiv 89/130/EEG, Euratom,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
För tillämpning av direktiv 89/130/EEG, Euratom skall inkomst från institut för kollektiv investering definieras dels som erhållen ränta från inlåning och värdepapper, dels som utdelning på aktier vilka innehas av instituten för kollektiv investering. Denna inkomst kan delas ut till aktieägare eller läggas till kapitalet.
Om utdelning sker, skall denna inkomst föras till aktieägarnas inkomstfördelningskonto som kapital- och företagarinkomster (post R40 i gällande ENS).
Om det inte sker någon utdelning av inkomsten, skall denna behandlas som en inkomst utbetald av institutet för kollektiv investering till dess aktieägare, som dessa omedelbart återinvesterar i institutet för kollektiv investering. Detta innebär att inkomsten måste bokföras som kapital- och företagarinkomster på samma sätt som när det gäller utdelning av inkomst. Motsvarande summa kommer att bokföras på aktieägarnas finanskonto under posten aktier.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 17 februari 1997 om förfarandet för bestyrkande av överensstämmelse av byggprodukter enligt artikel 20.2 i rådets direktiv 89/106/EEG beträffande konstruktionsvirke o.d. med tillbehör (Text av betydelse för EES) (97/176/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 89/106/EEG av den 21 december 1988 om tillnärmning av medlemsstaternas lagar och andra författningar om byggprodukter (1), ändrat genom direktiv 93/68/EEG (2), särskilt artikel 13.4 i detta, och med beaktande av följande:
Kommissionen skall välja det av de två förfaranden enligt artikel 13.3 i direktiv 89/106/EEG för bestyrkande av överensstämmelse av en produkt, som är "minst betungande och samtidigt förenligt med kraven på säkerhet". Detta innebär att det är nödvändigt att besluta huruvida en tillverkningskontroll i fabriken under tillverkarens ansvar är erforderlig och tillräcklig för bestyrkande av överensstämmelse för en bestämd produkt eller produktgrupp, eller om det av orsaker som rör uppfyllandet av de kriterier som avses i artikel 13.4 krävs att ett godkänt certifieringsorgan deltar.
Enligt artikel 13.4 i direktiv 89/106/EEG krävs att det förfarande som sålunda bestämts anges i uppdragen och i de tekniska specifikationerna. Det är därför önskvärt att definiera de produkter eller produktgrupper som används i uppdragen och i de tekniska specifikationerna.
De två förfarandena i artikel 13.3 beskrivs i detalj i bilaga III till direktiv 89/106/EEG. Det är därför nödvändigt att, i enlighet med bilaga III, klart specificera de metoder med vilka de två förfarandena skall genomföras för varje produkt eller produktgrupp, eftersom bilaga III anger att vissa system i första hand skall användas.
Det förfarande som avses i artikel 13.3 a motsvarar de system som anges i det första alternativet utan fortlöpande övervakning, samt i det andra och det tredje alternativet i punkt 2 ii i bilaga III och det förfarande som avses i artikel 13.3 b motsvarar de system som anges i punkt 2 i i bilaga III samt i det första alternativet med fortlöpande övervakning i punkt 2 ii i bilaga III.
Det åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga byggkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
För de produkter och produktgrupper som anges i bilaga I skall överensstämmelsen bestyrkas genom ett förfarande där tillverkaren ensam ansvarar för ett tillverkningskontrollsystem i fabriken som säkerställer att produkten överensstämmer med de relevanta tekniska specifikationerna.
Artikel 2
För de produkter som anges i bilaga II skall överensstämmelsen bestyrkas genom ett förfarande där, förutom ett tillverkningskontrollsystem i fabriken som genomförs av tillverkaren, även ett godkänt certifieringsorgan deltar vid bedömningen och övervakningen av tillverkningskontrollen eller av själva produkten.
Artikel 3
Förfarandet för bestyrkande av överensstämmelse enligt bilaga III skall anges i uppdragen för harmoniserade standarder.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 2 oktober 1997 om ändring av beslut 93/53/EEG om inrättande av en vetenskaplig kommitté för ursprungsbeteckningar, geografiska beteckningar och särartsskydd (Text av betydelse för EES) (97/656/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, och
med beaktande av följande: Det är lämpligt att närmare fastställa de villkor som skall gälla för medlemmarna i kommittén i deras tjänsteutövande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Enda artikel
Beslut 95/53/EEG ändras på följande sätt:
1. Den första meningen i artikel 6.1 skall ersättas med följande:
"Medlemmarna skall utses för en period på tre år."
2. Artikel 6.2 skall ersättas med följande:
"Efter utgången av treårs- eller tvåårsperioden skall medlemmarna, ordföranden och vice ordföranden sitta kvar tills de ersätts eller deras mandat förnyas."
3. Artikel 9 skall ersättas med följande:
2. De får inte för yrkesmässiga syften använda de uppgifter som kommit till deras kännedom under och efter deras mandat som medlemmar i kommittén."
Medlemmarna skall åta sig att undvika alla intressekonflikter under det att de utövar sina uppdrag."
KOMMISSIONENS BESLUT av den 11 december 1997 om upphävande av kommissionens beslut 97/613/EG och om införande av särskilda villkor för import av pistaschmandlar och vissa produkter som är framställda av dessa, som har sitt ursprung i eller försänds från Iran (Text av betydelse för EES) (97/830/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 93/43/EEG (1) av den 14 juni 1993 om livsmedelshygien, särskilt artikel 10.1 i detta, och med beaktande av följande:
Kommissionens beslut 97/613/EG (2) av den 8 september 1997 om ett tillfälligt förbud mot import av pistaschmandlar och vissa produkter som är framställda från dessa, som har sitt ursprung i eller försänds från Iran gäller fram till den 15 december 1997 och bör upphävas.
Pistaschmandlar som har sitt ursprung i Iran eller som försänds från Iran har i många fall visat sig innehålla alltför höga halter av aflatoxin B1.
Vetenskapliga livsmedelskommittén har konstaterat att aflatoxin B1, även i mycket små mängder, orsakar levercancer och att ämnet dessutom är genotoxiskt.
Detta utgör en allvarlig fara för folkhälsan i gemenskapen och det är absolut nödvändigt att vidta skyddsåtgärder på gemenskapsnivå.
De undersökningar som genomförts av de hygieniska förhållandena i Iran har visat att det krävs förbättrad hygienpraxis, och att pistaschmandlarna måste kunna spåras. Undersökningsgruppen lyckades inte kontrollera alla steg i hanteringen av pistaschmandlarna för export. De iranska myndigheterna har dock gjort åtaganden, i synnerhet beträffande förbättringar i fråga om produktion, hantering, sortering, bearbetning, förpackning och transport. Därför är det lämpligt att pistaschmandlar och produkter som är framställda av dessa, som har sitt ursprung i eller försänds från Iran, underkastas vissa särskilda villkor i syfte att säkerställa en hög skyddsnivå för folkhälsan.
Pistaschmandlar och produkter som är framställda av dessa, som har sitt ursprung i eller försänds från Iran får importeras under förutsättning att dessa särskilda villkor uppfylls.
Pistaschmandlar och vissa produkter som är framställda av dessa skall ha producerats, sorterats, hanterats, bearbetats, förpackats och transporterats i överensstämmelse med god hygienisk sed. Det är nödvändigt att fastställa halten av aflatoxin B1 och den totala aflatoxinhalten i prover tagna från sändningen omedelbart innan den lämnar Iran.
De iranska myndigheterna måste tillhandahålla dokumenterade bevis rörande villkoren för produktion, sortering, hantering, bearbetning, förpackning och transport samt resultaten av laboratorieundersökningar av sändningen beträffande halten av aflatoxin B1 och den totala aflatoxinhalten; denna dokumentation måste åtfölja varje sändning av pistaschmandlar som har sitt ursprung i Iran eller som försänds från Iran.
Partier med pistaschmandlar som har sitt ursprung i eller försänds från andra länder utanför EU bör underkastas analyser för att fastställa pistaschmandlarnas halter av aflatoxin B1 och den totala aflatoxinhalten, oberoende av varifrån pistaschmandlarna kommer. De samordnade programmen för officiell kontroll av livsmedel bör därför kompletteras.
Samråd har ägt rum med medlemsstaterna den 29 oktober 1997 och den 10 november 1997.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Detta beslut upphäver beslut 97/613/EG av den 8 september 1997 om ett tillfälligt förbud mot import av pistaschmandlar och vissa produkter som är framställda från dessa, som har sitt ursprung i eller försänds från Iran.
Artikel 2
1. Medlemsstaterna får importera
- pistaschmandlar som omfattas av KN-nummer 0802 50 00,
- rostade pistaschmandlar som omfattas av KN-numren 2008 19 13 och 2008 19 93,
som har sitt ursprung i eller som försänds från Iran, under förutsättning att sändningen åtföljs av officiella provtagnings- och analysresultat samt av ett hälsointyg enligt bilaga I, ifyllt, undertecknat och kontrollerat av en företrädare för det iranska hälsoministeriet.
2. Pistaschmandlar och produkter som är framställda från dessa, och som har sitt ursprung i, eller sänds från Iran, skall endast införas i gemenskapen via en av de införselorter som anges i bilaga II.
3. Varje sändning skall identifieras med en kod som motsvarar koden på provtagnings- och analysresultaten från den officiella provtagningen och analysen, och på det hälsointyg som avses i punkt 1.
4. De behöriga myndigheter i varje medlemsstat skall säkerställa att importerade pistaschmandlar som har sitt ursprung i, eller sänds från Iran, underkastas dokumentkontroller i syfte att säkerställa att sändningarna överensstämmer med de krav för hälsointyg och provtagningsresultat som avses i punkt 1.
5. De behöriga myndigheterna skall säkerställa att prover tas från varje sändning och att dessa analyseras för att fastställa halten av aflatoxin B1 och den totala aflatoxinhalten, och skall informera kommissionen om resultaten av dessa analyser.
Artikel 3
Detta beslut skall tas upp till förnyad behandling senast den 31 oktober 1998, för att bedöma huruvida de särskilda villkor som avses i artikel 2 ger ett tillräckligt skydd av folkhälsan i gemenskapen. Vid översynen skall också fastställas om det finns fortsatt behov av de särskilda villkoren.
Artikel 4
Medlemsstaterna skall vidta de åtgärder som krävs för att följa detta beslut. De skall underrätta kommissionen om detta.
Artikel 5
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS DIREKTIV 97/37/EG av den 19 juni 1997 om anpassning av bilaga I och II till Europaparlamentets och rådets direktiv 96/74/EG om benämningar på textilier till den tekniska utvecklingen (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets direktiv 96/74/EG av den 16 december 1996 om benämningar på textilier (1), särskilt artikel 16.1 i detta, och
med beaktande av följande: Textilprodukter får endast införas på gemenskapsmarknaden om de uppfyller direktivets bestämmelser.
Detta direktiv om benämningar på textilier föreskriver etiketter eller märkning eller angivelse av benämningarna på produktens textilfibrer för att säkerställa att konsumenternas intressen säkras genom rätt information.
Endast textilfibrerna i förteckningen i bilaga I till nämnda direktiv får användas vid sammansättning av textilprodukter som är avsedda för gemenskapens inre marknad. Det är nödvändigt att anpassa bilagornas förteckningar över fibrer till den tekniska utvecklingen genom att tillföra nya fibrer som har införts på marknaden efter den senaste ändringen av direktivet.
Detta direktivs bestämmelser är i enlighet med det yttrande som Kommittén för direktiv om benämningen och märkningen av textilier har avgett.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till direktiv 96/74/EG ändras på följande sätt:
1) Nummer 2 ändras på följande sätt:
- I kolumnen "beteckning" förs "kashgora" in efter "guanaco".
- I kolumnen "beskrivning" läggs "kashgoraget" (en korsning mellan kashmirget och angoraget) till efter "guanaco".
2) Nummer 30 ändras på följande sätt:
- Texten i kolumnen "beteckning" skall vara "polyamid eller nylon".
3) Numren 31-41 ersätts med 34-44.
4) Ett nytt nr 31 införs enligt följande:
"fiber bildad av syntetiska linjära makromolekyler bestående av aromatiska grupper som binds samman med amid- eller imidbindningar, av vilka minst 85 % binds direkt till två aromatiska ringar och där imidbindningarna, om sådana finns, till antalet inte får överskrida antalet amidbindningar."
5) Ett nytt nr 32 införs enligt följande:
- Texten i kolumnen "beteckning" skall vara "polyimid".
6) Ett nytt nr 33 införs enligt följande:
"fiber av regenererad cellulosa som fås genom upplösning och en spinnprocess i organiskt lösningsmedel utan att derivats bildas".
- En hänvisning till fotnoten har bifogats efter texten i kolumnen "beteckning". Fotnotens text skall vara följande:
"Med `organiskt lösningsmedel` avses en blandning av organiska ämnen och vatten."
"fiber av regenererad cellulosa som erhålls genom en ändrad viskosprocess och som har en hög hållfasthet och en hög våtmodul. Hållfastheten (BC) i konditionerat provningstillstånd och den dragkraft (BM) som krävs för att åstadkomma en förlängning om 5 % i vått tillstånd är följande:
Artikel 2
Bilaga II till direktiv 96/74/EEG ändras på följande sätt:
1) Numren 31-41 ersätts med 34-44.
2) Ett nytt nr 31 införs enligt följande:
Texten i kolumnerna "benämning" och "procentsatser" skall vara följande:
>Plats för tabell>
3) Ett nytt nr 32 införs enligt följande:
Texten i kolumnerna "benämning" och "procentsatser" skall vara följande:
>Plats för tabell>
4) Ett nytt nr 33 införs enligt följande:
Texten i kolumnerna "benämning" och "procentsatser" skall vara följande:
>Plats för tabell>
Artikel 3
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa direktiv 96/74/EG senast den 1 juni 1998.
De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 97/52/EG av den 13 oktober 1997 om ändring av direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG om samordning av förfarandena vid tilldelning av kontrakt vid offentlig upphandling av tjänster, varor samt bygg- och anläggningsarbeten
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 57.2, 66 och 100a i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
i enlighet med det i artikel 189b i fördraget angivna förfarandet (3), och
med beaktande av följande: 1. Genom sitt beslut 94/800/EG av den 22 december 1994 om ingående, på Europeiska gemenskapens vägnar - såvitt avser frågor som omfattas av dess behörighet - av de överenskommelser som är resultatet av de multilaterala förhandlingarna inom Uruguayrundan (1986 1994) (4) godkände rådet på Europeiska gemenskapens vägnar bland annat avtalet om offentlig upphandling, nedan kallat "avtalet", vars syfte är att införa ett multilateralt system av väl avvägda rättigheter och skyldigheter när det gäller offentlig upphandling för att liberalisera och utvidga världshandeln. Detta avtal har inte direkt effekt.
2. Genom direktiven 92/50/EEG (5), 93/36/EEG (6) och 93/37/EEG (7) samordnades de nationella förfarandena vid tilldelning av offentliga tjänstekontrakt, varukontrakt respektive bygg- och anläggningskontrakt för att införa rättvisa konkurrensvillkor för sådana kontrakt i alla medlemsstater.
3. De upphandlande myndigheter som omfattas av avtalet rättar sig efter direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG, i dessas lydelse enligt det här direktivet, och tillämpar samma bestämmelser som gäller för tjänsteleverantörer, leverantörer och entreprenörer i tredje land som undertecknat avtalet, handlar i enlighet med avtalet.
4. Med tanke på de internationella rättigheter och åtaganden som ett godtagande av avtalet medför för Europeiska gemenskapen, bör det system som tillämpas på anbudsgivare och varor från tredje land som undertecknat avtalet vara det som anges i avtalet, vars räckvidd när det gäller direktiv 92/50/EEG inte omfattar tjänstekontrakt enligt bilaga I B, kontrakt om forsknings- och utvecklingstjänster enligt kategori 8 i bilaga I A därtill, kontrakt om telekommunikationstjänster enligt kategori 5 i bilaga I A därtill med referensnummer enligt den allmänna klassificeringen av produkter (CPC) 7524, 7525 och 7526 eller kontrakt om finansiella tjänster enligt kategori 6 i bilaga I A därtill i samband med utfärdande, försäljning, förvärv eller överförande av värdepapper eller andra finansiella instrument samt i samband med tjänster som utförs av centralbanker.
5. Vissa av avtalets bestämmelser medför fördelaktigare villkor för anbudsgivande företag än de som framgår av direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG.
6. När upphandlande myndigheter tilldelar ett kontrakt på sätt som avses med avtalet, måste möjligheterna att få tillgång till offentliga tjänste-, varu- samt bygg- och anläggningskontrakt som i enlighet med fördraget är tillgängliga för företag och produkter från medlemsstater, vara minst lika förmånliga som villkoren för tillgång till sådana offentliga upphandlingskontrakt inom Europeiska unionen som enligt bestämmelserna i avtalet tillämpas för företag och produkter med ursprung i tredje land som undertecknat avtalet.
7. Det är därför nödvändigt att anpassa och komplettera bestämmelserna i direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG.
8. Tillämpningen av dessa direktiv måste förenklas samtidigt som jämvikten i gemenskapens gällande lagstiftning om offentlig upphandling måste bibehållas så långt det är möjligt.
9. Därför bör tillämpligheten av vissa av anpassningarna i direktiv 92/50/EEG utökas till att gälla alla tjänster som omfattas av detta direktiv.
10. Upphandlande myndigheter får begära eller ta emot råd som kan användas för att upprätta specifikationer för ett bestämt upphandlingsförfarande under förutsättning att dessa råd inte hindrar konkurrensen.
11. Kommissionen bör tillhandahålla små och medelstora företag utbildnings- och informationsunderlag för att göra det möjligt för dem att fullt ut delta i det ändrade upphandlingsförfarandet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
A) ersätts punkterna 1 och 2 med följande text:
"1. a) Det här direktivet gäller för
- de offentliga kontrakt avseende tjänster som avses i artikel 3.3, de offentliga kontrakt avseende sådana tjänster som avses i bilaga I B, tjänster i kategori 8 i bilaga I A och telekommunikationstjänster i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, förutsatt att det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 200 000 ecu,
- de offentliga kontrakt avseende sådana tjänster som avses i bilaga I A, med undantag för tjänster i kategori 8 och telekommunikationstjänster i kategori 5, med CPD-referensnumren 7524, 7525 och 7526,
i) som tilldelas av de upphandlande myndigheter som anges i bilaga I till direktiv 93/36/EEG, förutsatt att det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 130 000 särskilda dragningsrätter (SDR) i ecu,
ii) som tilldelas av de upphandlande myndigheter som anges i artikel 1 b utom dem som nämns i bilaga I till direktiv 93/36/EEG och vilkas uppskattade värde, exklusive mervärdesskatt, uppgår till minst 200 000 SDR i ecu.
b) Motvärdena i ecu och nationella valutor för de tröskelvärden som fastställs i a skall i princip revideras vartannat år med verkan från den 1 januari 1996. Beräkningen av detta motvärde skall grundas på den genomsnittliga dagskursen för dessa valutor uttryck i ecu och för ecun uttryckt i SDR under de sista 24 månaderna fram till den sista augusti som föregår revisionen per den 1 januari.
Den beräkningsmetod som avses i den här punkten skall på förslag av kommissionen ses över av Rådgivande kommittén för offentlig upphandling, i princip två år efter det att den tillämpats för första gången.
c) De tröskelvärden som framgår av a och deras motvärden uttryckta i ecu och i nationella valutor skall offentliggöras i Europeiska gemenskapernas officiella tidning i början av november månad efter den revision som anges i b i det här stycket.
2. Vid beräkning av det uppskattade värdet av ett kontrakt skall den upphandlande myndigheten inkludera den uppskattade, sammanlagda ersättningen till tjänsteleverantören med beaktande av bestämmelserna i punkterna 3 7."
B) Punkt 8 utgår.
2. Artikel 12.1 och 12.2 ersätts med följande text:
"1. Den upphandlande myndigheten skall inom 15 dagar efter att ha mottagit en skriftlig begäran underrätta varje anbudssökande eller anbudsgivare vars ansökan eller anbud har förkastats om orsakerna till att hans ansökan eller anbud förkastats samt underrätta varje anbudsgivare som lämnat ett godtagbart anbud om utformningen av och de relativa fördelarna med det antagna anbudet samt namnet på den anbudsgivare som tilldelats kontraktet.
De upphandlande myndigheterna får emellertid besluta att viss information som rör tilldelningen av kontrakt och som nämns i första stycket inte skall lämnas ut om det bedöms att detta skulle hindra lagarnas tillämpning eller strida mot allmänintresset eller vara till skada för offentliga eller privata företags legitima kommersiella intressen eller för lojal konkurrens mellan tjänsteleverantörer.
2. De upphandlande myndigheterna skall så snart som möjligt underrätta de anbudssökande och anbudsgivarna om de beslut som fattas rörande tilldelningen av kontrakt, inklusive skälen till att de har beslutat att avstå från en upphandling för vilken anbud begärts eller att upprepa förfarandet; dessa upplysningar skall på begäran lämnas skriftligen. Myndigheterna skall även underrätta Byrån för Europeiska gemenskapernas officiella publikationer om dessa beslut."
3. Artikel 13.1 och 13.2 ersätts med följande text:
"1. Denna artikel skall tillämpas på formgivningstävlingar som anordnas som led i ett förfarande för att tilldela ett kontrakt om tjänster med ett uppskattat värde, exklusive mervärdesskatt, på minst
- det tröskelvärde som avses i artikel 7.1 a första strecksatsen för de tjänster som avses i bilaga I B, tjänsterna i kategori 8 i bilaga I A och telekommunikationstjänsterna i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, eller
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen i för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG, eller
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen ii för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, utom dem som nämns i bilaga I till direktiv 93/36/EEG.
2. Denna artikel skall tillämpas på alla formgivningstävlingar där det sammanlagda beloppet av tävlingspriserna och ersättningarna till deltagarna uppgår till minst
- det tröskelvärde som avses i artikel 7.1 a första strecksatsen för de tjänster som avses i bilaga I B, tjänsterna i kategori 8 i bilaga I A och telekommunikationstjänsterna i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, eller
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen i för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG, eller
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen ii för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, utom dem som nämns i bilaga I till direktiv 93/36/EEG."
4. Artikel 18.2 ersätts med följande text:
"2. Tidsfristen för mottagande av anbud enligt punkt 1 får ersättas av en tidsfrist som är tillräckligt lång för att de berörda parterna skall ha möjlighet att lägga in giltiga anbud, och som i allmänhet inte understiger 36 dagar, men som aldrig är kortare än 22 dagar räknat från dagen för avsändande av meddelandet om upphandling, om de upphandlande myndigheterna har avsänt det preliminära förhandsmeddelande som avses i artikel 15.1, utformat enligt förlagan i bilaga III A (förhandsinformation), till Europeiska gemenskapernas officiella tidning minst 52 dagar och högst tolv månader före insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 15.2, och om det preliminära förhandsmeddelandet dessutom innehåller minst den information som föreskrivs i förlagan i bilaga III B (öppet förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
5. Artikel 19.4 ersätts med följande text:
"4. Tidsfristen för mottagande av anbud enligt punkt 3 får förkortas till 26 dagar om de upphandlande myndigheterna har avsänt det preliminära förhandsmeddelande som avses i artikel 15.1, utformat enligt förlagan i bilaga III A (förhandsinformation), till Europeiska gemenskapernas officiella tidning minst 52 dagar och högst tolv månader före dagen för insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 15.2, och om det preliminära förhandsmeddelandet dessutom innehåller minst den information som föreskrivs i förlagan i bilaga III C (selektivt förfarande) eller, beroende på omständigheterna, i bilaga III D (förhandlat förfarande,) förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
6. I artikel 23 blir den nu befintliga texten punkt 1 och följande punkt läggs till:
"2. Anbud skall avges skriftligen, direkt eller per post. Medlemsstaterna får tillåta avgivande av anbud på alla andra sätt som gör det möjligt att säkerställa
- att varje anbud innehåller de upplysningar som krävs för att utvärdera det,
- att anbudets sekretess består i avvaktan på utvärderingen, och
- om det är nödvändigt av bevisskäl, att anbud så snart som möjligt bekräftas skriftligen eller genom översändande av en bestyrkt kopia,
- att öppnande av anbuden äger rum efter utgången av den tidsfrist som bestäms för avgivande av dessa."
7. Följande artikel förs in:
"Artikel 38a
1. För att möjliggöra bedömning av resultatet av tillämpningen av det här direktivet skall medlemsstaterna till kommissionen sända en statistisk rapport rörande de tjänstekontrakt som under föregående år tilldelats av de upphandlande myndigheterna, senast den 31 oktober 1997 och därefter senast den 31 oktober varje år.
2. Den statistiska rapporten skall innehålla åtminstone följande:
a) När det gäller de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG
- det uppskattade sammanlagda värdet för kontrakt som av varje upphandlande myndighet tilldelas under tröskelvärdet,
- antal och värden för kontrakt som av varje upphandlande myndighet tilldelas över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, tjänstekategori i enlighet med den terminologi som anges i bilaga I och nationalitet för den tjänsteleverantör som tilldelas kontraktet samt, i fråga om förhandlade förfaranden, med uppdelning enligt artikel 11 under angivande av antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
b) När det gäller övriga upphandlande myndigheter som avses med detta direktiv, antal och värden för kontrakt som av varje kategori av upphandlande myndighet tilldelas över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, tjänstekategori i enlighet med den terminologi som anges i bilaga I och nationalitet för den tjänsteleverantör som tilldelas kontraktet samt, i fråga om förhandlade förfaranden, med uppdelning enligt artikel 11 under angivande av antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
c) När det gäller de upphandlande myndigheter som framgår av bilaga I till direktiv 93/36/EEG, antal och sammanlagt värde för kontrakt som tilldelas av varje upphandlande myndighet enligt undantagen från avtalet. När det gäller övriga upphandlande myndigheter som omfattas av detta direktiv, det sammanlagda värdet för kontrakt som tilldelats av varje upphandlande myndighet enligt undantagen från avtalet.
d) Alla andra statistiska upplysningar som skall bestämmas i enlighet med förfarandet i artikel 40.3 och som begärs i enlighet med avtalet.
De statistiska rapporter som begärs enligt denna punkt skall inte avse kontrakt som rör tjänster i kategori 8 i bilaga I A, telekommunikationstjänster i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, eller tjänster i enlighet med bilaga I B, förutsatt att deras uppskattade värde, exklusive mervärdesskatt, är mindre än 200 000 ecu.
3. Kommissionen skall enligt det förfarande som anges i artikel 40.3 bestämma arten av de statistiska upplysningar som krävs enligt det här direktivet."
9. Bilaga III ersätts med den text som framgår av bilaga II till det här direktivet.
Artikel 2
Direktiv 93/36/EEG ändras på följande sätt:
1. I artikel 5
A) ersätts punkt 1 med följande text:
"1. a) Avdelningarna II, III och IV samt artiklarna 6 och 7 skall gälla offentliga varukontrakt som tilldelas av
i) de i artikel 1 b angivna upphandlande myndigheterna, inklusive kontrakt som tilldelas av de upphandlande myndigheterna inom försvarssektorn som anges i bilaga I i den mån det gäller varor som inte omfattas av bilaga II, om det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 200 000 särskilda dragningsrätter (SDR) i ecu,
ii) de upphandlande myndigheterna som anges i bilaga I, om det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 130 000 SDR i ecu. När det gäller upphandlande myndigheter inom försvarssektorn skall detta gälla bara för upphandling av produkter enligt bilaga II.
b) Det här direktivet gäller offentlig upphandling av varor vilkas uppskattade värde är lika med eller högre än det tröskelvärde som gäller vid tidpunkten för offentliggörande av meddelandet enligt artikel 9.2.
c) Motvärdet i ecu och nationella valutor för de tröskelvärden som avses i a skall i princip revideras vartannat år med verkan från och med den 1 januari 1996. Beräkningen av detta motvärde skall grundas på det dagliga genomsnittsvärdet för dessa valutor uttryckt i ecu och för ecun uttryckt i SDR under de sista 24 månaderna fram till den sista augusti som föregår revisionen per den 1 januari.
Den beräkningsmetod som anges i detta stycke skall på förslag av kommissionen ses över av Rådgivande kommittén för offentlig upphandling i princip två år efter det att den tillämpats för första gången.
d) De tröskelvärden som avses i a och deras motvärden uttryckta i ecu och nationella valutor skall regelbundet offentliggöras i Europeiska gemenskapernas officiella tidning i början av november efter den revision som avses i c första stycket."
B) läggs följande punkt till:
"7. De upphandlande myndigheterna skall se till att det inte förekommer någon diskriminering mellan olika leverantörer."
2. Artikel 7.1 och 7.2 ersätts med följande text:
"1. De upphandlande myndigheterna skall inom 15 dagar efter det att en skriftlig begäran inkommit underrätta varje anbudssökande eller anbudsgivare vars ansökan eller anbud har förkastats om orsakerna till att hans ansökan eller anbud förkastats samt underrätta varje anbudsgivare som lämnat ett godtagbart anbud om utformningen av och de relativa fördelarna med det antagna anbudet samt namnet på den anbudsgivare som tilldelats kontraktet.
De upphandlande myndigheterna får emellertid besluta att viss information som rör tilldelningen av kontrakt och som nämns i första stycket inte skall lämnas ut om det bedöms att detta skulle hindra lagarnas tillämpning eller strida mot allmänintresset eller vara till skada för offentliga eller privata företags legitima kommersiella intressen eller för lojal konkurrens mellan tjänsteleverantörer.
2. De upphandlande myndigheterna skall så snart som möjligt underrätta de anbudssökande och anbudsgivarna om de beslut som fattas rörande tilldelningen av kontrakt, inklusive skälen till att de har beslutat att avstå från en upphandling för vilken anbud begärts eller att upprepa förfarandet; dessa upplysningar skall på begäran lämnas skriftligen. Myndigheterna skall även underrätta Byrån för Europeiska gemenskapernas officiella publikationer om dessa beslut."
3. I artikel 10 skall följande punkt föras in:
"1 a. Tidsfristen för mottagande av anbud enligt punkt 1 får ersättas av en tidsfrist som är tillräckligt lång för att de berörda parterna skall ha möjlighet att avge giltiga anbud, och som i allmänhet inte skall understiga 36 dagar, men som aldrig skall vara kortare än 22 dagar räknat från dagen för avsändande av meddelandet om upphandling, om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 9.1, utformat enligt förlagan i bilaga IV A (förhandsinformation) till Europeiska gemenskapernas officiella tidning åtminstone 52 dagar och högst tolv månader före insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 9.2, och om förhandsmeddelandet dessutom innehåller åtminstone den information som föreskrivs i förlagan i bilaga IV B (öppet förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
4. I artikel 11 skall följande punkt föras in:
"3 a. Tidsfristen för mottagande av anbud enligt punkt 3 får förkortas till 26 dagar, om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 9.1, utformat enligt förlagan i bilaga IV A (Förhandsinformation), till Europeiska gemenskapernas officiella tidning åtminstone 52 dagar och högst tolv månader före dagen för insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 9.2, och om förhandsmeddelandet dessutom innehåller åtminstone den information som föreskrivs i förlagan i bilaga IV C (selektivt förfarande) eller, beroende på omständigheterna, i bilaga IV D (förhandlat förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
5. I artikel 15 skall följande punkt läggas till:
"3. Anbud skall avges skriftligen, direkt eller per post. Medlemsstaterna får tillåta avgivande av anbud på alla andra sätt som gör det möjligt att säkerställa
- att varje anbud innehåller de upplysningar som krävs för att utvärdera det,
- att anbudets sekretess består i avvaktan på utvärderingen, och
- om det är nödvändigt av bevisskäl, att anbud så snart som möjligt bekräftas skriftligen eller genom översändande av en bestyrkt kopia,
- att öppnande av anbuden äger rum efter utgången av den tidsfrist som bestäms för avgivande av dessa."
1. Kommissionen skall i samråd med Rådgivande kommittén för offentlig upphandling granska hur detta direktiv tillämpas, och den skall vid behov lägga fram nya förslag för rådet, särskilt i syfte att samordna medlemsstaternas åtgärder för att följa detta direktiv.
2. Kommissionen skall se över detta direktiv och varje ny åtgärd som kan ha tillkommit enligt vad som sägs i punkt 1, med hänsyn till resultaten av de nya förhandlingar som avses i artikel XXIV.7 i avtalet om offentlig upphandling, som ingåtts inom ramen för de multilaterala förhandlingarna i Uruguayrundan (*), nedan kallat "avtalet`, och den skall i förekommande fall lägga fram lämpliga förslag för rådet.
3. Kommissionen skall på grundval av gjorda rättelser, ändringar eller tillägg uppdatera bilaga I i enlighet med det förfarande som anges i artikel 32.2 och skall se till att den offentliggörs i Europeiska gemenskapernas officiella tidning.
1. För att möjliggöra en bedömning av resultatet av tillämpningen av detta direktiv skall medlemsstaterna till kommissionen översända en statistisk rapport rörande de varukontrakt som under det föregående året tilldelats av de upphandlande myndigheterna, senast den 31 oktober 1996, och när det gäller de upphandlande myndigheter som inte anges i bilaga I, senast den 31 oktober 1997 och därefter senast den 31 oktober varje år.
2. Den statistiska rapporten skall innehålla åtminstone följande:
a) När det gäller de upphandlande myndigheter som avses i bilaga I
- det beräknade sammanlagda värdet för kontrakt som av varje upphandlande myndighet tilldelas under tröskelvärdet,
- antal och värden för kontrakt som av varje upphandlande myndighet tilldelas över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, varukategori i enlighet med den terminologi som avses i artikel 9.1 och nationalitet för den varuleverantör som tilldelas kontraktet samt, i fråga om förhandlade förfaranden, med uppdelning enligt artikel 6 med uppgift om antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
b) När det gäller övriga upphandlande myndigheter som omfattas av detta direktiv, antal och värden för kontrakt som tilldelas av varje kategori av upphandlande myndighet över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, varukategori i enlighet med den terminologi som avses i artikel 9.1 och nationalitet för den varuleverantör som tilldelas kontraktet, fördelat enligt artikel 6 med uppgift om antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
c) När det gäller de upphandlande myndigheter som avses i bilaga I, antal och sammanlagt värde för kontrakt som tilldelas av varje upphandlande myndighet enligt undantagen från avtalet. När det gäller övriga upphandlande myndigheter som omfattas av detta direktiv, det sammanlagda värdet för kontrakt som tilldelas av varje kategori av upphandlande myndighet enligt undantagen från avtalet.
d) Alla andra statistiska upplysningar som skall bestämmas i enlighet med förfarandet i artikel 32.2 och som begärs i enlighet med avtalet.
3. Kommissionen skall enligt den förfarande som anges i artikel 32.2 bestämma arten av de statistiska upplysningar som krävs enligt det här direktivet."
8. Bilaga I ersätts med den text som framgår av bilaga I till det här direktivet, och bilaga IV ersätts med den text som framgår av bilaga III till det här direktivet.
Artikel 3
Direktiv 93/37/EEG ändras på följande sätt:
1. I artikel b
A) ersätts punkterna 1 och 2 med följande text:
"1. Det här direktivet gäller för
a) offentliga bygg- och anläggningsarbeten med ett uppskattat värde, exklusive mervärdesskatt, som uppgår till minst 5 000 000 särskilda dragningsrätter (SDR) i ecu.
b) offentliga bygg- och anläggningsarbeten som avses i artikel 2.1 när det uppskattade värdet exklusive mervärdesskatt uppgår till minst 5 000 000 ecu.
2. a) Motvärdet i ecu och nationella valutor för det tröskelvärde som fastställs i punkt 1 skall i princip revideras vartannat år med verkan från den 1 januari 1996. Beräkningen av detta motvärde skall grundas på den genomsnittliga dagskursen för ecun, uttryckt i SDR, och för dessa nationella valutor uttryckt i ecu under de sista 24 månaderna fram till den sista augusti som föregår revisionen per den 1 januari.
Det tröskelvärde som bestäms i punkt 1 och dettas motvärde uttryckt i ecu och i nationella valutor skall offentliggöras i Europeiska gemenskapernas officiella tidning i början av november efter den revision som avses i första stycket.
b) Den beräkningsmetod som anges under a skall på förslag av kommissionen ses över av Rådgivande kommittén för offentlig upphandling i princip två år efter dess första tillämpning."
B) Följande punkt läggs till:
"6. De upphandlande myndigheterna skall se till att det inte förekommer någon diskriminering mellan olika entreprenörer."
2. Artikel 8.1 och 8.2 ersätts med följande text:
"1. De upphandlande myndigheterna skall inom 15 dagar efter det att en skriftlig begäran inkommit underrätta varje anbudssökande eller anbudsgivare vars ansökan eller anbud har förkastats om orsakerna till att hans ansökan eller anbud förkastats samt underrätta varje anbudsgivare som lämnat ett godtagbart anbud om utformningen av och de relativa fördelarna med det antagna anbudet samt namnet på den anbudsgivare som tilldelats kontraktet.
De upphandlande myndigheterna får emellertid besluta att viss information som rör tilldelningen av kontrakt och som nämns i första stycket inte behöver lämnas ut om det bedöms att detta skulle hindra lagarnas tillämpning eller strida mot allmänintresset eller vara till skada för offentliga eller privata företags legitima kommersiella intressen eller för en sund konkurrens mellan entreprenörer.
2. De upphandlande myndigheterna skall så snart som möjligt underrätta de anbudssökande och anbudsgivarna om de beslut som fattats rörande tilldelningen av kontrakt, inklusive skälen till att de har beslutat att avstå från en upphandling för vilken anbud begärts eller att upprepa förfarandet; dessa upplysningar skall på begäran lämnas skriftligen. Myndigheterna skall även underrätta Byrån för Europeiska gemenskapernas officiella publikationer om dessa beslut."
3. Artikel 12.2 ersätts med följande text:
"2. Tidsfristen för mottagande av anbud enligt punkt 1 får ersättas av en tidsfrist som är tillräckligt lång för att de berörda parterna skall ha möjlighet att avge giltiga anbud, och som i allmänhet inte skall understiga 36 dagar, men som aldrig skall vara kortare än 22 dagar räknat från dagen för avsändandet av meddelandet om upphandling om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 11.1, utformat enligt förlagan i bilaga IV A (förhandsinformation), till Europeiska gemenskapernas officiella tidning åtminstone 52 dagar och högst tolv månader före insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 11.2, och om detta meddelande dessutom innehåller minst den information som föreskrivs i förlagan i bilaga IV B (öppet förfarande), förutsatt att denna information var tillgänglig vid tidpunkten för meddelandets offentliggörande."
4. Artikel 13.4 ersätts med följande text:
"4. Tidsfristen för mottagande av anbud enligt punkt 3 får förkortas till 26 dagar, om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 11.1, utformat enligt förlagan i bilaga IV A (Förhandsinformation), till Europeiska gemenskapernas officiella tidning minst 52 dagar och högst tolv månader före dagen för insändandet av det meddelande om upphandling som avses i artikel 11.2, och om förhandsmeddelandet dessutom innehåller minst den information som föreskrivs i förlagan i bilaga IV C (selektivt förfarande) eller, beroende på omständigheterna, i bilaga IV D (förhandlat förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
5. I artikel 18 blir den befintliga texten punkt 1 och följande punkt läggs till:
"2. Anbud skall avges skriftligen, direkt eller per post. Medlemsstaterna får tillåta avgivande av anbud på alla andra sätt som gör det möjligt att säkerställa
- att varje anbud innehåller de upplysningar som krävs för att utvärdera det,
- att anbudets sekretess består i avvaktan på utvärderingen, och
- om det är nödvändigt av bevisskäl, att anbud så snart som möjligt bekräftas skriftligen eller genom översändande av en bestyrkt kopia,
- att öppnande av anbuden äger rum efter utgången av den tidsfrist som gäller för avgivande av dessa."
6. Följande artikel förs in:
"Artikel 33a
"1. För att möjliggöra bedömning av resultatet av tillämpningen av detta direktiv skall medlemsstaterna till kommissionen översända en statistisk rapport rörande de kontrakt för bygg- och anläggningsarbeten som under det föregående året tilldelats av de upphandlande myndigheterna senast den 31 oktober 1997 och därefter senast den 31 oktober varje år.
2. Den statistiska rapporten skall åtminstone innehålla följande:
a) När det gäller de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG
- det beräknade sammanlagda värdet för kontrakt som tilldelats av varje upphandlande myndighet under tröskelvärdet,
- antal och värden för kontrakt som tilldelats av varje upphandlande myndighet över tröskelvärdet, med uppdelning, så långt som möjligt, efter förfarande, kategori av bygg- och anläggningsarbeten i enlighet med den terminologi som används i bilaga II och nationaliteten hos den entreprenör som tilldelats kontraktet samt, i fråga om förhandlande förfaranden, fördelat enligt artikel 7 med uppgift om antal och värden för de kontrakt som tilldelats varje medlemsstat och tredje land.
b) När det gäller de upphandlande myndigheter som omfattas av detta direktiv antal och värde för kontrakt som tilldelats av varje kategori av upphandlande myndigheter över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, kategori av bygg- och anläggningsarbeten i enlighet med den terminologi som används i bilaga II och nationaliteten för det företag som tilldelats kontraktet samt, i fråga om förhandlande förfaranden, med uppdelning enligt artikel 7 med uppgift om antal och värden för de kontrakt som tilldelats varje medlemsstat och tredje land.
c) När det gäller de upphandlande myndigheter som anges i bilaga I till direktiv 93/36/EEG, antal och sammanlagt värde för kontrakt som tilldelats av varje upphandlande myndighet enligt undantagen från avtalet. När det gäller övriga upphandlande myndigheter som avses med detta direktiv, det sammanlagda värdet för kontrakt som tilldelats av varje kategori av upphandlande myndighet enligt undantagen från avtalet.
d) Alla andra statistiska upplysningar som skall bestämmas i enlighet med förfarandet i artikel 35.3 och som begärs i överensstämmelse med avtalet.
3. Kommissionen skall enligt det förfarande som föreskrivs i artikel 35.3 bestämma arten av de statistiska upplysningar som krävs enligt detta direktiv."
8. Bilaga IV ersätts med den text som framgår av bilaga IV till det här direktivet.
Artikel 4
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 13 oktober 1998. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar de bestämmelser som avses i första stycket skall de innehålla en hänvisning till det här direktivet eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som regleras av det här direktivet samt en jämförelsetabell över bestämmelserna i detta direktiv och de antagna nationella bestämmelserna.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EG) nr 142/97 av den 27 januari 1997 om lämnande av uppgifter om vissa existerande ämnen i enlighet med rådets förordning (EEG) nr 793/93 (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 793/93 av den 23 mars 1993 om bedömning och kontroll av risker med existerande ämnen (1), särskilt artikel 12.2 i denna, och med beaktande av följande:
Kommissionen har behov av relevanta uppgifter om vissa ämnen för att kunna inleda de förfaranden för översyn som avses i artiklarna 69, 84 och 112 i anslutningsfördraget för bestämmelser som ännu inte tillämpas i de nya medlemsstaterna. Dessa upplysningar måste finnas tillgängliga innan alla de upplysningar som avses i artiklarna 3 och 4 i förordning (EEG) nr 793/93 finns att tillgå.
I artikel 12 föreskrivs att tillverkare eller importörer av vissa ämnen som kan utgöra en allvarlig risk för människor eller miljön, kan åläggas att lämna de uppgifter som de har tillgång till.
Med beaktande av kommissionens förordning (EEG) nr 1488/94 (2) om principer för bedömning av risker för människor och miljö av existerande ämnen i enlighet med förordning (EEG) nr 793/93.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som inrättats i enlighet med artikel 15 i förordning (EEG) nr 793/93.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De som tillverkar eller importerar ämnen som ingår i förteckningen i bilagan till denna förordning skall inom fyra månader efter det att förordningen träder i kraft till kommissionen lämna all relevant tillgänglig information om exponering av människor eller miljö för dessa ämnen.
Relevant information om exponering av människor eller miljön för ett ämne omfattar utsläpp av ämnet eller exponering av människor eller delar av miljön för ämnet under olika stadier av ämnets livscykel i enlighet med artikel 3.3 och bilaga 1 A till förordning (EG) nr 1488/94, där
- människor avser arbetstagare, konsumenter och andra som kommer i kontakt med ämnet via miljön,
- delar av miljön omfattar vatten, mark och luft, vilket också innefattar information om ämnets fördelning och omvandling i reningsverk och dess ackumulering i näringskedjan och
- ett ämnes livscykel omfattar tillverkning, transport, lagring, blandning till en beredning eller annan bearbetning, användning och bortskaffade eller återvinning.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
RÅDETS FÖRORDNING (EG) nr 552/97 av den 24 mars 1997 om tillfälligt upphävande av allmänna tullförmåner för Unionen Myanmar
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 3281/94 av den 19 december 1994 om tillämpning av ett fyraårigt system med allmänna tullförmåner (1995-1998) för vissa industriprodukter med ursprung i utvecklingsländerna (1), särskilt artikel 12.3 i denna,
med beaktande av rådets förordning (EG) nr 1256/96 av den 20 juni 1996 om tillämpningen av en flerårig ordning med allmänna tullförmåner under perioden 1 juli 1996-30 juni 1999 för vissa jordbruksprodukter med ursprung i utvecklingsländerna (2), särskilt artikel 12.3 i denna,
med beaktande av kommissionens förslag (3),
med beaktande av Europaparlamentets yttrande (4),
med beaktande av Ekonomiska och sociala kommitténs yttrande (5), och
med beaktande av följande: Enligt förordning (EG) nr 3281/94 och förordning (EG) nr 1256/96 omfattas Unionen Myanmar (nedan kallad Myanmar) av allmänna tullförmåner.
Enligt artikel 9 i förordning (EG) nr 3281/94 och artikel 9 i förordning (EG) nr 1256/96 kan förmånerna i fråga helt eller delvis tillfälligt upphävas under omständigheter som inbegriper utövande av någon form av tvångsarbete såsom det definieras i Genèvekonventionerna av den 25 september 1926 och den 7 september 1956 och i Internationella arbetsorganisationens (ILO) konventioner nr 29 och 105.
Den 7 juni 1995 ingav Fria fackföreningsinternationalen (ICFTU) och Europeiska fackliga samorganisationen (ETUC) ett gemensamt klagomål enligt artikel 9 i förordning (EG) nr 3281/94 till kommissionen och begärde ett tillfälligt upphävande av gemenskapens system med allmänna tullförmåner för Myanmar på grund av dess användning av tvångsarbete.
Den 2 januari 1997 anmälde ICFTU och ETUC till kommissionen att de utvidgade omfattningen av det gemensamma klagomål som de ingivit enligt förordning (EG) nr 3281/94 i syfte att det tillfälliga upphävandet av gemenskapens system med förmåner för Myanmar även görs enligt förordning (EG) nr 1256/96.
Kommissionen har i samråd med kommittén för förvaltningen av allmänna tullförmåner undersökt klagomålet av den 7 juni 1995 och de fakta som de klagande framlagt har bedömts vara tillräckliga för att inleda en undersökning. Kommissionen fattade beslut om detta i ett tillkännagivande av den 16 januari 1996 (6).
Myanmars myndigheter har officiellt underrättats om att undersökningen har inletts. De bestrider att de metoder som avses i klagomålet utgör tvångsarbete med hänvisning till de undantag som avses i artikel 2.2 i ILO:s konvention nr 29 och hävdar att dessa undantag omfattas av 1907 års Town Act och 1908 års Village Act enligt vilka det är tillåtet att ålägga befolkningen att utföra arbeten och tjänster. ILO bestrider denna tolkning och dess behöriga organ har begärt att lagarna i fråga snarast skall upphävas i syfte att göra dessa lagar förenliga med andan och ordalydelsen i konvention nr 29.
De skriftliga och muntliga uppgifter som kommissionen har inhämtat i samband med undersökningen som genomfördes i samråd med kommittén för förvaltningen av allmänna tullförmåner stödjer de påståenden som anges i klagomålet. Det framgår att myndigheterna i Myanmar rutinmässigt med tillgripande av tvång och upprepade våldsamma straffåtgärder har tillämpat tvångsarbete inte endast för militära operationer utan även för civila och militära infrastrukturbyggprojekt.
Kommissionen har, i syfte att komplettera de uppgifter som den har inhämtat i samband med undersökningen, uppmanat myndigheterna i Myanmar att samarbeta genom att tillåta en undersökningsdelegation inresa i landet. Myndigheterna i Myanmar har inte efterkommit denna uppmaning och eftersom villkoren i artikel 11.5 i förordning (EG) nr 3281/94 följaktligen är uppfyllda kan slutsatserna grundas på tillgängliga uppgifter.
All den bevisning som kommissionen har inhämtat i den undersökning som den har utfört efter ICFTU:s och ETUC:s ursprungliga klagomål samt de slutsatser som den har dragit på grundval av dessa uppgifter är tillräckligt omfattande för att utgöra ett välgrundat underlag för prövningen av det utvidgade klagomål som har inlämnats av dessa organisationer den 2 januari 1997. Detta gör det onödigt med en särskild undersökning för jordbrukssektorn. Kraven i artikel 9.2 i förordning (EG) nr 1256/96 är sålunda uppfyllda och villkoren i artikel 11.5 i den förordningen är uppfyllda.
Av de tillgängliga uppgifterna framgår alltså att det finns tillräckliga skäl att dra slutsatsen att ett upphävande av systemet med allmänna tullförmåner som har beviljats Myanmar är berättigat.
En rapport om undersökningens slutsatser har överlämnats till kommittén för förvaltningen av allmänna tullförmåner enligt artikel 12.1 i förordning (EG) nr 3281/94.
Det faktum att de fördömda metoderna varit rutinmässiga och omfattande gör att det är befogat att helt upphäva bestämmelserna.
Mot bakgrund av detta bör tillämpningen av allmänna tullförmåner för industriprodukter och jordbruksprodukter med ursprung i Myanmar tillfälligt upphävas till dess det fastställts att metoderna i fråga har upphört.
Varor som redan avsänts till Europeiska gemenskapen bör undantas från detta upphävande av förmåner under förutsättning att de avsänts före den dag när denna förordning träder i kraft.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De allmänna tullförmåner enligt förordning (EG) nr 3281/94 och förordning (EG) nr 1256/96 är härmed tillfälligt upphävda för Unionen Myanmar.
Artikel 2
Rådet skall, med kvalificerad majoritet, på förslag av kommissionen, låta upphäva tillämpningen av denna förordning då det på grundval av en rapport om tvångsarbete i Myanmar från kommissionen kan visas att de metoder som avses i artikel 9.1 första strecksatsen i förordning (EG) nr 3281/94 och artikel 9.1 första strecksatsen i förordning (EG) nr 1256/96 som har orsakat upphävandet av allmänna tullförmåner för Myanmar inte längre förekommer.
Artikel 3
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 659/97 av den 16 april 1997 om tillämpningsföreskrifter för förordning (EG) nr 2200/96 med avseende på interventionsordningen för frukt och grönsaker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker (1), särskilt artiklarna 30.6, 48 och 57 i denna, och
med beaktande av följande: I avdelning IV i förordning (EG) nr 2200/96 fastställs interventionsordningen för de produkter som avses i artikel 1.2 i denna. Tillämpningsföreskrifter till dessa bestämmelser bör därför fastställas.
Vad gäller produkter bör uttrycken "inte saluförts" och "återtagits från marknaden" likställas och ingå i samma definition. Det är också lämpligt att förtydliga att för produkter som återtas från marknaden behöver förpackningskraven inte vara uppfyllda.
Det är nödvändigt att fastställa regleringsår för de produkter som anges i bilaga II till förordning (EG) nr 2200/96.
För att tillämpa de begränsningar som föreskrivs i artiklarna 23 och 24 i förordning (EG) nr 2200/96 är det lämpligt att definiera den "saluförda kvantiteten" av en produkt som saluförs en producentorganisation med hänsyn till den faktiska produktion som producentorganisationen i fråga är upphov till, produktionen från andra producentorganisationer liksom produktionen från producenter som inte är anslutna till någon producentorganisation.
I artikel 28 i förordning (EG) nr 2200/96 förskrivs att medlemsstaterna måste meddela de priser som noteras på de representativa marknaderna för vissa bestämda produkter och för vissa perioder. Följaktligen bör en förteckning upprättas över dessa marknader och över berörda produkter.
I artikel 26 i förordning (EG) nr 2200/96 fastställs gemenskapskompensationen för återtagande av de produkter som anges i bilaga II till den förordningen. Det är lämpligt att föreskriva ett system för utbetalning för att på så sätt hela tiden iaktta de begränsningar som föreskrivs i artikel 23 i förordning (EG) nr 2200/96.
För att undvika oriktigheter vid tillämpningen av ordningen och garantera öppenhet och insyn bör producentorganisationerna i förväg meddela varje återtagande till kontrollmyndigheterna. Om ett sådant meddelande inte har lämnats får produkten avsättas först efter tillstånd från medlemsstaten. Dessutom måste ett kommunikationssystem inrättas, både för producentorganisationerna och för medlemsstaterna.
Det är lämpligt att fastställa, i enlighet med vad som förskrivs i artikel 25 i förordning (EG) nr 2200/96, de frister för att framlägga de åtgärder som medlemsstaterna vidtar för att skydda miljön vid återtagande.
I artikel 30.1 a första andra och tredje strecksatsen i ovannämnda förordning föreskrivs att frukt och grönsaker som återtas från marknaden i enlighet med artikel 23.1 i den förordningen och som förblivit osålda, får delas ut gratis, både inom gemenskapen och utom gemenskapen, som humanitärt bistånd till vissa nödlidande befolkningskategorier med hjälp av välgörenhetsorganisationer. Det är i detta syfte lämpligt att föreskriva att dessa välgörenhetsorganisationer skall godkännas på förhand.
Bestämmelserna i kommissionens förordning (EEG) nr 3587/86 (3), senast ändrad genom förordning (EG) nr 1363/95 (4), (EEG) nr 827/90 (5), senast ändrad genom förordning (EG) nr 771/95 (6), (EEG) nr 2103/90 (7), ändrad genom förordning (EG) nr 1363/95, (EEG) nr 2276/92 (8), senast ändrad genom förordning (EG) nr 1363/95 och (EG) nr 113/97 (9), som har blivit föråldrade eller som skall ersättas av bestämmelserna i denna förordning, bör upphöra att gälla.
De bestämmelser som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för frukt och grönsaker samt från Kommittén för den europeiska utvecklings- och garantifonden för jordbruket.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I denna förordning fastställs tillämpningsföreskrifter för interventionsordning som avses i avdelningen IV i förordning (EG) nr 2200/96, och gäller för de produkter som avses i artikel 1.2 i den förordningen.
Artikel 2
1. Med produkter som "återtagits från marknaden" eller produkter som "inte saluförts" avses enligt denna förordning sådana produkter som inte sålts genom en producentorganisation, i enlighet med den interventionsordning som avses i förordning (EG) nr 2200/96.
2. Produkterna som återtagits från marknaden bör överensstämma med gällande normer om sådana normer har fastställts i enlighet med artikel 2 i förordning (EG) nr 2200/96. I detta fall är dock normerna för förpackning inte tillämpliga.
Artikel 3
1. För varje produkt skall den av en producentorganisation "saluförda kvantitet" som nämns i artikel 23.3 i förordning (EG) nr 2200/96 vara summan av
a) medlemmarnas produktion som faktiskt sålts genom eller bearbetats av producentorganisationen,
b) den produktion som medlemmarna i producentorganisationen sålde direkt enligt de villkor som avses i artikel 11.1 c 3 första och fjärde strecksatsen i förordning (EG) nr 2200/96,
c) den produktion som framställts av medlemmar i andra producentorganisationer och som saluförts genom den berörda producentorganisationen i enlighet med artikel 11.1 c 3 andra och tredje strecksatsen i förordning (EG) nr 2200/96.
Den saluförda kvantitet som avses i första stycket omfattar inte den produktion som saluförts av de av producentorganisationens medlemmar som får sälja i enlighet med artikel 11.1 c.3 andra och tredje strecksatsen i förordning (EG) nr 2200/96.
2. Den saluförda produktion som avses i artikel 23.4 i förordning (EG) nr 2200/96 skall likställas med den saluförda kvantiteten definierad enligt punkt 1.
Artikel 4
Regleringsåren för produkter som omfattas av gemenskapskompensation för återtagande i enlighet med artikel 23.3 i förordning (EG) nr 2200/96 anges i bilaga I till denna förordning.
Regleringsåren för produkter som avses i artikel 1.2 i förordning (EG) nr 2200/96 andra än de som avses i första stycket, sträcker sig från den 1 januari till den 31 december.
Artikel 5
2. Ansökan som avses i punkt 1 skall minst gälla en period om en månad. Den skall åtföljas av dokument som intygar kvantiteten av varje saluförd produkt och kvantiteten av varje produkt som inte saluförts genom producentorganisationen samt innehåller detaljerade uppgifter om
a) medlemmarnas produktion som faktiskt sålts genom eller bearbetats av producentorganisationen,
b) den produktion som medlemmarna i andra producentorganisationer salufört genom den berörda producentorganisationen i enlighet med artikel 11.1 c 3 andra och tredje strecksatsen i förordning (EG) nr 2200/96,
c) den produktion som tillförts av var och en av de odlare som inte tillhör någon producentorganisation enligt villkoren i artikel 24 i förordning (EG) nr 2200/96.
3. Vid behandlingen av varje ansökan skall medlemsstaterna för de sammanlagda kvantiteter som inte saluförts efter inledningen av varje regleringsår i fråga kontrollera att de begränsningar som föreskrivs i artiklarna 23 och 24 i förordning (EG) nr 2200/96 efterlevs. Om ett överskridande sker skall gemenskapskompensation för återtagande endast utgå under förutsättning att dessa begränsningar respekteras med hänsyn till den kompensation som redan utgått. De överskridande kvantiteterna skall återtas vid behandlingen av nästa ansökan.
Artikel 6
Utan att det påverkar tillämpningen av artikel 22 i denna förordning när det gäller utbetalning av kompensation för återtagande av produkter som inte anges i bilaga II till förordning (EG) nr 2200/96 samt utbetalning av det tillägg till gemenskapens ersättning för återtagande som föreskrivs i artikel 15.3 a och 15.3 b i förordning (EG) nr 2200/96, skall bestämmelserna i förordning (EG) nr 411/97 tillämpas.
Artikel 7
1. De representativa marknader som avses i artikel 28.1 i förordning (EG) nr 2200/96 skall motsvaras av dem som anges i bilaga II till denna förordning.
2. Medlemsstaterna skall en gång i veckan på elektronisk väg meddela kommissionen de på de representativa marknaderna för varje marknadsdag noterade dagspriserna för de produkter och för de perioder som anges i bilaga III till denna förordning. Kommissionen skall vidarebefordra dessa upplysningar till medlemsstaterna.
Artikel 8
1. Producentorganisationerna eller deras sammanslutningar skall minst 24 timmar i förväg underrätta de behöriga nationella myndigheterna om varje återtagande samt tillhandahålla en detaljerad förteckning över de produkter som avses för intervention, den kvantitet som beräknas för varje produkt.
2. Följande uppgifter skall av producentorganisationerna eller deras sammanslutningar meddelas till medlemsstaterna, vilka i sin tur skall vidarebefordra dem till kommissionen:
a) De tillgängliga lagren av äpplen och päron den första dagen i varje månad.
b) Vid början av varje regleringsår uppgifterna om de uppodlade arealerna för varje produkt och eventuellt för varje sort.
Artikel 9
1. Före den 10 i varje månad skall medlemsstaterna på elektronisk väg till kommissionen översända en uppskattning fördelad per produkt av de produkter som inte saluförts under föregående månad.
2. Vid slutet av varje regleringsår skall medlemsstaterna för varje berörd produkt meddela kommissionen de uppgifter som anges i bilaga IV. Dessa uppgifter skall meddelas
a) senast den 30 juni som följer på varje regleringsår för tomater, auberginer, blomkål, aprikoser, persikor, nektariner, vindruvor, meloner och vattenmeloner samt för produkter utanför bilaga II till förordning (EG) nr 2200/96, och
b) senast den 30 november som följer på varje regleringsår för citroner, päron, äpplen, satsumas, clementiner och söta apelsiner.
3. Om medlemsstaterna inte lämnar in de uppgifter som avses i punkt 2 och om de meddelade uppgifterna med hänsyn till de objektiva fakta som kommissionen förfogar över verkar oriktiga, kan kommissionen i avvaktan på att ovan nämnda uppgifter läggs fram tillfälligt upphöra med den utbetalning av förskotten på de beräknade utgifter som avses i artikel 5.2 a i rådets förordning (EEG) nr 729/70 (10).
Artikel 10
Artikel 11
1. De produkter som återtagits från marknaden under ett visst regleringsår får ställas till förfogande för välgörenhetsorganisationer som godkänts av medlemsstaterna på deras begäran för gratis utdelning i enlighet med bestämmelserna i artikel 30.1 a första och tredje strecksatsen i förordning (EG) nr 2200/96.
2. För att kunna bli godkända skall välgörenhetsorganisationerna förbinda sig att
a) följa bestämmelserna i denna förordning,
b) föra särskilda räkenskaper över den aktuella verksamheten,
c) underkasta sig de kontroller som föreskrivs av gemenskapsrätten.
3. Medlemsstaterna skall godkänna välgörenhetsorganisationer i minst en av följande kategorier:
a) Välgörenhetsorganisationer som har tillstånd att genomföra utdelning på medlemsstatens territorium av produkter som har återtagits från marknaden.
Medlemsstaterna skall till kommissionen lämna in förteckningar över de godkända välgörenhetsorganisationer som avses i första stycket b och c och kommissionen skall i sin tur se till att de offentliggörs i Europeiska gemenskapernas officiella tidning, serie C.
Artikel 12
De av medlemsstaterna utvalda institutioner som avses i artikel 30.1 a andra strecksatsen i förordning (EG) nr 2200/96 måste uppfylla villkoren i artikel 11.2 i denna förordning.
Artikel 13
Medlemsstaterna skall vidta nödvändiga åtgärder för att underlätta kontakter och transaktioner mellan de berörda producentorganisationerna och de välgörenhetsorganisationer som godkänts i enlighet med artikel 11.2.
Vid slutet av varje regleringsår skall medlemsstaterna till kommissionen vidarebefordra de uppgifter om gratis utdelning som avses i bilaga VI.
Artikel 14
1. Gratis utdelning som sker utanför gemenskapen inom ramen för humanitärt bistånd skall genomföras av sådana välgörenhetsorganisationer som avses i artikel 11.3 c, enligt punkterna 2 och 3 i denna artikel.
2. För avsända produkter utgår inget exportbidrag. På tulldokumentet för export, transiteringshandlingen samt det kontrolldokument T 5 som eventuellt utfärdats skall uppgiften "utan bidrag" anges.
Artikel 15
1. Transportkostnader knutna till insatser för gratis utdelning av alla produkter som återtagits från marknaden skall betalas av garantisektionen inom Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) på grundval av schablonbelopp som fastställs utifrån avståndet mellan platsen för återtagandet och leveransplatsen och som anges i bilaga V.
Om gratis utdelning sker utanför gemenskapen skall schablonbeloppen som avses i bilaga V täcka avståndet mellan platsen för återtagandet och den plats där sändningen lämnar gemenskapen.
2. Transportkostnaderna skall betalas till den avsändare som faktiskt har burit transportkostnaderna i fråga.
Utbetalningen av beloppen skall ske på villkor att intyg läggs fram som bekräftar
- namnet på de mottagande organisationerna,
- kvantiteten av aktuella produkter,
- ett övertagandeintyg utfärdat av välgörenhetsorganisationen,
- vilka transportmedel som använts.
Artikel 16
1. När det gäller återtagna äpplen och citrusfrukter skall sorterings- och förpackningskostnader i samband med gratis utdelning betalas av garantisektionen inom EUGFJ och inom gränsen för de belopp som anges i bilaga V.2, om det rör sig om gratis utdelning inom ramen för ett avtal mellan de berörda producent- och välgörenhetsorganisationerna.
2. Enligt punkt 1 skall producentorganisationerna vid regleringsårets början ingå avtal med de välgörenhetsorganisationer som godkänts i enlighet med artikel 11.2 och 11.3 samt underrätta de behöriga nationella myndigheterna om dessa avtal så snart de ingåtts. Dessa myndigheter får fastställa en frist för slutandet av sådana avtal.
3. Dessa avtal får slutas på villkor att det finns produkter som återtagits från marknaden. Kvantiteterna som anges i avtalen får med hänsyn till situationen på marknaden ökas under regleringsåret.
4. Avtalen skall slutas för ett enda regleringsår i den mening som avses i förordning (EG) nr 2200/96 och skall innehålla uppgifter om
- den för varje produkt sannolika utdelningskvantiteten,
- de planerade transportmedlen,
- den planerade leveranstakten,
- den överenskomna överlåtelseplatsen,
- kravet att producentorganisationen tillhandahåller produkter som storlekssorterats på förhand och förpackats i emballage med en vikt på högst 25 kg.
- en uppskattning av antalet stödmottagare per administrativ enhet.
5. Medlemsstaterna skall senast en månad efter det att avtalen slutits meddela kommissionen de uppgifter som avses i punkt 4.
6. Ersättning för sorterings- och förpackningskostnader skall utbetalas till de producentorganisationer som har sorterat och förpackat produkterna och skall utgå på villkor att intyg läggs fram som bekräftar
- namnet på de mottagande organisationerna,
- kvantiteten berörda produkter,
- de faktiska kostnaderna för förpackning och sortering,
- ett övertagandeintyg som utfärdats av välgörenhetsorganisationen.
Artikel 17
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att säkerställa att bestämmelserna i avdelning IV i förordning 2200/96 efterlevs, särskilt de som föreskrivs i punkterna 2, 3 och 4.
2. Medlemsstaterna skall minst en gång per regleringsår genomföra fysiska kontroller och dokumentkontroller av alla producentorganisationernas återtagande transaktioner. Dessa kontroller skall för varje produkt gälla minst 20 % av den totala återtagna kvantiteten.
De skall dessutom förvissa sig om att de produkter som inte saluförts överensstämmer med gällande normer, om sådana normer har fastställts med tillämpning av artikel 2.2 i förordning (EG) nr 2200/96.
Vid tillämpning av artikel 30.2 i förordning (EG) nr 2200/96, skall medlemsstaterna kontrollera alla återtagna kvantiteter.
3. Medlemsstaterna skall genomföra dokumentkontroller av interventionerna för att effektivt fastställa att redovisningen utförs på ett korrekt sätt samt att betalningsvillkoren uppfylls för gemenskapskompensation för återtagande eller om finansiering genom driftsfonden, som avses i artikel 15.1 i förordning (EG) nr 2200/96.
Kontrollerna skall genomföras för varje producentorganisation minst en gång per regleringsår och den skall för varje produkt omfatta minst 10 % av betalningsansökningarna.
4. Om kontrollerna visar på väsentliga oriktigheter skall de behöriga myndigheterna genomföra ytterligare kontroller det pågående regleringsåret och öka antalet kontroller det påföljande regleringsåret.
Artikel 18
a) att verksamheten i fråga utförs på ett korrekt sätt,
b) välgörenhetsorganisationernas slutliga användning av produkterna, särskilt genom att kräva av dessa ett övertagandeintyg som intygar användningen av produkterna, och
c) produkternas slutliga bestämmelseort.
2. Kontrollen enligt punkt 1 består av dokumentkontroller och fysiska kontroller, vilka skall avse berörda producentorganisationer och välgörenhetsorganisationer. Kontrollerna får bestå av stickprovskontroller som genomförs varje regleringsår och de skall avse minst 10 % av de utdelade kvantiteterna.
3. Beträffande utdelning inom gemenskapen och utan att det påverkar bestämmelserna i artikel 39 i förordning (EG) nr 2200/96 skall de behöriga nationella myndigheterna genomföra kontroller av produkternas användning och slutliga bestämmelse på det territorium där gratisutdelningen sker.
4. På begäran av medlemsstaten skall kommissionen bistå medlemsstaten vid kontrollen av de gratisutdelningar som genomförs utanför gemenskapen.
Artikel 19
1. Den som mottar gemenskapernas kompensation för återtagande eller finansiering genom driftsfonden är skyldig att återbetala dubbelt så mycket som de belopp som felaktigt betalats ut plus ränta för den tid som förflutit mellan utbetalningen och mottagarens återbetalning om det vid kontroll enligt artikel 17 visar sig att
a) de produkter som inte saluförts inte överensstämmer med de normer som avses i artikel 2 i förordning (EG) nr 2200/96,
b) de produkter som inte saluförts inte har avsatts i enlighet med artikel 30 i förordning (EG) nr 2200/96,
c) avsättningen av produkter som inte saluförts medför allvarliga skador för miljön.
2. De återtagna beloppen samt räntan skall betalas till den behöriga utbetalande organisationen och avräknas de kostnader som finansieras av EUGFJ.
3. I händelse av uppsåtlig falskdeklaration eller av grov vårdslöshet skall den berörda producentorganisationen inte erhålla gemenskapskompensation för återtagande under det regleringsår för vilket oegentligheten konstaterats.
Artikel 20
1. Om det vid kontroller i enlighet med artikel 18 konstateras oegentligheter som kan tillskrivas producentorganisationer godkända välgörenhetsorganisationer eller institutionerna som avses i artiklarna 11 och 12 skall bestämmelserna i punkt 2-7 i denna artikel tillämpas.
2. Godkännandet av den välgörenhetsorganisation som avses i artikel 11.2 dras in. Indragningen skall verkställas omedelbart, den skall gälla under minst ett regleringsår samt förlängas med hänsyn till hur allvarlig oegentligheten är.
3. De institutioner som anges i artikel 12 har inte rätt till gratis utdelning under nästa regleringsår.
4. Välgörenhetsorganisationen eller den institution som tagit emot produkten som återtagits från marknaden skall återbetala värdet av de produkter som ställts till dess förfogande ökat med en ränta beräknad på grundval av den tid som förflutit mellan mottagandet av produkten och mottagarens återbetalning.
Den avsändare som har fått transportkostnaderna täckta som avses i artikel 15 skall återbetala den dubbla summan av de belopp som erhållits för transportkostnader, ökad med en ränta beräknad på grundval av den tid som förflutit mellan utbetalningen och mottagarens återbetalning.
6. Räntesatsen för denna ränta skall vara den som tillämpas av Europeiska monetära institutet för dess transaktioner i ecu som offentliggörs i Europeiska gemenskapernas officiella tidning C-serien, och som gäller den dag den felaktiga utbetalningen gjordes, ökad med tre procentenheter.
7. De återtagna beloppen samt räntan skall betalas till det behöriga utbetalande organet och avräknas från de utgifter som finansieras av EUGFJ.
Artikel 21
Artikel 22
De producentorganisationer som ansökt om godkännande av ett operativt program i enlighet med artiklarna 3 eller 15 i förordning (EG) nr 411/97 får som en tillfällig åtgärd för 1997 på egen risk och i enlighet med artikel 15.3 b i förordning (EG) nr 2200/96 bevilja ett tillägg till gemenskapens ersättning för återtagande.
Artikel 23
Förordningarna (EEG) nr 3587/86, (EEG) nr 827/90, (EEG) nr 2103/90, (EEG) nr 2276/92 samt (EG) nr 113/97 upphör att gälla.
Artikel 24
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 888/97 av den 16 maj 1997 om ändring av vissa bestämmelser i de normer som fastställts för färsk frukt och färska grönsaker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker (1), särskilt artiklarna 2.2 och 10 i denna, och
med beaktande av följande: I artikel 2 i förordning (EG) nr 2200/96 fastställs att kommissionen, när den antar normer för färsk frukt och färska grönsaker, skall beakta Ekonomiska kommissionens för Europa (FN) internationella normer.
Gemenskapens normer för frukt och grönsaker är utspridda på en rad gemenskapsbestämmelser. Det är nödvändigt att harmonisera vissa av dessa bestämmelser för att uppnå en enhetlig tillämpning av dessa normer och av kontrollen av deras överensstämmelse.
I Ekonomiska kommissionens för Europa internationella normer för färsk frukt och färska grönsaker fastställs tydligt hur packaren och avsändaren skall anges på förpackningen. Dessa internationella bestämmelser bör, i synnerhet för den juridiska tydlighetens skull, införlivas i gemenskapens alla normer för färsk frukt och färska grönsaker.
De förordningar i vilka normer för kronärtskockor, bönor, ärtor, blomkål och vitlök föreskrivs innehåller inga bestämmelser om angivelse av ursprungsland på förpackningen. Bestämmelser av denna art i gällande internationella normer bör införas i dessa förordningar.
En kategori III har fastställts i de förordningar i vilka normer för purjolök, aubergine, zucchini, tomater, lök, endiver, körsbär, jordgubbar, brysselkål, bordsdruvor, trädgårdssallad, endivsallad, gurkor, citrusfrukter, äpplen och päron har fastställts. Denna kategori III tillämpades enbart i undantagsfall och har förlorat sin betydelse för färsk frukt och färska grönsaker. De internationella normerna innehåller ingen sådan kategori och för enkelhetens skull bör den tas bort i gemenskapens normer.
I rådets förordning nr 211/66/EEG av den 14 december 1966 om utökning av de gemensamma kvalitetsnormerna för vissa frukt och grönsaksslag med en kompletterande kvalitetsklass (2), senast ändrad genom kommissionens förordning (EEG) nr 3596/90 (3), fastställs också en kategori III för blomkål. Av samma skäl som ovan bör förordning nr 211/66/EEG upphävas.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för frukt och grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) i de förordningar som anges i bilaga I skall ändras på följande sätt:
Texten i A "Identifiering" skall ersättas med följande:
"Packare och/eller avsändare. Namn och adress eller officiellt utfärdat eller godkänt märke. Om en kod (ett märke) används skall "packare och/eller avsändare (eller motsvarande förkortning)" anges vid denna kod (detta märke)."
b) i de förordningar som anges i bilaga II skall ändras på följande sätt:
Texten i C "Produktens ursprung" skall ersättas med följande:
"Ursprungsland och eventuellt produktionsområde eller nationell, regional eller lokal benämning."
2. I de förordningar som anges i bilaga III skall all hänvisning till kategori III utgå.
3. Förordning nr 211/66/EEG skall upphöra att gälla.
Artikel 2
Denna förordning träder i kraft den 1 juli 1997.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 1054/97 av den 11 juni 1997 om klassificeringen av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 866/97 (2), särskilt artikel 9 i denna, och med beaktande av följande:
För att åstadkomma en enhetlig tillämpning av den Kombinerade nomenklatur som intagits i bilagan till ovannämnda förordning bör bestämmelser antas avseende klassificering av de varor som intagits i bilagan till den här förordningen.
De allmänna reglerna för hur Kombinerade nomenklaturen skall tolkas har fastställts i förordning (EEG) nr 2658/87. Dessa regler skall också tillämpas på all annan nomenklatur som baseras på denna, även om detta gäller endast delvis eller om underuppdelningar eventuellt gjorts som tillägg till den, och som fastställts genom särskilda gemenskapsbestämmelser för tillämpningen av tullmässiga eller andra åtgärder inom ramen för varuutbytet.
Med tillämpning av dessa allmänna regler måste de varor som beskrivs i första kolumnen i tabellen i bilagan till den här förordningen hänföras till de nummer i Kombinerade nomenklaturen som anges i andra kolumnen med stöd av den motivering som anges i tredje kolumnen.
Om inte annat följer av gällande bestämmelser i gemenskapen avseende systemet för dubbelkontroll samt övervakning på gemenskapsnivå, i förväg eller i efterhand, av textilvaror som importeras till gemenskapen, är det lämpligt att bindande tulltaxeupplysningar i fråga om klassificering av varor i Kombinerade nomenklaturen som lämnats av tullmyndigheterna i medlemsstaterna och som inte överensstämmer med den här förordningen får fortsätta att åberopas av innehavaren under en period av 60 dagar, i enlighet med bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen (3), senast ändrad genom förordning (EG) nr 82/97 (4).
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från sektionen för tulltaxe- och statistiknomenklatur inom tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i första kolumnen i tabellen i bilagan hänförs till de nummer i Kombinerade nomenklaturen som anges i andra kolumnen i samma tabell.
Artikel 2
Om inte annat följer av gällande bestämmelser i gemenskapen avseende systemen för dubbelkontroll samt övervakning på gemenskapsnivå, i förväg eller i efterhand, av textilvaror som importeras till gemenskapen får bindande tulltaxeupplysningar i fråga om klassificering av varor i Kombinerade nomenklaturen, som lämnats av tullmyndigheterna i medlemsstaterna och som inte överensstämmer med den här förordningen, fortsätta att åberopas, i enlighet med bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 under en period av 60 dagar.
Artikel 3
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1059/97 av den 11 juni 1997 om anpassning av den årliga maximala fiskeansträngningsnivån för vissa fiskevatten
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2027/95 av den 15 juni 1995 om en förvaltningsordning för fiskeansträngningen för vissa fiskezoner och fisketillgångar inom gemenskapen (1), särskilt artikel 4 andra strecksatsen i denna, och
med beaktande av följande: I artikel 4 andra strecksatsen i förordning (EG) nr 2027/95 föreskrivs att kommissionen på en medlemsstats begäran skall vidta lämpliga åtgärder så att denna medlemsstat skall kunna utnyttja sina kvoter i enlighet med bestämmelserna i artikel 6.2 tredje stycket i rådets förordning (EG) nr 685/95 av den 27 mars 1995 om administreringen av fiskeinsatsen med avseende på vissa fiskezoner och -resurser i gemenskapen (2).
Nederländerna har begärt att kommissionen skall anpassa den årliga maximala fiskeansträngningsnivå som beviljats den nederländska flottan för vissa kvoter som de har tilldelats i enlighet med rådets förordning (EG) nr 390/97 av den 20 december 1996 om fastställande, för vissa fiskbestånd och grupper av fiskbestånd, av totala tillåtna fångstmängder under 1997 och av vissa villkor för fångsten (3), senast ändrad genom förordning (EG) nr 711/97 (4).
Med beaktande av rådets förordning, skall följande träda i kraft omedelbart så att Nederländerna kan använda sin tilldelade kvot.
Förvaltningskommittén för fiskeresurser har avgivit sitt yttrande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Den årliga maximala fiskeansträngningsnivån för Nederländerna för fiske med släpredskap, bottenlevande arter, som anges i bilaga I till förordning (EG) nr 2027/95 skall anpassas i enlighet med vad som anges i bilagan.
Artikel 2
Denna förordning träder i kraft dagen efter det att den offentliggörs i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1365/97 av den 16 juli 1997 om ändring av förordning (EG) nr 716/96 om undantagsåtgärder till stöd för nötköttsmarknaden i Förenade kungariket
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött (1), senast ändrad genom kommissionens förordning (EG) nr 2222/96 (2), särskilt artikel 23 i denna, och
med beaktande av följande: I kommissionens förordning (EG) nr 716/96 (3), senast ändrad genom förordning (EG) nr 2423/96 (4), föreskrivs undantagsåtgärder till stöd för nötköttsmarknaden i Förenade kungariket, särskilt genom att utbetalning till producenten av 0,9 ecu per kg levande vikt tillåts för djur som slaktas enligt den plan som föreskrivs i förordningen. Med hänsyn till prisutvecklingen i Förenade kungariket bör detta belopp justeras för kor samtidigt som en högsta tillåten vikt föreskrivs för djur som slaktas enligt planen. Denna högsta tillåtna vikt bör fastställas med hänsyn till den genomsnittliga vikten för kor. Följaktligen bör även gemenskapens bidrag, uttryckt i ecu per djur, justeras.
Förvaltningskommittén för nötkött har inte yttrat sig inom den tid som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Det pris som den behöriga myndigheten i Förenade kungariket skall betala till producenterna eller deras ombud enligt artikel 1.1 skall vara:
- 0,8 ecu per kg levande vikt när det gäller kor, och
- 0,9 ecu per kg levande vikt när det gäller alla andra djur.
Ingen betalning utgår för djur vars levande vikt överskrider 560 kg, i förekommande fall beräknad genom tillämpning av koefficienterna i punkt 2.
2. Där det är nödvändigt att väga berörda djur efter slakt för att beräkna vad den levande vikten skulle ha varit, skall man multiplicera slaktvikten efter avblodning, avhudning, urtagning samt avlägsnande av klövar och hud med en koefficient på
- 2, när det gäller kor, och
- 1,70 när det gäller alla andra djur.
3. Gemenskapen skall medfinansiera den utgift som Förenade kungariket haft för de inköp som avses i artikel 1.1 till ett pris av 291 ecu per inköpt ko och 328 ecu per inköpt djur för alla andra djur som har destruerats i enlighet med bestämmelserna i artikel 1.
Ett förskott på 80 % av det medfinansierade beloppet skall i enlighet med artikel 1.2 betalas ut efter det att de uppköpta djuren slaktats.
4. Om det köp som avses i artikel 1.1 avser ett kastrerat nötkreatur av hankön, skall utbetalningen av hela det pris som avses i punkt 1 endast göras om det sålda djuret inte omfattas av den ansökan om säsongsutjämningsbidrag som avses i artikel 4c i förordning (EEG) nr 805/68.
Producenten eller hans ombud förbinder sig att försäkra att detta bidrag inte har sökts för djuret i fråga.
Om denna förbindelse inte görs skall det pris som skall betalas enligt punkt 1 för djuret i fråga nedsättas till ett belopp motsvarande det belopp som tillämpas för säsongsutjämningsbidraget. Om en premieansökan lämnas in för djuret i fråga, skall den berörda producenten tvingas betala tillbaka ett belopp motsvarande det belopp som tillämpas för säsongsutjämningsbidraget av det pris han erhållit för djuret i fråga. I båda dessa fall skall den andel medfinansiering från gemenskapen som avses i punkt 3 nedsättas med ett belopp motsvarande det belopp som skall tillämpas för säsongsutjämningsbidraget.
5. Den omräkningskurs som skall tillämpas är den jordbruksomräkningskurs som gäller den första dagen i den månad då djuret i fråga köps."
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
RÅDETS FÖRORDNING (EG) nr 2046/97 av den 13 oktober 1997 om samarbete mellan nordliga och sydliga länder i kampen mot narkotika och narkotikamissbruk
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 130 w i detta,
med beaktande av kommissionens förslag (1),
i enlighet med förfarandet i artikel 189 c i fördraget (2), och med beaktande av följande:
Verkningarna av en ekonomi som baseras på framställning av narkotika - eller som gör stora förtjänster på detta - på strukturen hos ett samhälle under utveckling, äventyrar en harmonisk integration av landet i världsekonomin.
Snedvridningen av de sociala strukturerna i utvecklingsländerna på grund av narkotikamissbruk och den industri som är knuten till detta, skadar den hållbara sociala utvecklingen och hindrar uppnåendet av målen för gemenskapens politik inom området för utvecklingssamarbete enligt artikel 130 u i fördraget.
Inom ramen för kampen mot utbudet av narkotika är det synnerligen väsentligt att fattigdomen i söder minskas radikalt och att befolkningen erbjuds ett lagligt alternativ till den olagliga odlingen.
Det är lämpligt att ge de utvecklingsländer som begär det ett institutionellt stöd för att de skall kunna bekämpa narkotikan mer effektivt.
I sitt meddelande av den 23 juni 1994 till Europaparlamentet och rådet, lade kommissionen fram sina riktlinjer för en åtgärdsplan för Europeiska unionen som rör kampen mot narkotika (1995-1999), särskilt på internationell nivå.
Europaparlamentet avgav ett yttrande om dessa riktlinjer den 15 juni 1995.
Den fjärde AVS-EG-konventionen och de avtal om samarbete, association eller partnerskap som har ingåtts mellan gemenskapen och utvecklingsländerna innehåller klausuler om samarbete i kampen mot narkotikamissbruk och illegal handel med narkotika, kontroll av handeln med prekursorer, kemiska produkter och psykotropa ämnen samt utbyte av relevant information, inklusive åtgärder när det gäller penningtvätt. Det finns också ett samband mellan kampen mot narkotika och narkotikamissbruk och målen för samarbetet mellan gemenskapen och utvecklingsländerna.
Den allmänna anslutningen till konventionen ersättande äldre konventioner rörande narkotika från 1961, till samma konvention ändrad enligt protokollet från 1972, till konventionen från 1971 om psykotropa ämnen och till konventionen 1988 mot olaglig hantering av narkotika och psykotropa ämnen, liksom en systematisk tillämpning på nationell och internationell nivå av bestämmelserna i dessa fördrag, utgör hörnstenen i en internationell strategi för att bekämpa missbruk och illegal handel med narkotika.
Europeiska gemenskapen är part i konventionen från 1988, särskilt i kraft av dess artikel 12, och har antagit gemenskapslagstiftning som syftar till kontroll över handeln med prekursorer, efter rekommendationer från den aktionsgrupp för kemiska produkter (GAPC) som skapades av G7 och ordföranden i EG-kommissionen 1989; en grupp som skulle kunna bli effektivare globalt sett om lämplig lagstiftning och lämpliga förfaranden antogs i andra delar av världen.
En effektiv kamp mot narkotika måste också omfatta åtgärder mot penningtvätt som härrör från narkotikahandel, såsom antagandet av en lämplig rättslig ram och lämpliga mekanismer i berörda länder.
De mänskliga rättigheterna måste respekteras när åtgärder genomförs i enlighet med denna förordning.
Europeiska gemenskapens medlemsstater har skrivit under den politiska deklarationen och det globala åtgärdsprogram som antogs av Förenta nationernas generalförsamling vid dess 17:e extramöte.
Ett finansiellt referensbelopp, i betydelsen enligt punkt 2 i förklaringen från Europaparlamentet, rådet och kommissionen av den 6 mars 1995 (3) har införts i den här förordningen för perioden 1998-2000 utan att detta påverkar den budgetansvariga myndighetens befogenheter enligt fördraget.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Inom ramen för sin politik för utvecklingssamarbete och med beaktande av de skadliga verkningarna på utvecklingsinsatserna som framställning, saluförande och konsumtion av narkotika har, skall gemenskapen genomföra samverkansåtgärder inom området narkotika och narkotikamissbruk i utvecklingsländerna, varvid företräde skall ges åt dem som har visat politisk vilja på högsta nivå att lösa sina problem med narkotika. Förekomsten av en sådan vilja kan manifesteras bl.a. genom ratificering av konventionen från 1961, ändrad genom protokollet från 1972, konventionen från 1971 och konventionen från 1988. Utvecklingsländernas engagemang skall ta sig uttryck bl.a. i genomförandet av inhemsk lagstiftning mot penningtvätt som härrör från illegal handel med narkotika.
Artikel 2
Det bistånd som ges i enlighet med denna artikel skall komplettera och förstärka bistånd som lämnas enligt andra instrument för utvecklingssamarbete.
Artikel 3
Gemenskapen skall prioritera begäran från ett samarbetsland om att stödja utarbetandet av en nationell övergripande plan för narkotikakontroll, i nära samarbete med Förenta nationernas program för narkotikakontroll (UNDCP). Dessa planer skall fastställa mål, strategier och prioriteringar i kampen mot narkotika och därtill knutna krav på resurser (inklusive finansiella krav), för att kunna skapa ett integrerat, tvärvetenskapligt angreppssätt som spänner över flera områden och kan ge bästa möjliga effektivitet i nationella program för narkotikakontroll och internationellt bistånd.
Att förebygga narkotikamissbruk och att minska efterfrågan bör ingå som åtgärder i en konsekvent politik som innefattar utbildning och objektiv information om följderna av narkotikamissbruk, främst riktad mot de unga.
Samarbete inom gemenskapen skall ha formen av en dialog som återspeglar de genuina kulturskillnader som påverkar synen på problem som är knutna till narkotikan; detta är avgörande för att se till att strategierna för narkotikakontroll blir socialt och politiskt möjliga att genomföra.
Artikel 4
Gemenskapen skall helst arbeta inom den strategiska ram som har lagts fast i de nationella planerna, och skall även stödja särskilda aktioner med mätbar inverkan (dvs. effektiva och påtagliga resultat inom en i förväg fastställd tidsperiod) på följande områden:
- Utveckling av den institutionella kapaciteten, särskilt för att:
- utvecklingsländerna skall kunna genomföra "National Drug Control Master Plans", och
- avtalen mellan gemenskapen och vissa utvecklingsländer skall kunna genomföras, särskilt när det gäller att bekämpa att kemiska prekursorer kommer på avvägar och kampen mot penningtvätt.
- Minska efterfrågan främst genom analys av fenomenet på lokal nivå, inrättandet av kontrollmekanismer riktade mot handeln med och konsumtionen av narkotika liksom av psykotropa ämnen, behandling och återanpassning av narkotikamissbrukare, och även att minska riskerna. Dessa aktioner bör integreras i den politik som förs på hälso- och utbildningsområdet, utveckling och kamp mot fattigdom och ekonomisk och social utslagning.
- Främja pilotprojekt för alternativ utveckling; genom denna process kan på lång sikt odling av illegal narkotika såväl bekämpas som elimineras genom lämpliga åtgärder för landsbygdsutveckling inom ramen för en hållbar ekonomisk tillväxt nationellt. Dessa projekt skall innefatta ekonomiska och sociala åtgärder som tar hänsyn till de faktorer som bidrar till den illegala framställningen och samtidigt åtgärder som kan underlätta ett bättre utnyttjande av handelsförmånerna. I detta sammanhang skall systematiska undersökningar genomföras om det är möjligt att ytterligare utnyttja andra finansiella gemenskapsinstrument (till exempel ALA) och Europeiska utvecklingsfonden för projekt för alternativ utveckling.
- finansiering av studier, seminarier och forum för erfarenhetsutbyte inom ovannämnda områden.
Särskild uppmärksamhet skall ägnas åt att få lokalbefolkningen och målgrupper att delta när aktionerna beslutas, planeras och genomförs.
Gemenskapen ger endast stöd till projekt i vilka respekten för de mänskliga rättigheterna garanteras.
Artikel 5
Samarbetsparter som är berättigade till finansiellt stöd enligt denna förordning skall vara regionala och internationella organisationer, särskilt UNDCP, lokala och i medlemsstaterna förankrade icke-statliga organisationer, nationella, regionala och lokala styrande organ och myndigheter, organisationer förankrade i lokalsamhället, institut samt offentliga och privata aktörer.
Artikel 6
1. De instrument som skall användas för åtgärderna enligt artiklarna 3 och 4 skall innefatta studier, tekniskt bistånd, utbildning eller andra tjänster, leveranser och anläggningar, liksom även revision samt utvärderings- och övervakningsuppdrag.
2. Gemenskapens finansiering kan, beroende på behoven för varje åtgärd, täcka såväl investeringskostnader, med undantag av fastighetsköp, som driftskostnader i utländsk eller inhemsk valuta. Med undantag av utbildningsprogrammen skall dock driftskostnaderna normalt täckas endast under inledningsfasen, för att sedan gradvis minska.
3. Ekonomiska bidrag från de parter som anges i artikel 5 skall sökas för alla samarbetsåtgärder. Bidrag skall begäras inom ramen för de berörda parternas möjligheter och med hänsyn till varje åtgärds art.
4. Ekonomiska bidrag från lokala samarbetsparter, i synnerhet till driftskostnaderna, skall sökas som en prioriterad åtgärd när det gäller projekt med syfte att sätta igång långsiktig verksamhet, för att på så sätt säkerställa att sådana projekt lever vidare då gemenskapsbidragen upphör.
5. Möjligheter till samfinansiering med andra bidragsgivare, i synnerhet medlemsstaterna, kan undersökas.
6. Kommissionen skall säkerställa att gemenskapskaraktären på det bistånd som ges i enlighet med denna förordning framhävs.
7. För att kunna uppnå fördragets mål om konsekvens och komplementaritet och i syfte att optimera effekten av alla dessa åtgärder kan kommissionen vidta alla de nödvändiga samordningsåtgärderna, i synnerhet
a) inrätta ett system för systematiskt utbyte och analys av information om finansierade åtgärder samt de åtgärder som gemenskapen och medlemsstaterna har för avsikt att finansiera,
b) samordning på plats av genomförandet av åtgärderna med hjälp av regelbundna möten och utbyte av information mellan kommissionens och medlemsstaternas företrädare i mottagarlandet.
8. I syfte att få största möjliga verkan så väl globalt som nationellt, skall kommissionen tillsammans med medlemsstaterna ta alla initiativ som krävs för att säkerställa god samordning och nära samarbete med mottagarländerna och bidragsgivarna samt andra internationella organ som berörs, i synnerhet de som ingår i Förenta nationernas organisation och då särskilt UNDCP.
Artikel 7
Det ekonomiska stöd som ges enligt denna förordning skall vara i form av gåvobistånd.
Artikel 8
Det finansiella referensbeloppet för att genomföra detta program är 30 miljoner ecu för perioden 1998-2000.
Årliga anslag skall beviljas av budgetmyndigheten inom budgetramarna.
Artikel 9
1. Kommissionen skall ansvara för bedömning, godkännande och förvaltning av de åtgärder som omfattas av denna förordning enligt gällande budgetförfaranden och andra gällande förfaranden, särskilt de som föreskrivs i budgetförordningen för Europeiska gemenskapernas allmänna budget.
2. Vid bedömningen av projekt och program skall följande faktorer beaktas:
- Effekten av och möjligheten att genomföra åtgärderna.
- Kulturella och sociala aspekter samt genus- och miljöaspekter.
- Vilken institutionell utveckling som är nödvändig för att projektmålen skall kunna uppnås.
- Erfarenheter av åtgärder av samma typ.
3. Beslut om finansiering som överskrider 2 miljoner ecu för enskilda åtgärder enligt denna förordning samt alla förändringar som ger en ökning på mer än 20 % av den summa som ursprungligen godkänts för en sådan åtgärd, skall fattas enligt det förfarande som föreskrivs i artikel 10.
Kommissionen skall kortfattat informera den kommitté som avses i artikel 10 om de finansieringsbeslut som den ämnar fatta avseende projekt och program vars kostnad understiger 2 miljoner ecu. Sådan information skall lämnas senast en vecka innan beslutet fattas.
4. Kommissionen bemyndigas att, utan dessförinnan höra den kommitté som avses i artikel 10, godkänna de ytterligare åtaganden som kan behövas för att täcka sådana överskridanden som kan förutses eller som har konstaterats i samband med dessa åtgärder om överskridandet uppgår till högst 20 % av det ursprungliga åtagande som fastställdes genom finansieringsbeslutet.
5. I alla överenskommelser eller kontrakt om finansiering som ingås enligt denna förordning, skall föreskrivas särskilt att kommissionen och revisionsrätten kan utföra kontroller på plats i enlighet med de sedvanliga villkor som kommissionen fastställer inom ramen för gällande bestämmelser, särskilt bestämmelserna i budgetförordningen för Europeiska gemenskapernas allmänna budget.
6. Om åtgärderna är föremål för finansieringsöverenskommelser mellan gemenskapen och mottagarlandet, skall i dessa föreskrivas att betalning av skatter, tullar och andra avgifter inte skall erläggas av gemenskapen.
7. Deltagande i anbudsförfaranden och i avtal skall vara öppet på lika villkor för alla fysiska och juridiska personer i medlemsstaterna och mottagarlandet. Det kan utsträckas till andra utvecklingsländer.
8. Leveranser skall härröra från medlemsstaterna, mottagarlandet eller andra utvecklingsländer. I vederbörligen styrkta undantagsfall kan leveranser härröra från andra länder.
9. Särskild uppmärksamhet skall ägnas
- strävan efter kostnadseffektivitet och en varaktig inverkan i samband med att projekten utformas, och
- klart definierade och övervakade mål samt genomförandeindikatorer för samtliga projekt.
Artikel 10
1. Kommissionen skall biträdas av den behöriga geografiska kommittén för utvecklingssamarbete.
2. Kommissionens företrädare skall förelägga kommittén ett utkast till de åtgärder som skall vidtas. Kommittén skall yttra sig över utkastet inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Medlemsstaternas röster skall vägas enligt bestämmelserna i samma artikel. Ordföranden får inte rösta.
Kommissionen skall själv anta de planerade åtgärderna om de är förenliga med kommitténs yttrande.
Om de planerade åtgärderna inte är förenliga med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
3. En gång om året skall en diskussion hållas på grundval av en framställning av kommissionens företrädare om de allmänna riktlinjerna för de åtgärder som skall vidtas under det kommande året inom de kommittéer som avses i punkt 1.
Artikel 11
1. Efter varje budgetår skall kommissionen överlämna en årsrapport till Europaparlamentet och rådet med en sammanfattning av de åtgärder som finansierats under budgetåret samt en utvärdering av hur denna förordning genomförts under denna period.
Sammanfattningen skall i synnerhet innehålla upplysningar om dem med vilka avtal eller kontrakt har slutits.
2. Kommissionen skall regelbundet utvärdera de åtgärder som gemenskapen finansierar för att fastställa om de mål som ställdes upp för dessa åtgärder har uppnåtts och för att ange riktlinjer för att förbättra framtida åtgärders effektivitet. Kommissionen skall överlämna en sammanfattning av de utvärderingar som gjorts till den kommitté som avses i artikel 10, vilka denna kommitté i förekommande skall kunna granska. Utvärderingsrapporterna skall finnas tillgängliga för de medlemsstater som önskar ta del av dem.
3. Kommissionen skall, senast en månad efter det att den fattat sitt beslut, informera medlemsstaterna om godkända åtgärder och projekt med uppgift om kostnad, art, mottagarland och parter.
Artikel 12
1. Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS BESLUT av den 25 februari 1998 om ett frågeformulär för medlemsstaternas rapporter om genomförande av rådets direktiv 94/67/EG om förbränning av farligt avfall (genomförande av rådets direktiv 91/692/EEG) (Text av betydelse för EES) (98/184/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/692/EEG av den 23 december 1991 om att standardisera och rationalisera rapporterna om genomförandet av vissa direktiv om miljön (1), särskilt artiklarna 5 och 6 i detta,
med beaktande av rådets direktiv 94/67/EG om förbränning av farligt avfall (2), och
med beaktande av följande: I artikel 17 i direktiv 94/67/EG fastställs att medlemsstaterna skall rapportera om genomförandet av detta direktiv i enlighet med artikel 5 i direktiv 91/692/EEG.
Rapporten skall utarbetas på grundval av frågeformulär eller mallar som kommissionen fastställer i enlighet med förfarandet i artikel 6 i direktiv 91/692/EG.
Den första rapporten kommer att omfatta åren från och med 1998 till och med 2000.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som upprättats i enlighet med artikel 6 i ovan nämnda direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Det frågeformulär som bifogas detta beslut, och som skall användas i samband med rådets direktiv 94/67/EG om förbränning av farligt avfall, antas härmed.
Artikel 2
Medlemsstaterna skall använda frågeformuläret som underlag när de utarbetar den rapport som de skall lämna till kommissionen i enlighet med artikel 5 i direktiv 91/692/EEG och artikel 17 i direktiv 94/67/EG.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 29 juli 1998 om ändring av rådets beslut 96/411/EG om förbättring av gemenskapens jordbruksstatistik [delgivet med nr K(1998) 2135] (Text av betydelse för EES) (98/514/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets beslut 96/411/EG av den 25 juni 1996 om förbättring av gemenskapens jordbruksstatistik (1), ändrat genom beslut 98/3/EG (2), särskilt artikel 8 i detta, och av följande skäl:
Att slå vakt om kvaliteten på landsbygdsmiljön är ett av målen för politiken för landsbygdens utveckling.
För detta ändamål bör beslut 94/411/EG ändras genom att dess bilaga II ersätts.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för jordbruksstatistik.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga II till beslut 96/411/EG skall ersättas med bilagan till detta beslut.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
RÅDETS BESLUT av den 20 juli 1998 om ingående av ett avtal om ömsesidigt erkännande mellan Europeiska gemenskapen och Kanada (98/566/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113, tillsammans med artikel 228.2 första meningen och 228.3 första stycket, samt artikel 228.4 i detta,
med beaktande av kommissionens förslag, och
av följande skål: Avtalet om ömsesidigt erkännande mellan Europeiska gemenskapen och Kanada, vilket undertecknades i London den 14 maj 1998, har framförhandlats och bör godkännas.
Vissa genomförandeuppgifter har anförtrotts den gemensamma kommitté som inrättas genom avtalet, särskilt befogenheten att ändra vissa aspekter av de sektoriella bilagorna till detta.
För att säkerställa att avtalet fungerar korrekt bör lämpliga interna förfaranden fastställas och det är nödvändigt att bemyndiga kommissionen att göra vissa ändringar av teknisk natur i avtalet och att fatta vissa beslut för dess genomförande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Avtalet om ömsesidigt erkännande mellan Europeiska gemenskapen och Kanada, inbegripet dess bilagor, godkänns härmed på Europeiska gemenskapens vägnar.
Texten till avtalet och bilagorna till det bifogas detta beslut.
Artikel 2
Rådets ordförande skall på gemenskapens vägnar överlämna den skrivelse som avses i artikel XIX i avtalet.
Artikel 3
1. Gemenskapen skall i den gemensamma kommitté som föreskrivs i artikel XI i avtalet och i de gemensamma sektoriella grupper som föreskrivs i artikel XII i avtalet och som inrättas genom de sektoriella bilagorna företrädas av kommissionen, som skall biträdas av den särskilda kommitté som utsetts av rådet. Kommissionen skall efter samråd med denna särskilda kommitté verkställa de utseenden, det informationsutbyte och de framställningar om kontroller som avses i artiklarna IX, X, XI.3 c och e, XII b och XIII i avtalet och i motsvarande bestämmelser i de sektoriella bilagorna.
2. Gemenskapens ståndpunkt vad gäller beslut som skall fattas av den gemensamma kommittén eller i förekommande fall av de gemensamma sektoriella grupperna skall, såvitt gäller ändringar i de sektoriella bilagorna (artikel XI.3 a och XI.4 i avtalet) och kontroll enligt artiklarna VIII och XI.4 c i avtalet av att gällande krav är uppfyllda, fastställas av kommissionen efter samråd med den särskilda kommitté som avses i punkt 1 i den här artikeln.
3. I samtliga övriga fall skall gemenskapens ståndpunkt i den gemensamma kommittén eller i de gemensamma sektoriella grupperna fastställas av rådet som skall fatta sina beslut med kvalificerad majoritet på förslag av kommissionen. Samma förfarande skall gälla för beslut som fattas av gemenskapen inom ramen för artiklarna XV.3 och XIX.4 i avtalet.
RÅDETS DIREKTIV 98/29/EG av den 7 maj 1998 om harmonisering av huvudbestämmelserna för kreditförsäkringar för medellånga och långa exportaffärer
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113 i detta,
med beaktande av kommissionens förslag, och
med beaktande av följande: (1) Kreditförsäkringar för medellånga och långa exportaffärer spelar en viktig roll i internationell handel och utgör ett viktigt handelspolitiskt instrument.
(2) Kreditförsäkringar för medellånga och långa exportaffärer spelar en viktig roll för handeln med utvecklingsländer och främjar dessa länders integrering med världsekonomin, vilket är ett mål för gemenskapens utvecklingspolitik.
(3) Skillnaderna mellan medlemsstaternas nu existerande statsstödda system för kreditförsäkringar för medellånga och långa exportaffärer med avseende på de huvudsakliga beståndsdelarna i försäkringsskyddet, premiebestämmelserna och täckningspolitiken kan leda till att konkurrensen mellan företag inom gemenskapen snedvrids.
(4) De åtgärder som föreskrivs i detta direktiv bör inte gå utöver vad som är nödvändigt för att uppnå det mål, som består i att åstadkomma den harmonisering som är nödvändig för att säkerställa att exportpolitiken grundas på enhetliga principer och att konkurrensen mellan företagen inom gemenskapen inte snedvrids.
(5) För att minska befintlig snedvridning av konkurrensen är det önskvärt att de olika statsstödda systemen för exportkreditförsäkringar harmoniseras enligt artikel 112 i fördraget, på grundval av enhetliga principer och på ett sådant sätt att de bildar en integrerad del av den gemensamma handelspolitiken.
(6) Regeringars (eller särskilda av regeringar kontrollerade institutioners) tillhandahållande av exportkreditgarantisystem eller exportkreditförsäkringssystem till premier som är otillräckliga för att täcka systemens långsiktiga kostnader och förluster betraktas som förbjudna exportsubventioner i det avtal om subventioner och utjämningsåtgärder som ingicks inom ramen för de multilaterala handelsförhandlingarna i Uruguayrundan (1986-1994) (1) (se artikel 3.1 a och bilaga I j till avtalet).
(7) Den premie som kreditförsäkraren tar ut bör motsvara den risk som försäkras.
(8) En harmonisering skulle gynna samarbete mellan de kreditförsäkrare som agerar på en stats vägnar eller med statligt stöd, och öka samarbetet mellan företag inom gemenskapen enligt artikel 130 i fördraget.
(9) Både harmonisering och samarbete är huvudsakliga och avgörande faktorer för gemenskapsexportens konkurrenskraft på marknader utanför gemenskapen.
(10) I kommissionens vitbok om den inre marknadens fullbordande som antogs av Europeiska rådet i juni 1985 betonas vikten av ett samarbetsvänligt klimat hos gemenskapens företag.
(11) Genom sitt beslut (2) av den 27 september 1960 inrättade rådet en arbetsgrupp för samordning av politiken för kreditförsäkringar, kreditgarantier och finansiella krediter.
(12) Den 15 maj 1991 gav den nämnda arbetsgruppen mandat till experter från var och en av de dåvarande medlemsstaterna vilka, under namnet Expertgruppen för den inre marknaden 1992, den 27 mars 1992, den 11 juni 1993 och den 9 februari 1994 lade fram rapporter, som innehöll ett antal förslag.
(13) Genom beslut 93/112/EEG (3) genomförde rådet OECD-överenskommelsen om riktlinjer för exportkrediter med offentligt stöd i gemenskapsrätten.
(14) Rådets direktiv 70/509/EEG av den 27 oktober 1970 om antagande av gemensamma kreditförsäkringsvillkor för medellånga och långa exportaffärer med offentliga köpare (4), och rådets direktiv 70/510/EEG av den 27 oktober 1970 om antagande av gemensamma kreditförsäkringsvillkor för medellånga och långa exportaffärer med privata köpare (5), bör ersättas med det här direktivet.
(15) Denna begynnande harmonisering av exportkreditförsäkringarna bör ses som ett steg i riktning mot samstämmighet mellan medlemsstaternas olika system.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Tillämpningsområde
Detta direktiv är tillämpligt på försäkringsskydd för affärer avseende export av varor och/eller tjänster med ursprung i en medlemsstat, under förutsättning att detta stöd ges, direkt eller indirekt, för en eller flera medlemsstaters räkning eller med stöd av en eller flera medlemsstater och omfattar en total riskperiod på minst två år, dvs. återbetalningsperioden inklusive tillverkningsperioden.
Detta direktiv gäller varken försäkringsskydd för anbud, förskottsbetalning eller fullgörandegarantier och inte heller försäkring för säkerhet för "retention money", så kallad retention payment bond. Det gäller inte heller försäkringsskydd för risker avseende byggutrustning och byggmaterial när dessa används lokalt för att fullgöra ett affärsavtal.
Artikel 2
Medlemsstaternas skyldigheter
Medlemsstaterna skall se till att alla institut, som direkt eller indirekt erbjuder försäkringsskydd i form av exportkreditförsäkringar, garantier eller refinansiering för medlemsstatens räkning eller med stöd av den medlemsstat som företräder själva regeringen eller som kontrolleras av och/eller handlar enligt bemyndigande av den regering som erbjuder försäkringsskydd, nedan kallade försäkringsgivare, erbjuder försäkringsskydd för affärer avseende export av varor och/eller tjänster i enlighet med bestämmelserna i bilagan, när exportaffärerna görs med länder utanför gemenskapen och finansieras med hjälp av köparkrediter eller leverantörskrediter eller betalas kontant.
Artikel 3
Genomförandebeslut
De beslut som avses i punkt 46 i bilagan skall fattas av kommissionen i enlighet med det förfarande som avses i artikel 4.
Artikel 4
Kommitté
Kommissionen skall biträdas av en kommitté som skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Den skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Medlemsstaternas röster skall vägas enligt bestämmelserna i samma artikel. Ordföranden får inte rösta.
Kommissionen skall besluta med omedelbar verkan. Om beslutet inte är förenligt med kommitténs yttrande skall kommissionen emellertid genast underrätta rådet. I sådana fall:
- Skall kommissionen uppskjuta verkställandet av de beslutade åtgärderna under en tid som inte överstiger en månad från den dag då rådet underrättats.
- Får rådet fatta ett annat beslut med kvalificerad majoritet inom den tid som anges i första strecksatsen.
Artikel 5
Rapport och översyn
Kommissionen skall senast den 31 december 2001 förelägga rådet en rapport om de erfarenheter som gjorts och den samstämmighet som uppnåtts vid tillämpning av bestämmelserna i detta direktiv.
Artikel 6
Förhållande till andra förfaranden
De förfaranden som föreskrivs i detta direktiv kompletterar dem som inrättas genom beslut 73/391/EEG (6).
Artikel 7
Upphävande
Direktiv 70/509/EEG och direktiv 70/510/EEG upphävs.
Artikel 8
Överföring
Artikel 9
Ikraftträdande
RÅDETS DIREKTIV 98/49/EG av den 29 juni 1998 om skydd av kompletterande pensionsrättigheter för anställda och egenföretagare som flyttar inom gemenskapen
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 51 och 235 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
av följande skäl: (1) En av de grundläggande friheterna i gemenskapen är fri rörlighet för personer. I fördraget föreskrivs att rådet enhälligt skall besluta om sådana åtgärder inom den sociala trygghetens område som är nödvändiga för att genomföra fri rörlighet för arbetstagare.
(2) Arbetstagarnas sociala skydd säkerställs genom lagstadgade system för social trygghet som supplerar kompletterande system för social trygghet.
(3) Den lagstiftning som rådet redan har antagit för att skydda rättigheterna på den sociala trygghetens område för de arbetstagare och deras familjemedlemmar som flyttar inom gemenskapen, det vill säga rådets förordningar (EEG) nr 1408/71 av den 14 juli 1971 om tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen (4) och (EEG) nr 574/72 av den 21 mars 1972 om tillämpning av förordning (EEG) nr 1408/71 om tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen (5), avser endast lagstadgade pensionssystem; det samordningssystem som föreskrivs i dessa förordningar omfattar inte kompletterande pensionssystem med undantag för system som täcks av begreppet "lagstiftning" enligt definitionen i artikel 1 j första stycket i förordning (EEG) nr 1408/71 eller med avseende på vilka en medlemsstat avger en förklaring enligt den artikeln.
(4) Rådet äger stor frihet när det gäller valet av vilka åtgärder som är bäst lämpade för att uppnå målet i artikel 51 i fördraget; det samordningssystem som avses i förordningarna (EEG) nr 1408/71 och (EEG) nr 574/72, och särskilt reglerna för sammanläggning, passar inte för kompletterande pensionssystem, med undantag för system som täcks av begreppet "lagstiftning" enligt definitionen i artikel 1 j första stycket i förordning (EEG) nr 1408/71 eller med avseende på vilka en medlemsstat avger en förklaring enligt den artikeln, och bör därför bli föremål för särskilda åtgärder, av vilka detta direktiv är den första, så att hänsyn kan tas till deras särskilda karaktär och kännetecken och till olikheterna mellan sådana system inom och mellan medlemsstaterna.
(5) Ingen pension eller förmån bör omfattas både av bestämmelserna i detta direktiv och av förordningarna (EEG) nr 1408/71 och (EEG) nr 574/72 och därför kan ett kompletterande pensionssystem, som ligger inom dessa förordningars räckvidd därför att en medlemsstat har avgett en förklaring av denna innebörd enligt artikel 1 j i förordning (EEG) nr 1408/71, inte omfattas av bestämmelserna i detta direktiv.
(6) I sin rekommendation 92/442/EEG av den 27 juli 1992 om samstämmighet mellan mål och politik på det sociala skyddets område (6) rekommenderar rådet medlemsstaterna att "vid behov främja ändringar av villkoren för förvärv av rätt till pension, särskilt kompletterande pensionsrättigheter, för att avskaffa hindren för anställdas rörlighet".
(7) Ett bidrag till att nå detta mål kan vara att arbetstagare, som flyttar eller vilkas arbetsplats flyttar från en medlemsstat till en annan, i fråga om skyddet för deras kompletterande pensionsrättigheter garanteras en behandling som är likvärdig med den som ges arbetstagare som stannar kvar eller vilkas arbetsplats stannar kvar inom samma medlemsstat.
(8) Den fria rörligheten för personer, som är en av de grundläggande rättigheterna i fördraget, är inte begränsad till anställda utan omfattar också egenföretagare.
(9) Fördraget innehåller inga andra befogenheter än de som finns i artikel 235 för att vidta lämpliga åtgärder på området social trygghet för egenföretagare.
(10) För att rätten till fri rörlighet skall kunna utövas på ett effektivt sätt bör arbetstagare och andra berättigade personer ha vissa garantier för lika behandling i fråga om bevarandet av sina intjänade pensionsrättigheter enligt kompletterande pensionssystem.
(11) Medlemsstaterna bör vidta de åtgärder som behövs för att se till att förmåner enligt kompletterande pensionssystem betalas ut till försäkringstagare och före detta försäkringstagare samt till andra personer som är berättigade enligt sådana system i alla medlemsstater, eftersom alla restriktioner för betalningar och kapitalrörelser är förbjudna enligt artikel 73 b i fördraget.
(12) För att underlätta utövandet av rätten till fri rörlighet bör, när så behövs, nationella bestämmelser i enlighet med avdelning II i förordning (EEG) nr 1408/71 anpassas så att det blir möjligt att fortsätta att betala in avgifter till ett kompletterande pensionssystem i en medlemsstat från eller för arbetstagare som är utsända till en annan medlemsstat.
(13) I detta avseende krävs enligt fördraget inte bara avskaffande av diskriminering av arbetstagare i medlemsstaterna på grund av medborgarskap utan även undanröjande av alla nationella bestämmelser som kan hindra dessa arbetstagares utövande av, eller göra det mindre attraktivt för dem att utöva, de grundläggande friheter som garanteras i fördraget, enligt Europeiska gemenskapernas domstols tolkning i flera på varandra följande domar.
(14) De arbetstagare som utövar sin rätt till fri rörlighet bör på ett adekvat sätt informeras av arbetsgivare, förvaltare eller andra som har ansvar för förvaltningen av de kompletterande pensionssystemen, särskilt vad gäller de val och de alternativ som erbjuds dem.
(15) Detta direktiv påverkar inte medlemsstaternas lagar ifråga om kollektiva åtgärder för att försvara yrkesintressen.
(16) På grund av mångfalden av kompletterande system för social trygghet bör gemenskapen endast ställa upp allmänna mål och därför är ett direktiv det lämpliga rättsliga instrumentet.
(17) I enlighet med subsidiaritets- och proportionalitetsprinciperna i artikel 3 b i fördraget kan målen för detta direktiv inte i tillräcklig utsträckning uppnås av medlemsstaterna utan de kan uppnås bättre på gemenskapsnivå. Detta direktiv går inte utöver vad som är nödvändigt för att uppnå dessa mål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
SYFTE OCH RÄCKVIDD
Artikel 1
Syftet med detta direktiv är att skydda rättigheterna för de försäkringstagare som omfattas av kompletterande pensionssystem och som flyttar från en medlemsstat till en annan och att därigenom bidra till att undanröja hinder för den fria rörligheten för anställda och egenföretagare inom gemenskapen. Detta skydd avser pensionsrättigheter enligt både frivilliga och obligatoriska kompletterande pensionssystem, med undantag av de system som omfattas av förordning (EEG) nr 1408/71.
Artikel 2
Detta direktiv skall tillämpas på försäkringstagare som omfattas av kompletterande pensionssystem och andra personer som är berättigade enligt sådana system och som har förvärvat eller håller på att förvärva rättigheter i en eller flera medlemsstater.
KAPITEL II
DEFINITIONER
Artikel 3
I detta direktiv används följande beteckningar med de betydelser som här anges:
a) kompletterande pension: ålderspension och, om det föreskrivs i bestämmelserna för ett i enlighet med nationell lagstiftning och praxis inrättat kompletterande pensionssystem, invaliditets- och efterlevandeförmåner som är avsedda att komplettera eller ersätta de förmåner som de lagstadgade systemen för social trygghet föreskriver för samma försäkringsfall,
b) kompletterande pensionssystem: alla i enlighet med nationell lagstiftning och praxis inrättade tjänstepensionssystem, såsom gruppförsäkringsavtal eller system med löpande inbetalning ("pay as you go") om vilka en eller flera branscher eller sektorer kommit överens, premiereservsystem eller utfästelser om pension som garanteras av bokförda reserver, eller alla kollektiva eller andra jämförbara system vilka är avsedda som en kompletterande pension för anställda eller egenföretagare,
c) pensionsrättigheter: alla förmåner som försäkringstagare och andra berättigade personer har rätt till enligt bestämmelserna i ett kompletterande pensionssystem och, i förekommande fall, enligt nationell lagstiftning,
d) intjänade pensionsrättigheter: alla rättigheter till förmåner som erhålls efter uppfyllande av de krav som ställs enligt reglerna för ett kompletterande pensionssystem och, i förekommande fall, enligt nationell lagstiftning,
e) utsänd arbetstagare: en person som är utsänd till en annan medlemsstat för att arbeta och som enligt villkoren i avdelning II i förordning (EEG) nr 1408/71 fortsätter att omfattas av ursprungsmedlemsstatens lagstiftning; utsändning skall tolkas i enlighet härmed,
f) avgift: alla betalningar som gjorts eller anses ha gjorts till ett kompletterande pensionssystem.
KAPITEL III
ÅTGÄRDER FÖR ATT SKYDDA KOMPLETTERANDE PENSIONSRÄTTIGHETER FÖR ARBETSTAGARE SOM FLYTTAR INOM GEMENSKAPEN
Artikel 4
Likabehandling i fråga om bevarande av pensionsrättigheter
Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa bevarande av intjänade pensionsrättigheter för de personer, som är försäkringstagare enligt ett kompletterande pensionssystem och för vilka avgifter inte längre betalas därför att de har flyttat från en medlemsstat till en annan medlemsstat, i samma utsträckning som för de försäkringstagare för vilka avgifter inte längre betalas men som bor kvar i samma medlemsstat. Denna artikel skall också tillämpas på andra personer som är berättigade enligt bestämmelserna för det kompletterande pensionssystemet i fråga.
Artikel 5
Gränsöverskridande betalningar
Medlemsstaterna skall se till att de kompletterande pensionssystemen till försäkringstagare och andra personer som är berättigade enligt dessa system i andra medlemsstater betalar ut alla förmåner som utfaller enligt dessa system, efter avdrag för de skatter och transaktionskostnader som kan vara tillämpliga.
Artikel 6
Avgifter till kompletterande pensionssystem från eller för utsända arbetstagare
1. Medlemsstaterna skall besluta om sådana åtgärder som behövs för att göra det möjligt att fortsätta att betala avgifter från eller för en utsänd arbetstagare som är försäkringstagare i ett kompletterande pensionssystem i en medlemsstat, under den tid som arbetstagaren är utsänd till en annan medlemsstat.
2. Om avgifter fortsatt betalas in till ett kompletterande pensionssystem i en medlemsstat i enlighet med punkt 1, skall den utsända arbetstagaren och, i förekommande fall, dennas arbetsgivare, vara undantagen från alla förpliktelser att betala in avgifter till ett kompletterande pensionssystem i en annan medlemsstat.
Artikel 7
Information till försäkringstagarna
Medlemsstaterna skall vidta åtgärder så att arbetsgivare, förvaltare eller andra, som har ansvar för förvaltningen av de kompletterande pensionssystemen, när försäkringstagarna flyttar till en annan medlemsstat förser dem med adekvat information i fråga om deras pensionsrättigheter och om de valmöjligheter som finns att tillgå för dem enligt systemet. Denna information skall minst motsvara den information som ges de försäkringstagare för vilka avgifter inte längre betalas men som bor kvar i samma medlemsstat.
KAPITEL IV
SLUTBESTÄMMELSER
Artikel 8
Medlemsstaterna kan föreskriva att bestämmelserna i artikel 6 skall tillämpas endast på utsändningar som påbörjas 25 juli 2001.
Artikel 9
Medlemsstaterna skall i sin nationella lagstiftning införa de bestämmelser som behövs för att alla, som anser sig förfördelade på grund av underlåtenhet att tillämpa bestämmelserna i detta direktiv, skall kunna föra talan vid domstol, efter att i förekommande fall ha vänt sig till andra behöriga myndigheter.
Artikel 10
1. Medlemsstaterna skall sätta i kraft de lagar och författningar som är nödvändiga för att följa detta direktiv senast 36 månader efter det att direktivet har trätt i kraft eller skall säkerställa att arbetsgivare och arbetstagare senast den dagen avtalar om de bestämmelser som krävs. Medlemsstaterna är skyldiga att vidta alla de åtgärder som krävs för att de alltid skall kunna garantera de resultat som föreskrivs i detta direktiv. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
De skall underrätta kommissionen om vilka nationella myndigheter som skall kontaktas vad avser tillämpningen av detta direktiv.
2. Medlemsstaterna skall senast 25 januari 2002 till kommissionen överlämna texten till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
3. På grundval av de upplysningar som medlemsstaterna lämnar skall kommissionen inom sex år efter detta direktivs ikraftträdande överlämna en rapport som till Europaparlamentet, rådet och Ekonomiska och sociala kommittén.
Rapporten skall behandla direktivets tillämpning och skall vid behov innehålla förslag till ändringar som kan behöva göras.
Artikel 11
RÅDETS DIREKTIV 98/57/EG av den 20 juli 1998 om bekämpning av Ralstonia solanacearum (Smith) Yabuuchi m.fl.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
av följande skäl: Skadegöraren Ralstonia solanacearum (Smith) Yabuuchi m.fl. var tidigare känd som Pseudomonas solanacearum (Smith) Smith. Ralstonia solanacearum (Smith) Yabuuchi m.fl. kommer förmodligen att bli det allmänt godtagna namnet på skadegöraren. I detta direktiv bör hänsyn tas till denna vetenskapliga utveckling.
Produktionen av potatis och tomater intar en viktig plats inom gemenskapens jordbruk. Potatis- och tomatskörden hotas ständigt av skadegörare.
Om odlingen av potatis och tomater skyddas mot sådana skadegörare skulle produktionskapaciteten upprätthållas och dessutom skulle jordbruksproduktionen öka.
Skyddsåtgärder mot införsel av skadegörare till en medlemsstats territorium skulle endast ha begränsad effekt om inte sådana skadegörare samtidigt och metodiskt bekämpades inom hela gemenskapen och hindrades från att sprida sig.
En av skadegörarna på potatis och tomat är Ralstonia solanacearum (Smith) Yabuuchi m.fl., den sjukdomsalstrande organism som orsakar mörk ringröta hos potatis och bakteriologisk vissnesjuka hos potatis och tomat. Sjukdomar som orsakats av denna sjukdomsalstrande organism har brutit ut i några delar av gemenskapen, och det existerar fortfarande några begränsade smittkällor.
Det föreligger en avsevärd risk för odlingen av potatis och tomater i hela gemenskapen om effektiva åtgärder inte vidtas med avseende på dessa grödor för att lokalisera denna skadegörare och avgöra dess utbredning, för att förhindra dess förekomst och spridning samt, om den påträffas, för att förhindra dess spridning och bekämpa den i syfte att utrota den.
För att säkerställa detta måste vissa åtgärder vidtas inom gemenskapen. Medlemsstaterna måste dessutom kunna vidta ytterligare eller strängare åtgärder, där detta är nödvändigt förutsatt att dessa inte hindrar handeln med potatis eller tomater inom gemenskapen än de som anges i rådets direktiv 77/93/EEG av den 21 december 1976 om skyddsåtgärder mot att skadegörare på växter eller växtprodukter förs in till medlemsstaterna (4). Sådana åtgärder måste anmälas till de andra medlemsstaterna och till kommissionen.
Åtgärderna måste beakta att systematiska officiella undersökningar är nödvändiga för att lokalisera den sjukdomsalstrande organismen. Sådana undersökningar bör omfatta besiktningar och där så är lämpligt stickprovskontroller och test, eftersom sjukdomen under vissa miljömässiga omständigheter kan förbli latent och obemärkt både i potatisens förökningsmaterial och i lagrade potatisknölar. Spridningen av den sjukdomsalstrande organismen inom förökningsmaterialet är inte den viktigaste faktorn, men eftersom den sjukdomsalstrande organismen kan spridas med ytvatten och genom vissa besläktade vilda växter av familjen Solanaceae, utgör bevattning av potatis- och tomatgrödor med angripet vatten en smittorisk för sådana grödor. Den sjukdomsalstrande organismen kan också övervintra i självsådda (övervintrade) potatis- och tomatplantor, och dessa kan utgöra en smittkälla då de för över smittan från en odlingssäsong till nästa. Den sjukdomsalstrande organismen sprids också genom att potatisplantor angrips vid kontakt med smittad potatis och vid kontakt med utrustning för sättning, upptagning och hantering eller med transport- och lagringsbehållare som har angripits av skadegöraren vid tidigare kontakt med smittad potatis.
Spridningen av den sjukdomsalstrande organismen kan minskas eller förhindras genom desinfektion av sådana föremål. Varje angrepp på utsädespotatis innebär en stor risk för att den sjukdomsalstrande organismen sprids. Utsädespotatisens latenta smitta utgör på liknande sätt en stor risk för att den sjukdomsalstrande organismen sprids, och detta kan förhindras genom användning av utsädespotatis som har producerats i ett officiellt godkänt program, där utsädespotatis har testats och konstaterats vara fri från smitta.
Den nuvarande kunskapen om de biologiska och epidemiologiska egenskaperna hos Ralstonia solanacearum (Smith) Yabuuchi m.fl. under europeiska förhållanden är ofullständig, och det förutses att en översyn av de föreslagna åtgärderna kommer att bli nödvändig om ett antal säsonger. Förbättringar av testprocedurerna förväntas också mot bakgrund av ytterligare forskning, särskilt kring testmetodernas sensibilitet och noggrannhet, för att optimala testmetoder skall kunna väljas ut och standardiseras.
För att närmare kunna besluta om dessa allmänna åtgärder, liksom om de strängare eller ytterligare åtgärder som medlemsstaterna vidtar för att förhindra att den sjukdomsalstrande organismen förs in till deras territorium, är det önskvärt att medlemsstaterna samarbetar nära med kommissionen inom Ständiga kommittén för växtskydd (nedan kallad kommittén).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Detta direktiv rör de åtgärder som i medlemsstaterna skall vidtas mot Ralstonia solanacearum (Smith) Yabuuchi m.fl., tidigare känd som Pseudomonas solanacearum (Smith) Smith (nedan kallad skadegöraren) för att, såvitt avser skadegörarens värdväxter, vilka förtecknas i del 1 i bilaga I, (nedan kallade det förtecknade växtmaterialet),
a) lokalisera skadegöraren och kartlägga dess utbredning,
b) förhindra dess förekomst och spridning, och
c) om det konstateras förekomst av den, förhindra dess spridning och bekämpa den i syfte att utrota den.
Artikel 2
1. Medlemsstaterna skall varje år genomföra systematiska officiella undersökningar för att kontrollera förekomst av skadegöraren på det förtecknade växtmaterialet med ursprung i deras territorium. För att identifiera andra möjliga smittkällor som hotar produktionen av det förtecknade växtmaterialet skall medlemsstaterna göra en riskbedömning och, om ingen risk för spridning av skadegöraren har konstaterats under den bedömningen skall de, i produktionsområdena för det förtecknade växtmaterialet, genomföra riktade officiella undersökningar för att kontrollera förekomst av skadegöraren på andra växter än det förtecknade växtmaterialet, även på vilda värdväxter av familjen Solanaceae samt på ytvatten som används för bevattning eller duschning av det förtecknade växtmaterialet och på flytande avfall som släpps ut från anläggningar för industriell bearbetning eller förpackning där det förtecknade växtmaterialet hanteras och som används för bevattning och duschning av det förtecknade växtmaterialet. Omfattningen av dessa riktade undersökningar skall bestämmas med beaktande av den konstaterade risken. Medlemsstaterna kan också utföra officiella undersökningar för att kontrollera förekomst av skadegöraren på annat material, t.ex. odlingssubstrat, jord och fast avfall från anläggningar för industriell bearbetning eller förpackning.
2. De officiella undersökningar som anges i punkt 1 skall genomföras
a) på det förtecknade växtmaterialet i enlighet med de uppgifter som anges i punkt 1 i avsnitt II i bilaga I,
b) på värdväxter som inte återfinns i det förtecknade växtmaterialet och på vatten, inklusive flytande avfall, i enlighet med lämpliga metoder, och stickprov skall, när så är lämpligt, tas och genomgå officiella eller officiellt övervakade laboratorietest, och
c) när så är lämpligt på annat material i enlighet med lämpliga metoder.
Ytterligare uppgifter om besiktningarna och om stickprovernas antal, ursprung och inledning samt om tidpunkten för deras insamling skall för dessa undersökningar beslutas av de ansvariga officiella organen enligt direktiv 77/93/EEG, på grundval av sunda vetenskapliga och statistiska principer och skadegörarens biologiska egenskaper samt med beaktande av de berörda medlemsstaternas särskilda produktionssystem för det förtecknade växtmaterialet och, i förekommande fall, för skadegörarens andra värdväxter.
3. Resultaten av och detaljerna i fråga om de officiella undersökningar som fastställs i punkt 1 skall varje år anmälas till de andra medlemsstaterna och till kommissionen i enlighet med bestämmelserna i punkt 2 i avsnitt II i bilaga I. Dessa anmälningar skall göras senast den 1 juni, med undantag av anmälningar om utsädespotatis som skall ges in före den 1 september. Detaljerna och resultaten ifråga om grödor skall avse föregående års produktion. Innehållet i dessa anmälningar kan överlämnas till kommittén.
4. Följande bestämmelse skall antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
- De lämpliga metoderna för de undersökningar och laboratorietest som avses i punkt 2 första stycket under b.
5. Följande bestämmelser får antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
- De lämpliga metoderna för de undersökningar som avses i punkt 2 första stycket under c.
- Närmare uppgifter om de undersökningar som avses i punkt 2 andra stycket, för att säkerställa jämförbara nivåer på medlemsstaternas garantier.
Artikel 3
Medlemsstaterna skall säkerställa att misstänkt förekomst eller bekräftad närvaro av skadegöraren på deras territorium rapporteras till deras egna ansvariga officiella organ.
Artikel 4
1. Vid varje fall av misstänkt förekomst av skadegöraren skall de ansvariga officiella organen i den berörda medlemsstaten eller de berörda medlemsstaterna säkerställa att officiella eller officiellt övervakade laboratorietest genomförs på det förtecknade växtmaterialet enligt den lämpliga metod som anges i bilaga II och enligt de villkor som anges i punkt 1 i bilaga III, eller, i andra fall, någon annan officiellt godkänt metod, för att bekräfta eller vederlägga den misstänkta förekomsten. Om misstanken bekräftas skall de krav som fastställs i punkt 2 i bilaga III gälla.
2. I avvaktan på bekräftelse eller vederläggande av misstänkt förekomst enligt punkt 1, i varje enskilt fall av misstänkt förekomst där antingen
i) de sjukdomssymptom som orsakas av skadegöraren har diagnostiserats och ett eller flera snabbscreeningtest har genomförts med positivt resultat på sätt som anges i avsnitt I punkt 1 och avsnitt II i bilaga II, eller
a) förbjuda flyttning av plantor och knölar från alla grödor, partier eller sändningar från vilka stickproven har tagits, förutom då det sker under deras övervakning och förutsatt att det har konstaterats att det inte finns någon identifierbar risk för att skadegöraren skall spridas,
b) vidta åtgärder för att spåra den misstänkta förekomstens ursprung,
c) införa lämpliga ytterligare försiktighetsåtgärder på grundval av hur stor risken bedöms vara, särskilt i förhållande till produktionen av det förtecknade växtmaterialet och flyttning av andra partier av utsädespotatis än sådana som avses under a, som har producerats på den odlingsplats där de stickprov, som avses under a, har tagits, för att hindra att skadegöraren på något sätt sprids.
3. I fall av misstänkt förekomst av skadegöraren skall, om det finns risk för angrepp på det förtecknade växtmaterialet eller ytvattnet från eller till en annan medlemsstat, den medlemsstat där misstanken har rapporterats omedelbart till den eller de andra berörda medlemsstaterna, beroende på den konstaterade risken, anmäla den nämnda misstänkta förekomsten, och de nämnda medlemsstaterna skall då samarbeta på lämpligt sätt. Den eller de medlemsstater som fått anmälan skall vidta försiktighetsåtgärder enligt punkt 2 c och i förekommande fall vidta ytterligare åtgärder enligt punkterna 1 och 2.
4. Följande bestämmelse får antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
- De åtgärder som anges i punkt 2 c.
Artikel 5
1. Om ett officiellt eller officiellt övervakat laboratorietest som, med avseende på det förtecknade växtmaterialet, använder den lämpliga metod som anges i bilaga II, eller i andra fall, någon annan officiellt godkänd metod, bekräftar skadegörarens förekomst i ett stickprov som tagits på grund av detta direktiv, skall de ansvariga officiella organen i en medlemsstat, med beaktande av sunda vetenskapliga principer, skadegörarens biologiska egenskaper och de särskilda systemen för produktion, marknadsföring och bearbetning av skadegörarens värdväxt i den medlemsstaten,
a) i fråga om det förtecknade växtmaterialet vidta följande åtgärder:
i) Genomföra en utredning för att, i enlighet med bestämmelserna i bilaga IV, fastställa angreppets omfattning och dess primärkälla eller -källor, med ytterligare test i enlighet med artikel 4.1 på åtminstone alla lager av utsädespotatis ur kloner som är närbesläktade.
ii) Förklara följande angripet: Det förtecknade växtmaterialet, sändningen och/eller partiet som stickprovet togs från, maskinerna, fordonet, fartyget, lagret, eller delar av dessa, och alla andra föremål, inklusive förpackningsmaterialet som har varit i kontakt med det förtecknade växtmaterial från vilket stickprovet togs. I förekommande fall även förklara följande som angripet: Det eller de fält, den eller de enheter för skyddad växtproduktion och den eller de produktionsplatser där det förtecknade växtmaterialet har skördats och från vilka stickprovet tagits. I fråga om de stickprov som tagits under växtsäsongen förklara följande för angripet: Det eller de fält, den eller de produktionsplatser, och i förekommande fall den eller de enheter för skyddad växtproduktion som stickprovet togs ifrån.
iii) I enlighet med bestämmelserna i punkt 1 i bilaga V fastställa omfattningen av troliga angrepp genom kontakt före eller efter skörd, genom produktionsmässig anknytning, bevattning eller duschning eller genom klonsläktskap med det angivna angreppet.
iv) Avgränsa ett område på grundval av förklaringen om angreppet enligt punkt ii, fastställa omfattningen av det troliga angreppet enligt punkt iii och skadegörarens möjliga spridning, i enlighet med bestämmelserna i punkt 2 i i bilaga V.
b) I fråga om grödor från värdväxter som inte nämns under a, då det har konstaterats att det finns en risk vid produktionen av det förtecknade växtmaterialet vidta följande åtgärder:
i) Genomföra en utredning i enlighet med punkt a i.
ii) Förklara de av skadegörarens värdväxter som provet har tagits från för angripna.
iii) Fastställa det troliga angreppet och avgränsa ett område i enlighet med punkterna a iii respektive a iv i förhållande till produktionen av det förtecknade växtmaterialet.
c) I fråga om ytvatten (även flytande avfall från anläggningar för industriell bearbetning eller förpackning där det förtecknade växtmaterialet hanteras) och besläktade vilda värdväxter av familjen Solanaceae, då det har konstaterats att produktionen av det förtecknade växtmaterialet utgör en risk genom bevattning, duschning eller översvämning med ytvattnet vidta följande åtgärder:
i) Genomföra en utredning som omfattar en officiell undersökning vid lämpliga tidpunkter på prov av ytvattnet och, om sådana finns, på vilda värdväxter av familjen Solanaceae för att fastställa angreppets omfattning.
ii) Förklara det ytvatten som provet eller proven har tagits från för angripet i den utsträckning som det är lämpligt och på grundval av undersökningen enligt punkt i.
iii) Fastställa det troliga angreppet och avgränsa ett område på grundval av förklaringen om angreppet enligt punkt ii och skadegörarens möjliga spridning med beaktande av bestämmelserna i punkt 1 och 2 ii i bilaga V.
2. Medlemsstaterna skall, i enlighet med bestämmelserna i punkt 3 i bilaga V, omedelbart till de andra medlemsstaterna och till kommissionen anmäla varje angrepp som fastställs enligt punkterna 1 a ii och 1 c ii och uppgifterna om avgränsning av områden enligt punkt 1 a iv och, där så är tillämpligt, enligt punkt 1 c iii. Innehållet i denna anmälan enligt detta stycke får överlämnas till kommittén.
Medlemsstaterna skall samtidigt till kommissionen överlämna en tilläggsanmälan enligt 3 a i bilaga V. Innehållet i denna anmälan enligt detta stycke skall omedelbart överlämnas till kommitténs ledamöter.
3. Till följd av den anmälan som avses i punkt 2 och dess beståndsdelar, skall de andra medlemsstater som anges i anmälan genomföra en utredning i enlighet med punkt 1 a i och, där så är tillämpligt, punkt 1 c i och om så är lämpligt vidta ytterligare åtgärder i enlighet med punkterna 1 och 2.
Artikel 6
1. Medlemsstaterna skall föreskriva att det förtecknade växtmaterial som förklarats för angripet enligt artikel 5.1 a ii inte får planteras och att det, under övervakning av och med godkännande av deras ansvariga officiella organ, skall underkastas någon av bestämmelserna i punkt 1 i bilaga VI, så att det kan fastställas att det inte finns någon identifierbar risk för att skadegöraren sprids.
2. Medlemsstaterna skall föreskriva att det förtecknade växtmaterial som förklarats troligen angripet enligt artikel 5.1 a iii och 5.1 c iii inbegripet det förtecknade växtmaterial för vilket en risk har konstaterats föreligga, och som producerats på produktionsplatser som förklarats troligen angripna enligt artikel 5.1 a iii inte får planteras och att det, under övervakning av deras ansvariga officiella organ, skall användas på lämpligt sätt eller bortförskaffas enligt punkt 2 i bilaga VI, så att det kan fastställas att det inte finns någon identifierbar risk för att skadegöraren sprids.
3. Medlemsstaterna skall föreskriva att alla maskiner, fordon, fartyg, lager, eller delar av dessa, och alla andra föremål, inklusive förpackningsmaterial, som har förklarats angripna enligt artikel 5.1 a ii eller förklarats troligen angripna enligt artikel 5.1 a iii och 5.1 c iii, antingen skall förstöras eller saneras med lämpliga metoder som fastställs i punkt 3 i bilaga VI. Efter saneringen skall inga sådana föremål längre betraktas som angripna.
4. Utan att det påverkar tillämpningen av de åtgärder som genomförs enligt punkterna 1 3 skall medlemsstaterna föreskriva att ett antal åtgärder skall genomföras enligt punkterna 4.1 och 4.2 i bilaga VI inom det område som avgränsas enligt artikel 5.1 a iv och 5.1 c iii. Uppgifter om dessa åtgärder skall varje år anmälas till de andra medlemsstaterna och till kommissionen. Innehållet i denna anmälan för överlämnas till kommittén.
Artikel 7
1. Medlemsstaterna skall föreskriva att utsädespotatis skall uppfylla kraven i direktiv 77/93/EEG och att de i direkt led skall härstamma ur potatismaterial som erhållits enligt ett officiellt godkänt program och som har konstaterats vara fritt från skadegöraren vid officiella eller officiellt övervakade tester då den lämpliga metod, som anges i bilaga II, har använts.
De ovannämnda testerna skall utföras av en medlemsstat
a) i de fall då bekräftade fynd av skadegöraren har gjorts i dess egen produktion av utsädespotatis
i) genom tester av tidigare generationer inklusive det ursprungliga klonurvalet och systematiska tester av det ursprungliga klonurvalet av utsädespotatisen, eller
ii) genom tester av allt ursprungligt klonurval av utsädespotatis eller tidigare generationer inklusive det ursprungliga klonurvalet i de fall då inget släktskap genom klon har påvisats och
b) i andra fall, antingen av varje planta i det ursprungliga klonurvalet eller av representativa stickprov av basutsädespotatis eller tidigare generationer.
2. Följande bestämmelser får antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
- Tillämpningsföreskrifterna i punkt 1, andra stycket, punkt a.
- De bestämmelser om representativa stickprov som föreskrivs i punkt 1, andra stycket, punkt b.
Artikel 8
Medlemsstaterna skall förbjuda innehav och hantering av skadegöraren.
Artikel 9
Utan att det påverkar tillämpningen av bestämmelserna i direktiv 77/93/EEG får bestämmelserna bevilja undantag från de åtgärder som avses i artiklarna 6 och 8 i det här direktivet i enlighet med bestämmelserna i direktiv 95/44/EG i experimentellt eller vetenskapligt syfte och för växtförädling (5).
Artikel 10
Artikel 11
Ändringar i bilagorna till detta direktiv mot bakgrund av nya vetenskapliga eller tekniska rön skall antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG. När det gäller de metoder som anges i bilaga II och åtgärderna i punkt 4.1 och 4.2 i bilaga VI till detta direktiv, skall kommissionen förbereda en rapport där metoderna och åtgärderna granskas mot bakgrund av gjorda erfarenheter som vunnits, och rapporten skall överlämnas till kommittén före den 1 januari 2002.
Artikel 12
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 21 augusti 1999. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning till detta direktiv när de offentliggörs. Närmare föreskrifter för hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall omedelbart till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv. Kommissionen skall underrätta de övriga medlemsstaterna om detta.
Artikel 13
RÅDETS DIREKTIV 98/93/EG av den 14 december 1998 om ändring av direktiv 68/414/EEG om en skyldighet för medlemsstaterna i EEG att inneha minimilager av råolja och/eller petroleumprodukter
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 103 a.1 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
av följande skäl: (1) Den 20 december 1968 antog rådet direktiv 68/414/EEG om en skyldighet för medlemsstaterna i EEG att inneha minimilager av råolja och/eller petroleumprodukter (4).
(2) Råolja och petroleumprodukter som importeras spelar fortfarande en viktig roll i gemenskapens energiförsörjning. Varje svårighet, även om den är tillfällig, som leder till att leveranserna av dessa produkter begränsas, eller till att deras pris stiger avsevärt på de internationella marknaderna skulle kunna orsaka allvarliga störningar i gemenskapens ekonomiska verksamhet. Gemenskapen måste därför vara i stånd att upphäva eller åtminstone minska de skadeverkningar som skulle kunna uppstå i sådana fall. Det är nödvändigt att uppdatera direktiv 68/414/EEG så att det anpassas till den verklighet som råder på gemenskapens inre marknad och till utvecklingen på oljemarknaderna.
(3) Genom direktiv 73/238/EEG (5) fattade rådet beslut om lämpliga åtgärder - däribland uttag ur oljelager - som skall vidtas om det uppstår svårigheter i fråga om försörjningen av råolja och petroleumprodukter till gemenskapen. Medlemsstaterna har åtagit sig liknande skyldigheter i avtalet om ett "Internationellt energiprogram".
(4) Det är viktigt att öka försörjningssäkerheten för olja.
(5) Lagerhållningen av olja måste vara så organiserad att den inte förhindrar att den inre marknaden fungerar väl.
(6) Bestämmelserna i detta direktiv påverkar inte den fullständiga tillämpningen av fördraget, särskilt bestämmelserna om den inre marknaden och konkurrens.
(7) I enlighet med subsidiaritetsprincipen och proportionalitetsprincipen fastställd i artikel 3b i fördraget går det lättare att på gemenskapsnivå uppnå målet att upprätthålla en hög nivå av försörjningssäkerhet för olja i gemenskapen genom säkra system, som är öppna för insyn och som bygger på solidaritet mellan medlemsstaterna, och som samtidigt uppfyller bestämmelserna om den inre marknaden och om konkurrens. Detta direktiv sträcker sig inte utöver vad som behövs för att uppnå detta mål.
(8) Lagren måste stå till medlemsstaternas förfogande om det uppstår svårigheter med oljeförsörjningen. Medlemsstaterna bör ha befogenhet och möjlighet att kontrollera användningen av lagren så att de utan dröjsmål kan göras tillgängliga för de områden där behovet av oljeleveranser är störst.
(9) Lagerhållningen bör vara så organiserad att lagrens tillgänglighet och förbrukarnas tillgång till lagren säkerställs.
(10) Lagerhållningssystemen bör bygga på öppenhet för insyn för att säkerställa att den börda som lagerhållningsskyldigheten innebär fördelas rättvist och utan någon diskriminering. Medlemsstaterna kan göra information om kostnaden för att hålla oljelager tillgänglig för berörda parter.
(11) I syfte att organisera lagerhållningen får medlemsstaterna använda sig av ett system med ett lagerhållande organ eller en enhet som skall förvalta alla eller en del av de lager som utgör lagerhållningsskyldigheten. Eventuell överskjutande del bör hållas av raffinaderier och andra marknadsaktörer. Partnerskap mellan staten och branschen är nödvändigt för att lagerhållningssystemen skall fungera effektivt och säkert.
(12) En inhemsk utvinning bidrar i sig till försörjningssäkerhet. För medlemsstater med inhemsk oljeutvinning kan utvecklingen på oljemarknaden motivera ett lämpligt undantag från skyldigheten att hålla oljelager. I enlighet med subsidiaritetsprincipen får medlemsstaterna befria företag från skyldigheten att hålla lager i en omfattning som inte överstiger den kvantitet produkter som dessa företag framställer från råolja som utvunnits i medlemsstaten.
(13) Det är lämpligt att tillämpa tillvägagångssätt som gemenskapen och medlemsstaterna redan följer inom ramen för sina internationella skyldigheter och avtal. På grund av förändringar i oljeförbrukningsmönstret har flygbränsle för internationell luftfart blivit ett viktigt inslag i denna förbrukning.
(14) Det finns ett behov av att anpassa och förenkla gemenskapens system för statistisk rapportering av oljelager.
(15) Oljelager kan i princip hållas var som helst i gemenskapen och därför är det lämpligt att göra det enklare att upprätta lager utanför det nationella territoriets gränser. Det är nödvändigt att beslut om att hålla lager utanför det nationella territoriets gränser fattas av den berörda medlemsstatens regering i enlighet med dess behov och med hänsyn till försörjningssäkerheten. För lager som hålls tillgängliga för andra företag eller organ/enheter behövs utförligare bestämmelser för att garantera att de är tillgängliga och åtkomliga vid händelse av oljeförsörjningssvårigheter.
(16) För att säkerställa att den inre marknaden fungerar smidigt är det önskvärt att främja användningen av avtal mellan medlemsstater när det gäller minimilagerhållning för att främja användningen av lageranläggningar i andra medlemsstater. Beslut att ingå sådana avtal skall fattas av de berörda medlemsstaterna.
(17) Det är lämpligt att bygga ut den administrativa tillsynen av lagren och att inrätta verkningsfulla system för kontroll och verifiering av lagren. Införandet av ett sådant kontrollsystem kräver ett sanktionssystem.
(18) Genom direktiv 72/425/EEG ökades den referenstid som anges i artikel 1 första stycket i direktiv 68/414/EEG från 65 till 90 dagar och villkor för genomförandet av denna utökning fastlades. Det direktivet har gjorts obsolet genom det här direktivet. Direktiv 72/425/EEG bör därför upphävas.
(19) Det är lämpligt att med jämna mellanrum informera rådet om läget beträffande beredskapslagren i gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 68/414/EEG ändras på följande sätt:
1. Medlemsstaterna skall anta de lagar och andra författningar som är lämpliga för att, om inte annat följer av bestämmelserna i artikel 7, inom gemenskapen, alltid hålla sina lager av petroleumprodukter på en nivå som för varje typ av petroleumprodukter, enligt förteckningen i artikel 2, motsvarar minst 90 dagars genomsnittlig, daglig inhemsk förbrukning under det föregående kalenderåret enligt artikel 4.
2. Den del av den inhemska förbrukningen som täcks av petroleumprodukter baserade på utvinning inom den berörda medlemsstaten får dras av upp till högst 25 % från nämnda förbrukning. Fördelningen inom medlemsstaterna av resultatet av ett sådant avdrag skall beslutas av den berörda medlemsstaten." 2. Artikel 2 skall utgå.
3. Nuvarande artikel 3 skall betecknas artikel 2 och skall kompletteras med följande stycke:
3. För att kunna uppfylla kraven i punkterna 1 och 2 får medlemsstaterna besluta att använda sig av ett lagerhållande organ eller en enhet med ansvar för att hålla alla lagren eller en del av dessa.
"Artikel 4
Medlemsstaterna skall till kommissionen överlämna ett statistiskt sammandrag över de lager som finns i slutet av varje månad, upprättat enligt artiklarna 5 och 6 och med närmare angivande av antalet dagar med genomsnittlig förbrukning under det föregående kalenderåret som dessa lager representerar. Detta sammandrag skall överlämnas senast den tjugofemte dagen i den andra månaden efter den månad som sammandraget avser.
En medlemsstats lagerhållningsskyldighet skall baseras på det föregående kalenderårets inhemska förbrukning. Vid början av varje kalenderår skall medlemsstaterna göra en ny beräkning av sin lagerhållningsskyldighet senast den 31 mars varje år och säkerställa att de uppfyller sina nya skyldigheter så snart som möjligt och i vart fall senast den 31 juli varje år.
I det statistiska sammandraget skall lager av jetbränsle av fotogentyp särredovisas under kategori II." 6. Artikel 5 skall ersättas med följande:
"Artikel 5
Obligatoriska lager enligt artikel 1 får hållas i form av råolja, halvfabrikat och färdiga produkter.
I det statistiska sammandraget av lagren som föreskrivs i artikel 4, skall färdiga produkter redovisas efter sin verkliga vikt. Råolja och halvfabrikat skall redovisas
- fördelade i förhållande till de kvantiteter av varje produktkategori som erhållits under föregående kalenderår från den berörda statens raffinaderier, eller
- på grundval av raffinaderiernas produktionsprogram i den berörda staten under innevarande år, eller
- på grundval av förhållandet mellan den totala kvantitet som tillverkats under föregående kalenderår i den berörda staten av de produkter som omfattas av lagringsskyldigheten och den totala mängd råolja som använts under det året. Det föregående skall gälla högst 40 % av den totala lagringsskyldigheten för de första och andra kategorierna (motorbensin och tunn eldningsolja) och högst 50 % för den tredje kategorin (tjocka eldningsoljor).
Blandningsprodukter får, när de är avsedda för bearbetning till de färdiga produkter som anges i artikel 2, tjäna som ersättning för de produkter för vilka de är avsedda." 7. Artikel 6 skall ändras enligt följande:
a) Punkt 1 skall ersättas med följande:
"1. Vid beräkning av nivån på de minimilager som föreskrivs i artikel 1 skall endast de kvantiteter räknas in i det statistiska sammandraget som hålls i enlighet med artikel 3.1". b) Punkt 2 skall ersättas med följande:
"2. För genomförandet av detta direktiv får lager, enligt avtal mellan regeringar, upprättas inom en medlemsstats territorium för företag eller organ/enheter som är etablerade i en annan medlemsstat. Beslut om att hålla en del av sina lager utanför sitt nationella territorium skall fattas av den berörda medlemsstatens regering.
I dessa fall skall den medlemsstat på vars territorium lagren hålls inom ramen för ett sådant avtal inte hindra att dessa lager överförs till de andra medlemsstaterna, för vars räkning lagren hålls enligt avtalet. Den skall kontrollera dessa lager i enlighet med förfarandena som närmare anges i det avtalet men inte räkna in dem i sitt statistiska sammandrag. Den medlemsstat för vars räkning lagren hålls får räkna in dem i sitt statistiska sammandrag.
I dessa fall skall varje medlemsstat, tillsammans med det statistiska sammandrag som föreskrivs i artikel 4, överlämna en rapport till kommissionen om de lager som hålls på medlemsstatens eget territorium till förmån för en annan medlemsstat, liksom om de lager som hålls i andra medlemsstater till dess egen förmån. I båda fallen skall rapporten innehålla uppgift om var lagren är belägna och/eller om de företag som håller lagren, lagrade kvantiteter och produktkategorier - eller uppgift om att det rör sig om råolja.
Utkast till de avtal som nämns i första stycket skall överlämnas till kommissionen, som får lämna sina kommentarer till de berörda regeringarna. När avtalen väl har ingåtts skall de anmälas till kommissionen, som skall underrätta de övriga medlemsstaterna om dem.
Avtalen skall uppfylla följande villkor:
- De skall avse råolja samt alla petroleumprodukter som omfattas av detta direktiv.
- De skall fastställa villkor och tillvägagångssätt för lagerhållning som är inriktade på att trygga kontrollen av lagren och deras tillgänglighet.
- De skall närmare ange de förfaranden som skall användas för att kontrollera och identifiera de lager som föreskrivs, bland annat metoder för att utföra inspektioner och för samarbetet under dessa.
- De skall normalt gälla under obegränsad tid.
- De skall, om en part kan säga upp avtalet, föreskriva att sådan uppsägning inte skall gälla i händelse av en försörjningskris och att kommissionen under alla förhållanden skall erhålla förhandsinformation om uppsägning sker.
När lager, upprättade enligt sådana avtal, inte ägs av det företag, det organ/enhet som har skyldighet att hålla lager, utan hålls tillgängliga för företaget, organet/enheten av ett annat företag, organ/enhet, skall följande villkor uppfyllas:
- Det företag, organ eller den enhet som har rätt till lagren skall ha kontraktsenlig rätt att förvärva dessa lager under avtalsperioden. Sättet att fastställa priset för detta förvärv skall överenskommas mellan de berörda parterna.
- Minsta avtalsperiod skall vara 90 dagar.
- Uppgifter om var lagren är belägna och/eller om de företag som håller lagren tillgängliga för det företag, organ/enhet som har rätt till dem, liksom lagrade kvantiteter och produktkategorier eller uppgift om att det rör sig om lagrad råolja, skall anges.
- Den faktiska tillgången till lagren för det företag, organ/enhet som har rätt till dem måste, när som helst under avtalsperioden, garanteras av det företag, organ/enhet som håller lagren tillgängliga för det företag, organ eller den enhet som har rätt till dem.
- Det företag, organ/enhet som håller lagren för det företag, organ/enhet som har rätt till dem, skall vara underkastad lagstiftningen i den medlemsstat på vars territorium lagren befinner sig, när det gäller den medlemsstatens lagliga befogenheter att kontrollera och verifiera förekomsten av lagren." c) Punkt 3 andra stycket skall ersättas med följande:
"Följaktligen skall särskilt följande uteslutas från det statistiska sammandraget: inhemsk råolja som ännu inte utvunnits, mängder som skall användas till bunkring för havsgående fartyg, mängder i direkt transitering, frånsett de i punkt 2 angivna lagren, mängder i rörledningar, tankbilar och tankvagnar på järnväg, i lagertankar på detaljistmarknaden samt hos små förbrukare. De mängder som innehas av de väpnade styrkorna och de som innehas av oljebolag för deras räkning skall också uteslutas från det statistiska sammandraget." 8. Följande artikel skall införas:
"Artikel 6a
Medlemsstaterna skall anta alla bestämmelser som är nödvändiga och vidta alla åtgärder som är nödvändiga för att säkerställa kontrollen och övervakningen av lagren. De skall inrätta system för verifiering av lagren i enlighet med bestämmelserna i detta direktiv."
9. Följande artikel skall införas:
"Artikel 6b
Medlemsstaterna skall bestämma vilka straff som skall gälla för överträdelser av de nationella bestämmelser som antas i enlighet med detta direktiv och vidta alla åtgärder som är nödvändiga för att säkerställa genomförandet av dessa bestämmelser. Straffen skall vara effektiva, proportionerliga och avskräckande."
Artikel 2
Direktiv 72/425/EEG skall upphävas med verkan från och med den 31 december 1999.
Artikel 3
1. Medlemsstaterna skall före den 1 januari 2000 sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 4
På grund av Hellenska republikens särskilda situation garanteras den en ej förnybar extra period på tre år för att tillämpa detta direktivs skyldigheter vad gäller att låta mängder som används till bunkring av internationellt flyg ingå när det gäller att beräkna inhemsk förbrukning.
Artikel 5
Kommissionen skall regelbundet till rådet överlämna en rapport om läget beträffande lagren i gemenskapen, inbegripet, när så är lämpligt, om behovet av en harmonisering för att säkerställa en effektiv kontroll och övervakning av lagren. Den första rapporten skall överlämnas till rådet under det andra året efter det datum som fastställs i artikel 3.1.
Artikel 6
KOMMISSIONENS FÖRORDNING (EG) nr 121/98 av den 16 januari 1998 om ändring av bilagorna I, II och III i rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (1), senast ändrad genom kommissionens förordning (EG) nr 1850/97 (2), särskilt artikel 6, 7 och 8 i denna, och med beaktande av följande:
I enlighet med förordning (EEG) nr 2377/90 måste gränsvärden för högsta tillåtna restmängder successivt fastställas för samtliga farmakologiskt verksamma substanser som används inom gemenskapen i veterinärmedicinska läkemedel som är avsedda att ges till livsmedelsproducerande djur.
Gränsvärden bör fastställas först efter det att Kommittén för veterinärmedicinska läkemedel har granskat all relevant information beträffande säkerheten med restmängder av ämnet i fråga för den som konsumerar livsmedel med animaliskt ursprung samt restmängdernas påverkan på den industriella bearbetningen av livsmedel.
Vid fastställandet av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung är det nödvändigt att ange de djurarter i vilka restmängder kan förekomma, vilka mängder som kan förekomma i var och en av de relevanta vävnaderna från det behandlade djuret (målvävnad) samt vilket slag av restmängd som är relevant vid övervakningen av restmängder (restmarkör).
För kontroll av resthalter bör enligt tillämplig gemenskapslagstiftning gränsvärden vanligtvis fastställas för målvävnaderna lever eller njure. I den internationella handeln avlägsnas dock ofta lever och njure från slaktkroppen, och gränsvärden bör därför alltid fastställas även för muskel- eller fettvävnader.
För veterinärmedicinska läkemedel som är avsedda för äggläggande fåglar, mjölkdjur eller honungsbin, måste gränsvärden även fastställas för ägg, mjölk eller honung.
Danofloxacin, cefazolin och trimetoprim skall införas i bilaga I till förordning (EEG) nr 2377/90.
Lini oleum, folsyra, betain och cefazolin skall införas i bilaga II till förordning (EEG) nr 2377/90.
För att möjliggöra komplettering av vetenskapliga studier, bör giltighetstiden för temporära MRL, tidigare definierad i bilaga III i förordning (EEG) nr 2377/90, förlängas för penetamat.
En tidsfrist på 60 dagar bör tillåtas innan denna förordning träder i kraft så att medlemsstaterna kan göra de nödvändiga anpassningarna till bestämmelserna i denna förordning av tillstånden att släppa ut de berörda veterinärmedicinska läkemedlen på marknaden, vilka beviljats enligt rådets direktiv 81/851/EEG (3), senast ändrat genom direktiv 93/40/EEG (4).
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I, II och III till förordning (EEG) nr 2377/90 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den kraft den sextionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 179/98 av den 23 januari 1998 om ändring av rådets förordning (EG) nr 3051/95 om säkerhetsorganisation för roll-on/roll-off-passagerarfartyg (ro-ro-fartyg)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 3051/95 av den 8 december 1995 om säkerhetsorganisation för roll-on/roll-off-passagerarfartyg (ro-ro-fartyg) (1), särskilt artikel 9 i denna, och
med beaktande av följande: I förordning (EG) nr 3051/95 föreskrivs att företag och medlemsstater skall följa bestämmelserna i Internationella säkerhetsorganisationskoden, som antogs av Internationella sjöfartsorganisationen (IMO) genom församlingens resolution A.741 (18) av den 4 november 1993, för ro-ro-fartyg i trafik till eller från hamnar i medlemsstater inom gemenskapen.
För att säkerställa ett enhetligt genomförande av Internationella säkerhetsorganisationskoden (ISM), antog IMO genom resolution A.788 (19) av den 23 november 1995 riktlinjer om myndigheters genomförande av Internationella säkerhetsorganisationskoden (ISM-koden).
Det är nödvändigt att ta hänsyn till utvecklingen på det internationella planet genom att införa närmare bestämmelser om utfärdandet av interimistiska dokument och certifikat, formulär för ISM-dokument och ISM-certifikat samt vissa standarder avseende ISM-certifieringsarrangemang.
Det är lämpligt att säkerställa att giltigheten för vissa dokument och certifikat som redan utfärdats inte påverkas.
Förordning (EG) nr 3051/95 bör ändras till följd av detta.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som inrättats enligt artikel 12 i rådets direktiv 93/75/EEG (2), senast ändrat genom kommissionens direktiv 97/34/EG (3).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 496/98 av den 27 februari 1998 om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 2509/97 (2), särskilt artikel 9 i denna, och med beaktande av följande:
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från sektionen för tulltaxe- och statistiknomenklatur inom tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 539/98 av den 9 mars 1998 medförande ändring av förordning (EEG) nr 3077/78 om godkännande av intyg för humle som importeras från tredje land som likvärdiga med gemenskapsintyg
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1696/71 av den 26 juli 1971 om den gemensamma organisationen av marknaden för humle (1), senast ändrad genom förordning (EG) nr 1554/97 (2), särskilt artikel 5.2 i denna, och
med beaktande av följande: Genom kommissionens förordning (EEG) nr 3077/78 (3), senast ändrad genom förordning (EG) nr 2132/95 (4), godkänns intyg för humle som importeras från vissa tredje länder såsom likvärdiga med gemenskapsintygen samt upprättas en förteckning över de förvaltningar i dessa länder som har befogenhet att utfärda likvärdiga intyg, liksom en förteckning över de produkter som omfattas. Till följd av de uppgifter som Polen har lämnat in är det nödvändigt att ändra bilagan till förordning (EEG) nr 3077/78.
Det åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för humle.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till denna förordning skall ersätta bilagan till förordning (EEG) nr 3077/78.
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 726/98 av den 31 mars 1998 om ändring av förordning (EG) nr 2543/95 om tillämpningsföreskrifter för ordningen med exportlicenser inom olivoljesektorn
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter (1), senast ändrad genom förordning (EG) nr 1581/96 (2), särskilt artiklarna 2 och 3 i denna, och
med beaktande av följande: I kommissionens förordning (EG) nr 2543/95 (3), ändrad genom förordning (EG) nr 2126/96 (4), föreskrivs särskilda tillämpningsföreskrifter för ordningen med exportlicenser inom olivoljesektorn. För att förbättra det sätt på vilket ordningen fungerar bör vissa särskilda tillämpningsföreskrifter fastställas för licenser utan förutfastställelse av bidraget, bl.a. vad gäller säkerhetsbeloppet och ordningen för inlämnande av ansökningar och utfärdande av licenser. Erfarenheten visar att det också är lämpligt att anpassa beloppet för säkerheten liksom tidsfristen både för inlämnandet av licensansökningar och för utfärdandet av dessa. Det är lämpligt att föreskriva att de åtgärder som vidtas när det finns risk för att de normala avsättningskvantiteterna överskrida endast får gälla exportlicenser med förutfastställelse av bidraget. För att på ett bättre sätt kunna följa exportförloppet måste de upplysningar medlemsstaterna skall lämna in preciseras.
Enligt artikel 5.1 fjärde strecksatsen i kommissionens förordning (EEG) nr 3719/88 av den 16 november 1988 om gemensamma tillämpningsföreskrifter för systemet med import- och exportlicenser och förutfastställelselicenser för jordbruksprodukter (5), senast ändrad genom förordning (EG) nr 1404/97 (6), krävs ingen licens för export vid en säkerhet på högst 5 ecu. Det låga säkerhetsbeloppet för export utan bidrag innebär att mycket skulle kunna exporteras utan licens, vilket skulle försvaga kontrollen av kvantiteterna i fråga. För att undvika den risken bör särskilda villkor gälla i nämnda fall.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för oljor och fetter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 2543/95 ändras på följande sätt:
1. I artikel 2.2 skall "elva" ersättas med "tolv".
2. Artikel 2 skall ändras på följande sätt:
1. Punkt 3 skall ersättas med följande:
"3. Beloppet för säkerheten för exportlicenserna skall fastställas till
a) 10 ecu per 100 kg netto för licenser med förutfastställelse av bidraget,
b) 1 ecu per 100 kg netto i övriga fall."
2. Följande punkt skall läggas till:
"4. Genom undantag från artikel 5.1 fjärde strecksatsen i förordning (EEG) nr 3719/88 skall ingen licens krävas vid export av en kvantitet på 50 kg eller mindre."
3. Artikel 3 skall ändras på följande sätt:
1. Punkt 1 skall ersättas med följande:
"1. Ansökningar om exportlicenser med förutfastställelse av bidraget skall inlämnas hos den behöriga myndigheten från och med tisdag till och med torsdag varje vecka. Ansökningar som inlämnas en måndag eller fredag skall behandlas som om de vore inlämnade närmast följande tisdag."
2. Första stycket i punkt 2 skall ersättas med följande:
"2. Exportlicenserna med förutfastställelse av bidraget skall utfärdas första arbetsdagen från och med tisdagen den vecka som följer efter den period som avses i punkt 1, såvida inte kommissionen under tiden har vidtagit någon av de särskilda åtgärder som avses i punkt 3."
3. Den sista meningen i punkt 3 skall ersättas med följande:
"Dessa åtgärder skall gälla exportlicenser med förutfastställelse av bidraget, och får variera mellan produktkoderna i nomenklaturen över exportbidrag för jordbruksprodukter."
4. I artikel 3.5 sista strecksatsen skall "måndagen" ersättas med "tisdagen" och följande mening läggas till:
"I de fall den enhetliga procentsatsen för godkännande på under 80 % endast gäller de licenser som är bidragsberättigande, får operatören begära att en licens som inte berättigar till bidrag skall utfärdas inom samma tidsfrist för den kvantitet som inte har godkänts."
5. Följande stycke skall läggas till:
"6. Ansökningarna om exportlicenser utan förutfastställelse av bidraget skall lämnas in till de behöriga myndigheterna från måndag till fredag varje vecka. Licenserna skall utfärdas omedelbart."
4. Artikel 5 skall ändras på följande sätt:
1. I punkt 1 första stycket skall "torsdag" ersättas med "fredag".
2. Punkt 1 a skall ersättas med följande:
"a) de ansökningar om exportlicenser med förutfastställelse av bidraget, vilka har lämnats in från och med tisdag till och med torsdag i enlighet med artikel 3.1."
3. I punkt 1 b skall "måndagen innan" ändras till "från och med föregående period fredag till och med torsdag, med separat angivelse för licenser med förutfastställelse av bidraget i förhållande till licenser utan förutfastställelse av bidraget".
4. I punkt 2 skall den del av meningen som föregår den första strecksatsen ersättas med följande:
"Det meddelande om ansökningar som avses i punkt 1 a och, vad gäller tillämpningen av artikel 3.5 de upplysningar som avses i punkt 1 b, skall innehålla följande:"
5. I punkt 2 tredje strecksatsen skall "i förekommande fall" läggas till framför "tillämplig".
6. I punkt 2 skall följande stycke läggas till:
"Dessa upplysningar skall anges separat om licenser för livsmedelshjälp utfärdas."
7. I punkt 3 skall följande läggas till:
". . . ., och ange det regleringsår under vilket licensen utfärdades."
5. I bilagan skall delarna B och D ersättas med de som anges i bilagan till denna förordning.
Artikel 2
KOMMISSIONENS FÖRORDNING (EG) nr 1011/98 av den 14 maj 1998 om ändring av förordning (EEG) nr 1722/93 om tillämpningsföreskrifter för rådets förordningar (EEG) nr 1766/92 och (EEG) nr 1418/76 om produktionsbidrag inom spannmåls- respektive rissektorn
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1766/92 av den 30 juni 1992 om den gemensamma organisationen av marknaden för spannmål (1), senast ändrad genom kommissionens förordning (EG) nr 923/96 (2), särskilt artikel 7.3 i denna,
med beaktande av rådets förordning (EG) nr 3072/95 av den 22 december 1995 om den gemensamma organisationen av marknaden för ris (3), ändrad genom förordning (EG) nr 192/98 (4), särskilt artikel 7 i denna, och
med beaktande av följande: I kommissionens förordning (EEG) nr 1722/93 av den 30 juni 1993 om tillämpningsföreskrifter för rådet förordningar (EEG) nr 1766/92 och (EEG) nr 1418/76 om produktionsbidrag inom spannmåls- respektive rissektorn (5), senast ändrad genom kommissionens förordning (EG) nr 1516/95 (6), föreskrivs att det vid beräkning av produktionsbidrag skall göras åtskillnad mellan stärkelse av majs, vete, potatis och ris, å ena sidan, och stärkelse av korn och havre, å andra sidan. I praktiken har visat sig att det inte längre är nödvändigt att fastställa ett särskilt belopp för stärkelse av korn och havre, och att det enhetliga bidragsbeloppet hädanefter kan tillämpas på all stärkelse utan risk för att otillbörlig kompensation ges.
Särskilda åtgärder kan förväntas när regleringsåret ändras, vilket innebär att såväl bidragslicensernas giltighetstid som beloppet för det enhetliga bidraget förändras.
För att den särskilda säkerheten skall kunna frisläppas för framför allt förestrad och företrad stärkelse är det lämpligt att fastställa de huvudsakliga krav som måste vara uppfyllda. De särskilda bestämmelser som gäller för dessa produkter bör även fortsättningsvis kompletteras med vissa åtgärder inriktade på effektiviteten i kontroller och på sanktioner i fall då villkoren för bearbetning och användning inte iakttas.
I förordningen förskrivs för närvarande att medlemsstaterna varje månad till kommissionen skall överlämna de statistiska uppgifter som både omfattar de kvantiteter stärkelse som har fått produktionsbidrag och de produkter i vilka stärkelse har använts. Det har blivit uppenbart att detta informationslämnande sker onödigt ofta och att det vore lämpligt att ersätta det med kvartalsvisa meddelanden.
Förvaltningskommittén för spannmål har inte yttrat sig inom den tid som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"Artikel 3
1. När ett bidrag beviljas skall det fastställas en gång i månaden. Om marknadspriserna för majs och/eller vete i gemenskapen eller på världsmarknaden varierar betydligt, får det bidrag som beräknas i enlighet med punkt 2 ändras så att hänsyn tas till sådana svängningar.
2. Bidraget per ton stärkelse av majs, vete, korn, havre, potatis, ris eller brutet ris skall beräknas framför allt på grundval av skillnaden mellan
i) marknadspriset på majs i gemenskapen, giltigt i fem dagar före den dag det fastställs, med hänsyn tagen till priserna för vete, och
ii) genomsnittet av de representativa cif-importpriser för Rotterdam, vilket används för att beräkna importavgiften för majs och som konstaterats under de fem dagar som föregår den första tillämpningsdagen,
multiplicerad med koefficienten 1,60.
3. Det bidrag som skall utbetalas skall beräknas i enlighet med punkt 2 och multipliceras med koefficienten i bilaga II, vilken motsvarar KN-numret för den stärkelse som faktiskt används för att framställa de godkända produkterna.
4. De beslut som föreskrivs i denna artikel skall fattas av kommissionen enligt förfarandet i artikel 23 i förordning (EEG) nr 1766/92."
2) I artikel 6 skall punkterna 3 och 4 ersättas med följande:
"3. Bidragslicensen skall innefatta de upplysningar som anges i artikel 5.2, och dessutom bidragssatsen och den sista dag då licensen är giltig, som skall vara den sista dagen i den femte månaden efter den månad då licensen utfärdades.
De licenser som utfärdats efter en ansökan inlämnad under juli, augusti och fram till och med den 24 september skall dock endast vara giltiga under 30 dagar från och med den dag de utfärdas, och får inte löpa längre än till och med den 30 september.
4. Den bidragssats som är tillämplig och anges i licensen skall vara den som gäller den dag då ansökan inkommer.
Om någon av de kvantiteter stärkelse som anges i licensen bearbetas under det regleringsår för spannmål som följer på det år då ansökan inkom, skall dock det bidrag som skall utbetalas för den stärkelse som bearbetas under det nya regleringsåret justeras med skillnaden mellan det interventionspris som tillämpas under den månad då bidragslicensen utfärdas och det som tillämpas under bearbetningsmånaden, multiplicerad med koefficienten 1,60. Den omräkningskurs som skall användas för att uttrycka bidragsbeloppet i nationell valuta skall vara den som gäller den dag då stärkelsen bearbetas."
3) I artikel 9.2 skall följande stycke läggas till:
"Det primära kravet, enligt artikel 20 i förordning (EEG) nr 2220/85, är att produkten skall användas eller exporteras i enlighet med de respektive bestämmelserna i artikel 10.1 a och 10.1 b i denna förordning. Användningen eller exporten skall ske inom tolv månader efter det att licensens giltighet har löpt ut. En förlängning av detta slutdatum med som mest sex månader får övervägas på grundval av en välgrundad begäran som lagts fram för den behöriga myndigheten."
4) I artikel 10.4 skall följande stycke läggas till:
"De köpare som per kvartal använder en kvantitet på mindre än 1 000 kg av produkterna enligt detta KN-nummer får emellertid undantas från denna bestämmelse."
5) Artikel 12 skall ersättas med följande: "Artikel 12
Inom tre månader från utgången av varje kvartal skall medlemsstaterna underrätta kommissionen om typen, kvantiteterna och ursprunget (majs, vete, potatis, korn, havre eller ris) av den stärkelse för vilken bidrag har utbetalats och om typen och kvantiteterna av de produkter till vilka stärkelsen har använts."
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1549/98 av den 17 juli 1998 om komplettering av bilagan till förordning (EG) nr 1107/96 beträffande registrering av geografiska beteckningar och ursprungsbeteckningar enligt förfarandet i artikel 17 i rådets förordning (EEG) nr 2081/92 (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING,
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska beteckningar och ursprungsbeteckningar för jordbruksprodukter och livsmedel (1), senast ändrad genom kommissionens förordning (EG) nr 1068/97 (2), särskilt artikel 17.2 i denna, och av följande skäl:
För vissa beteckningar som medlemsstaterna har meddelat i enlighet med artikel 17 i förordning (EEG) nr 2018/92 har det begärts kompletterande uppgifter för att säkerställa att dessa beteckningar uppfyller kraven i artiklarna 2 och 4 i nämnda förordning. Efter granskning av dessa kompletterande uppgifter har det visat sig att dessa beteckningar stämmer överens med artiklarna i nämnda förordning. De bör därför registreras och läggas till i bilagan till kommissionens förordning (EG) nr 1107/96 (3), senast ändrad genom förordning (EG) nr 644/98 (4).
Till följd av de tre nya medlemsstaternas anslutning räknas den tidsfrist på sex månader som föreskrivs i artikel 17 i förordning (EEG) nr 2081/92 från deras anslutningsdag. Vissa av de beteckningar som meddelats av medlemsstaterna överensstämmer med artiklarna 2 och 4 i nämna förordning och bör därför registreras.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för geografiska och ursprungsbeteckningar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (EG) nr 1107/96 skall kompletteras med beteckningarna i bilagan till denna förordning.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1900/98 av den 4 september 1998 om ändring av bilaga I till rådets förordning (EEG) nr 2092/91 om ekologisk produktion av jordbruksprodukter och uppgifter därom på jordbruksprodukter och livsmedel
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2092/91 av den 24 juni 1991 om ekologisk produktion av jordbruksprodukter och uppgifter därom på jordbruksprodukter och livsmedel (1), senast ändrad genom kommissionens förordning (EG) nr 1488/97 (2), särskilt artikel 13 första och andra strecksatsen i denna, och
av följande skäl: Bestämmelser om egenskaperna hos substrat till svampproduktion bör införas i bilaga I så att det blir möjligt att tillåta ekologisk svampproduktion i medlemsstaterna enligt samma produktionsvillkor.
De jordbruksrelaterade komponenterna i dessa substrat bör i princip komma från jordbruksföretag där en ekologisk produktionsmetod används.
Vissa komponenter, särskilt halm och gödsel, kan dock för tillfället inte erhållas i tillräckligt stora mängder från ekologisk produktion. Därför bör en lämplig övergångsperiod fastställas så att producenterna kan anpassa sig till de nya kraven.
I artikel 7.2 tredje strecksatsen ges möjligheten att fastställa särskilda krav på märkning av produkter som framställts med hjälp av vissa produkter som anges i bilaga II till förordning (EEG) nr 2092/91. För just denna produktionstyp är det lämpligt att för en övergångsperiod föreskriva en märkning med upplysningar om det icke-ekologiska ursprunget hos komponenterna i substratet.
Det bör dock övervägas ytterligare förbättringar av bestämmelserna i denna förordning. Detta gäller särskilt bestämmelserna om villkoren för användning, inbegripet villkoren för högsta tillåtna procentandel gödsel som inte kommer från jordbruksföretag där en ekologisk produktionsmetod används samt mycelets egenskaper och ursprung. Det förberedande arbetet bör inledas i tillräckligt god tid så att det kan avslutas innan övergångsperioden går ut.
Övergångsperiodens varaktighet kan komma att ses över om situationen på något sätt förändras när det gäller tillgången på halm och gödsel från ekologisk odling.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som avses i artikel 14 i förordning (EEG) nr 2092/91.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till förordning (EEG) nr 2092/91 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
1. Denna förordning träder i kraft den 1 december 1998.
2. Trots vad som sägs i bestämmelserna i punkt 5.1 och 5.2 i bilaga I får medlemsstaterna under en övergångsperiod som löper ut den 1 december 2001 använda
- produkter som anges i punkt 5.1 a i bilagan och som inte kommer från jordbruksföretag där en ekologisk produktionsmetod används, men som uppfyller de krav som anges i del A första till fjärde strecksatsen i bilaga II till förordning (EEG) nr 2092/91, och/eller
- produkter som anges i punkt 5.2 i bilagan och som inte kommer från jordbruksföretag där en ekologisk produktionsmetod används, men som vid behov uppfyller de krav som anges i del A i bilaga II till förordning (EEG) nr 2092/91,
om de produkter som anges i punkt 5.1 a och 5.2 inte kan erhållas från jordbruksföretag där en ekologisk produktionsmetod används och behovet godkänts av kontrollmyndigheten eller kontrollorganet.
I dessa fall skall märkningen och annonseringen innehålla uppgiften "Svamp som odlats på substrat från extensivt jordbruk som är tillåtet i ekologiskt jordbruk under en övergångsperiod". Ordet "ekologiskt" får inte i denna uppgift, för övrigt på etiketten eller i annonseringen vara mer framträdande än något annat ord i uppgiften.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EG, EKSG, EURATOM) nr 2460/98 av den 12 november 1998 om ändring av förordning nr 7/66/Euratom, 122/66/EEG om fastställande av en lista över de orter för vilka transportbidrag kan beviljas, detta bidrags maximala belopp samt reglerna för dess beviljande
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av ett gemensamt råd och en gemensam kommission för Europeiska gemenskaperna,
med beaktande av kommissionens förslag, och
med beaktande av följande: Med beaktande av rådets förordning (EG, EKSG, Euratom) nr 2458/98 av den 12 november 1998 om ändring av förordning (EEG, Euratom, EKSG) nr 259/68 om fastställande av tjänsteföreskrifter för tjänstemännen i Europeiska gemenskaperna och anställningsvillkor för övriga anställda i dessa gemenskaper samt andra förordningar som skall tillämpas på dessa tjänstemän och anställda vad avser fastställande av löner, pensioner och andra ekonomiska ersättningar i euro (1), bör förordningarna nr 7/66/Euratom och nr 122/66/EEG (2) ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I förordningarna nr 7/66/Euratom, nr 122/66/EEG skall "belgiska franc" ersättas med "euro" och beloppen i belgiska franc ersättas med motsvarande belopp i euroenheter till den av rådet fastställda omräkningskursen.
De regler för avrundning av penningbelopp som fastställs i rådets förordning (EG) nr 1103/97 av den 17 juni 1997 om vissa bestämmelser som har samband med införandet av euron (3) skall tillämpas.
Artikel 2
KOMMISSIONENS FÖRORDNING (EG) nr 2521/98 av den 24 november 1998 om ändring av förordning (EG) nr 577/97 om vissa tillämpningsföreskrifter för rådets förordning (EG) nr 2991/94 om regler för bredbara fetter och rådets förordning (EEG) nr 1898/87 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2991/94 av den 5 december 1994 om regler för bredbara fetter (1), särskilt artikel 8 i denna,
med beaktande av rådets förordning (EEG) nr 1898/87 av den 2 juli 1987 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter (2), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 4.2 i denna, och
av följande skäl: I artikel 2.1 i kommissionens förordning (EG) nr 577/97 av den 1 april 1997 om vissa tillämpningsföreskrifter för rådets förordning (EG) nr 2991/94 om regler för bredbara fetter och rådets förordning (EEG) nr 1898/87 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter (3), senast ändrad genom förordning (EG) nr 1298/98 (4), föreskrivs regler för uppgifter om totala fetthalter i bredbara fetter med undantag för de produkter som avses i förordning (EG) nr 2991/94 med en lägsta fetthalt på 80 %. I artikel 2.3 i förordning (EG) nr 577/97 och i bilaga II till den förordningen fastställs en metod för kontroll av att dessa regler iakttas. Den dag då metoden skall börja tillämpas har skjutits fram till den 1 januari 1999 för att användarna skall ha tid att inhämta erfarenheter från användningen av metoden och för att möjliggöra grundliga studier av metodens genomförbarhet med hjälp av de resultat som kommissionen fått ta del av.
Granskningen av de uppgifter som har lämnats har visat att de toleranser som föreskrivs för kontrollen av fetthalten är alltför snäva. Det har visat sig vara befogat att fördubbla toleranserna för genomsnittet av de prov som tagits samt för de enskilda proven. Under dessa omständigheter kan inte kravet på att resultatet av varje prov skall ligga inom de gränser som fastställs i bilagan till förordning (EG) nr 2991/94 bibehållas. Det bör föreskrivas att de genomsnittliga fetthalter som fastställs skall motsvara dessa gränser.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandena från berörda förvaltningskommittéer.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) Punkterna 1.b och c skall ersättas med följande:
"b) Den genomsnittliga fetthalten får inte avvika med mer än en procentenhet från den angivna halten. Fetthalten i de enskilda proven får avvika med endast två procentenheter från den angivna halten.
c) I alla dessa fall skall den genomsnittliga fetthalten ligga inom de gränser som fastställs i bilagan till förordning (EG) nr 2991/94."
b) Punkt 2 skall ersättas med följande:
Artikel 2
RÅDETS FÖRORDNING (EG) nr 2531/98 av den 23 november 1998 om Europeiska centralbankens tillämpning av minimireserver
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av protokoll nr 3 om stadgan för Europeiska centralbankssystemet och Europeiska centralbanken (nedan kallad stadgan), särskilt artikel 19.2 i denna,
med beaktande av Europeiska centralbankens (nedan kallad ECB) rekommendation (1),
med beaktande av Europaparlamentets yttrande (2),
med beaktande av kommissionens yttrande (3)
i enlighet med det förfarande som anges i artikel 106.6 i Fördraget om upprättandet av Europeiska gemenskapen (nedan kallat fördraget) samt i artikel 42 i stadgan, och på de villkor som anges i artikel 43.1 i stadgan och punkt 8 i protokoll nr 11 om vissa bestämmelser angående Förenade konungariket Storbritannien och Nordirland, och av följande skäl:
(1) Artikel 19.2, jämförd med artikel 43.1, i stadgan, punkt 8 i protokollet nr 11 om vissa bestämmelser angående Förenade konungariket Storbritannien och Nordirland och punkt 2 i protokollet nr 12 om vissa bestämmelser angående Danmark, skall inte medföra att en icke deltagande medlemsstat får några rättigheter eller skyldigheter.
(2) Enligt artikel 19.2 i stadgan skall rådet bland annat fastställa basen för minimireserverna och den högsta tillåtna kvoten mellan dessa reserver och basen för dem.
(3) Enligt artikel 19.2 i stadgan skall rådet även fastställa lämpliga sanktioner vid åsidosättande av dessa skyldigheter, och i den här förordningen fastställs specifika sanktioner. I den här förordningen hänvisas det till rådets förordning (EG) nr 2532/98 av den 23 november 1998 om Europeiska centralbankens befogenhet att förelägga sanktioner (4) när det gäller principer och förfaranden samt anges ett förenklat förfarande för sanktioner avseende vissa typer av regelöverträdelser. Om bestämmelserna i rådets förordning (EG) nr 2532/98 skulle gå emot de bestämmelser i den här förordningen som ger ECB befogenhet att förelägga sanktioner skall bestämmelserna i den här förordningen gälla.
(4) Enligt artikel 19.1 i stadgan får ECB-rådet fastställa regler för att beräkna och fastställa de minimireserver som krävs.
(5) För att systemet med åläggande av minimireserver skall kunna vara ett effektivt verktyg för förvaltning av penningmarknaden och monetär styrning måste det ha en sådan struktur att ECB har förmåga och flexibilitet nog att tillämpa krav på reserver mot bakgrund av och med hänsyn tagen till förändringar i fråga om de ekonomiska och finansiella förhållandena i de deltagande medlemsstaterna. I detta avseende måste ECB vara flexibel nog att reagera för ny betalningsteknik, såsom utvecklingen av elektroniska pengar. För att begränsa möjligheterna att kringgå kraven på minimireserver får ECB tillämpa dem på skyldigheter som härrör från poster utanför balansräkningen, särskilt poster som - antingen enskilt eller i kombination med andra poster i eller utanför balansräkningen - är jämförbara med skyldigheter som är upptagna i balansräkningen.
(6) I arbetet med att fastställa detaljerade regler för åläggandet av minimireserver - inbegripet fastställandet av faktiska reservkvoter, av eventuell avkastning på reserverna, av eventuella undantag från kravet på minimireserver och av eventuella ändringar av kraven på en viss grupp eller vissa grupper av institut - måste ECB sträva efter att uppnå de mål för Europeiska centralbankssystemet (nedan kallat ECBS) som anges i artikel 105.1 i fördraget och som avspeglas i artikel 2 i stadgan. Detta innebär bland annat att ECB måste sträva efter att undvika betydande, icke önskvärda effekter i fråga om undanträngning eller disintermediering. Åläggandet av sådana krav på minimireserver kan utgöra en beståndsdel i utformningen och genomförandet av gemenskapens monetära politik, något som anges som en av ECBS:s grundläggande uppgifter i första strecksatsen i artikel 105.2 i fördraget, och som avspeglas i första strecksatsen i artikel 3.1 i stadgan.
(7) De sanktioner som föreskrivs vid åsidosättande av skyldigheterna enligt den här förordningen påverkar inte ECBS:s möjligheter att fastställa lämpliga bestämmelser för genomförande och påföljder i förhållande till sina motparter, inbegripet möjligheten att helt eller delvis utestänga ett institut från penningpolitiska transaktioner vid allvarligt åsidosättande av kraven på minimireserver.
(8) ECBS och ECB har anförtrotts uppgiften att förbereda de penningpolitiska instrumenten så att de kan ha trätt i kraft fullt ut när den tredje etappen av den ekonomiska och monetära unionen inleds (nedan kallad tredje etappen). Ett väsentligt inslag i dessa förberedelser är att innan den tredje etappen inleds ha antagit de ECB-förordningar enligt vilka instituten måste hålla minimireserver från och med den 1 januari 1999. Det är önskvärt att under 1998 underrätta marknadsaktörerna om de detaljerade bestämmelser som ECB kan anse sig behöva anta för att genomföra systemet med minimireserver. Det är därför nödvändigt att från och med dagen för den här förordningens ikraftträdande utrusta ECB med föreskrivande befogenheter.
(9) Bestämmelserna i den här förordningen kan tillämpas i sin helhet på ett verkningsfullt sätt endast om de deltagande medlemsstaterna vidtar nödvändiga åtgärder så att deras myndigheter har befogenhet att fullt ut bistå och samarbeta med ECB vad gäller insamling och kontroll av uppgifter i enlighet med vad som krävs i den här förordningen och i enlighet med artikel 5 i fördraget.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2) nationell centralbank: en deltagande medlemsstats centralbank,
3) institut: varje enhet i en deltagande medlemsstat som ECB enligt villkoren i artikel 19.1 i stadgan kan ålägga att hålla minimireserver,
4) reservkvot: den andel i procent av basen för minimireserverna som ECB får fastställa i enlighet med artikel 19.1 i stadgan,
5) sanktioner: böter, viten, straffränta och räntelös insättning.
Artikel 2
Rätt att undanta institut
ECB kan på icke-diskriminerande grunder undanta institut från kraven på minimireserver enligt kriterier som fastställs av ECB.
Artikel 3
Bas för minimireserver
1. I basen för de minimireserver som ECB enligt artikel 19.1 i stadgan kan ålägga institut att hålla skall, om inte annat följer av bestämmelserna i punkterna 2 och 3, ingå
i) institutets skyldigheter genom mottagande av medel, tillsammans med
ii) institutets skyldigheter som härrör från poster utanför balansräkningen; i basen skall dock inte ingå
iii) skyldigheter som ett institut helt eller delvis har gentemot andra institut enligt villkor som fastställs av ECB, och inte heller
iv) skyldigheter gentemot ECB eller gentemot nationella centralbanker.
2. För skyldigheter i form av omsättningsbara skuldförbindelser kan ECB som alternativ till bestämmelsen i punkt 1 iii ovan föreskriva att ett instituts skyldigheter gentemot ett annat institut helt eller delvis skall undantas från basen för det fordringsägande institutets minimireserver.
3. ECB kan på icke-diskriminerande grunder tillåta att vissa typer av tillgångar undantas från kategorier av skyldigheter som ingår i basen för minimireserverna.
Artikel 4
Reservkvoter
1. Reservkvoterna, som ECB får fastställa enligt artikel 19.1 i stadgan, får inte överstiga 10 % av någon relevant skyldighet som utgör en del av basen för minimireserverna, men kan vara 0 %.
2. Med förbehåll av punkt 1 kan ECB på icke-diskriminerande grunder fastställa skilda reservkvoter för vissa kategorier av skyldigheter som ingår i basen för minimireserverna.
Artikel 5
Föreskrivande befogenheter
När det gäller artiklarna 2, 3 och 4 skall ECB, när så är lämpligt, anta förordningar eller beslut.
Artikel 6
Rätt att inhämta och verifiera uppgifterna
1. ECB skall ha rätt att från institut inhämta de uppgifter som behövs för genomförandet av kravet på minimireserver. Sådana uppgifter skall vara insynsskyddade.
2. ECB skall ha rätt att med avseende på korrekthet och kvalitet kontrollera den information som instituten tillhandahåller för att visa att de uppfyller kraven på minimireserver. ECB skall underrätta instituten om sitt beslut att verifiera eller inhämta uppgifter.
3. Rätten att verifiera uppgifter skall inbegripa rätten att
a) begära att dokument överlämnas,
b) granska institutens räkenskaper och register,
c) ta kopior av eller göra utdrag ur sådana räkenskaper och register, och
d) begära skriftliga eller muntliga förklaringar.
Om ett institut förhindrar inhämtandet och/eller kontrollen av information skall den deltagande medlemsstat i vilken de relevanta lokalerna är belägna ge det bistånd som krävs, däribland säkerställa tillträde till institutets lokaler så att de ovannämnda rättigheterna kan utövas.
4. ECB får delegera verkställandet av de rättigheter som avses i punkterna 1-3 till de nationella centralbankerna. I enlighet med första strecksatsen i artikel 34.1 i stadgan skall ECB ha befogenhet att i en förordning ytterligare precisera villkoren för utövande av kontrollrätten.
Artikel 7
Sanktioner vid åsidosättande av kraven
1. Om ett institut underlåter att hålla alla eller delar av de minimireserver som krävs enligt den här förordningen och de ECB-förordningar eller ECB-beslut som är knutna till denna förordning, får ECB förelägga institutet endera av följande sanktioner:
a) En räntebetalning uppgående till högst fem procentenheter över ECBS:s marginallåneränta eller två gånger ECBS:s marginallåneränta; i båda fallen skall betalningen beräknas på det belopp varmed det berörda institutets reserver understiger kravet på minimireserver.
b) Ett åläggande av det berörda institutet att göra en räntelös insättning i ECB eller de nationella centralbankerna till ett belopp av högst tre gånger det belopp varmed institutets reserver understiger kravet på minimireserver. Insättningens löptid skall inte överstiga den period under vilken institutet underlåter att hålla minimireserverna.
2. När en sanktion föreläggs enligt punkt 1 skall principerna och förfarandena i förordning (EG) nr 2532/98 tillämpas. Artikel 2.1 och 2.3 och artikel 3.1-3.4 i den förordningen skall dock inte vara tillämpliga, och de tidsfrister som avses i artikel 3.6-3.8 skall förkortas till femton dagar.
3. Om ett institut underlåter att fullgöra skyldigheter enligt den här förordningen eller enligt ECB-förordningar eller ECB-beslut som är knutna till denna förordning, utöver de skyldigheter som avses i punkt 1, skall förordning (EG) nr 2532/98 tillämpas när det gäller sanktioner för sådan underlåtenhet och vad gäller gränser och villkor för sådana sanktioner.
Artikel 8
Slutbestämmelser
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
VERKSTÄLLANDE KOMMITTÉNS BESLUT
av den 16 december 1998
om införande av ett enhetligt formulär för inbjudan eller åtagandeförklaring
(SCH/Com-ex (98) 57)
VERKSTÄLLANDE KOMMITTÉN HAR FATTAT DETTA BESLUT
med beaktande av artikel 132 i konventionen om tillämpning av Schengenavtalet,
med beaktande av artikel 9 i samma konvention, och av följande skäl:
Det ligger i alla Schengenstaters intresse att inom ramen för sin gemensamma politik avseende rörligheten för personer fastställa enhetliga regler för utfärdande av viseringar för att undvika eventuella negativa följder när det gäller inresor till territoriet och den inre säkerheten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Enligt kapitel V punkt 1.4 i de gemensamma konsulära anvisningarna "Prövning av övriga för ansökan nödvändiga verifikationer" skall ett enhetligt formulär användas som bevis för att bostad finns.
Detta formulär medger en stor flexibilitet när det gäller användningen och skall anpassas till den rättsliga situationen för varje avtalsslutande part eftersom Schengenstaterna för närvarande använder mycket olika formulär för olika typer av åtaganden.
Dessa skillnader ökar särskilt risken för missbruk och därför skall ett dokument införas med särskilda kännetecken till skydd mot förfalskning.
Följande delar av dokumentet skall således vara enhetliga:
- Utseendet och strukturen.
- Säkerhetsdetaljerna i dessa dokument.
Det enhetliga formuläret skall användas under 1999 i de stater som tillämpar Schengenkonventionen där detta slags bevis föreskrivs i den nationella lagstiftningen.
1. Följande punkt skall läggas till i kapitel V punkt 1.4 i de gemensamma konsulära anvisningarna: "I de fall då det enligt Schengenstaternas nationella lagstiftning föreligger krav på inbjudningar av privatpersoner eller affärsmän, åtagandeförklaringar eller bevis för att bostad finns skall dessa dokument framläggas i form av ett enhetligt formulär(1)."
2. De avtalsslutande parterna i Schengenavtalet skall fylla i det enhetliga formuläret i enlighet med bestämmelserna i den nationella lagstiftningen.
3. Det enhetliga formulär som skall användas av de avtalsslutande parterna i Schengenavtalet för inbjudningar, åtagandeförklaringar och bevis för att bostad finns skall utarbetas centralt enligt anvisningarna i bilaga A (teknisk beskrivning av säkerhetsdetaljerna) och bilagorna A1 och A2 (modellformulär). De obligatoriska enhetliga uppgifterna i det enhetliga formuläret anges i bilaga B.
4. De modelldokument som utarbetats av de avtalsslutande parterna skall bifogas de gemensamma konsulära anvisningarna som bilaga 15.
5. Frankrike skall förse Schengenstaterna med de filmer som behövs för att framställa formulären. Kostnaderna skall delas mellan de avtalsslutande parterna.
6. Dokumentets säkerhetsmässiga utformning skall kontrolleras regelbundet (eventuellt vartannat år). Säkerhetsdetaljerna skall anpassas vartannat år oberoende av de ändringar av allmän karaktär som visar sig nödvändiga om formuläret förfalskas eller om åtgärder för att skydda de tekniska säkerhetsdetaljerna har blivit kända.
7. Dokumentet skall utarbetas på minst tre språk.
8. Detta beslut träder i kraft när de avtalsslutande parterna har meddelat att åtgärderna har genomförts. Berlin den 16 december 1998. C. H. Schapper
KOMMISSIONENS BESLUT av den 25 januari 1999 om förfarandet för bestyrkande av överensstämmelse av byggprodukter enligt artikel 20.2 i rådets direktiv 89/106/EEG beträffande värmeisoleringsprodukter [delgivet med nr K(1999) 115] (Text av betydelse för EES) (1999/91/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 89/106/EEG av den 21 december 1988 om tillnärmning av medlemsstaternas lagar och andra författningar om byggprodukter (1), ändrat genom direktiv 93/68/EEG (2), särskilt artikel 13.4 i detta, och av följande skäl:
Kommissionen skall välja det av de två förfaranden, enligt artikel 13.3 i direktiv 89/106/EEG för bestyrkande av överensstämmelse av en produkt, som är "minst betungande och samtidigt förenligt med kraven på säkerhet". Detta innebär att det är nödvändigt att besluta om huruvida en tillverkningskontroll i fabriken under tillverkarens ansvar är ett nödvändigt och tillräckligt villkor för bestyrkande av överensstämmelse för en bestämd produkt eller produktgrupp, eller om det av orsaker som rör uppfyllandet av de kriterier som avses i artikel 13.4 krävs att ett godkänt certifieringsorgan deltar.
Enligt artikel 13.4 krävs att det förfarande som sålunda bestämts skall anges i uppdragen och i de tekniska specifikationerna. Det är därför önskvärt att definiera de produkter eller produktgrupper som används i uppdragen och i de tekniska specifikationerna.
De två förfaranden som avses i artikel 13.3 beskrivs i detalj i bilaga III till direktiv 89/106/EEG. Det är därför nödvändigt att klart ange de metoder genom vilka de två förfarandena skall genomföras, i enlighet med bilaga III, för varje produkt eller produktgrupp, eftersom bilaga III anger att vissa system i första hand skall användas.
Det förfarande som avses i artikel 13.3 a motsvarar de system som anges i det första alternativet utan fortlöpande övervakning, samt i det andra och det tredje alternativet i punkt 2 ii i bilaga III och det förfarande som avses i artikel 13.3 b motsvarar de system som anges i punkt 2 i i bilaga III, samt i det första alternativet med fortlöpande övervakning i punkt 2 ii i bilaga III.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga byggkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
För de produkter och produktgrupper som anges i bilaga I skall överensstämmelsen bestyrkas genom ett förfarande där tillverkaren ensam ansvarar för ett system för tillverkningskontroll i fabriken som säkerställer att produkten överensstämmer med de tillämpliga tekniska specifikationerna.
Artikel 2
För de produkter som anges i bilaga II skall överensstämmelsen bestyrkas genom ett förfarande där, förutom ett system för tillverkningskontroll i fabriken som genomförs av tillverkaren, även ett godkänt certifieringsorgan tar del i bedömningen och övervakningen av tillverkningskontrollen eller av själva produkten.
Artikel 3
Förfarandet för bestyrkande av överensstämmelse enligt bilaga III skall anges i uppdragen för harmoniserade standarder.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS DIREKTIV 1999/68/EG
av den 28 juni 1999
om ytterligare bestämmelser för de listor över sorter av prydnadsväxter som förs av leverantörer i enlighet med rådets direktiv 98/56/EG
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 98/56/EG av den 20 juli 1998 om saluföring av förökningsmaterial av prydnadsväxter(1), särskilt artikel 9.4 i detta, och av följande skäl:
1. I kommissionens direktiv 93/78/EEG(2) fastställs genomförandebestämmelser för listor över sorter av prydnadsväxter som förs av leverantörer i enlighet med rådets direktiv 91/682/EEG(3).
2. Direktiv 91/682/EEG skall upphöra att gälla från och med den 1 juli 1999 och ersättas med direktiv 98/56/EG.
3. I enlighet med artikel 9.4 i direktiv 98/56/EG får ytterligare genomförandebestämmelser antagas för de listor över sorter av prydnadsväxter som förs av leverantör och som innehåller teknisk beskrivning och benämningar.
4. Ett system för sortbeskrivning finns redan på gemenskapsnivå inom ramen för gemenskapens växtförädlarrätt.
5. Detta system innehåller också uppgifter om upprätthållande av sorter och om skillnader i förhållande till de mest liknande sorterna.
6. Med hänsyn till utvecklingen av gemenskapens lagstiftning om växtförädlarrätt bör det garanteras att sortbeskrivning enligt direktiv 98/56/EG överensstämmer med denna lagstiftning.
7. Direktiv 93/78/EEG bör upphöra att gälla.
8. De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga kommittén för förökningsmaterial av prydnadsväxter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I detta direktiv fastställs ytterligare genomförandebestämmelser för de listor över sorter av prydnadsväxter och förökningsmaterial av prydnadsväxter som förs av leverantörer i enlighet med artikel 9.1 fjärde strecksatsen i direktiv 98/56/EG.
Artikel 2
1. De listor som förs av leverantörer skall innehålla följande:
i) Sortens namn, i tillämpliga fall tillsammans med dess allmänt kända synonymer.
ii) Uppgifter om upprätthållande av sort och om det förökningssystem som tillämpas.
iii) Sortbeskrivning, åtminstone på grundval av de egenskaper och dessas yttringar såsom de beskrivs i enlighet med bestämmelserna för de ansökningar som skall fyllas i för gemenskapens växtförädlarrätt där denna är tillämplig.
iv) Om möjligt, uppgifter om hur sorten skiljer sig från de sorter som mest liknar den.
2. Punkt 1 ii och iv skall inte omfatta någon leverantör vars verksamhet inskränker sig till utsläppande på marknaden av förökningsmaterial av prydnadsväxter.
Artikel 3
Direktiv 93/78/EEG skall upphöra att gälla från och med det datum som avses i artikel 4 i detta direktiv.
Artikel 4
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv den 31 december 1999. De skall genast underrätta kommissionen om detta.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Medlemsstaterna skall besluta om hur en sådan hänvisning skall göras.
3. Medlemsstaterna skall underrätta kommissionen om de viktigaste bestämmelserna i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 5
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 1999/92/EG
av den 16 december 1999
om minimikrav för förbättring av säkerhet och hälsa för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär (femtonde särdirektivet enligt artikel 16.1 i direktiv 89/391/EEG)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 137 i detta,
med beaktande av kommissionens förslag(1), som överlämnats efter samråd med Rådgivande kommittén för arbetarskyddsfrågor och Kommissionen för säkerhet och hälsa för gruvindustrin och andra utvinningsindustrier,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
enligt förfarandet i artikel 251 i fördraget, och mot bakgrund av det gemensamma utkast som godkändes av förlikningskommittén den 21 oktober 1999(3), och
av följande skäl:
1. I artikel 137 i fördraget föreskrivs att rådet genom direktiv får anta minimikrav för att, främst i fråga om arbetsmiljön främja förbättringar för att garantera en högre skyddsnivå för arbetstagares säkerhet och hälsa.
2. Enligt den artikeln skall dessa direktiv undvika sådana administrativa, finansiella och rättsliga ålägganden som motverkar tillkomsten och utvecklingen av små och medelstora företag.
3. Målsättningen att förbättra arbetstagarnas säkerhet, arbetshygieniska förhållanden och hälsa på arbetsplatsen får inte underordnas rent ekonomiska överväganden.
4. En förutsättning för att kunna säkerställa arbetstagarnas säkerhet och hälsa är att minimikraven för förbättring av säkerhet och hälsa för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär iakttas.
5. Detta direktiv är ett särdirektiv i den mening som avses i artikel 16.1 i rådets direktiv 89/391/EEG av den 12 juni 1989 om åtgärder för att främja förbättringar av arbetstagarnas säkerhet och hälsa i arbetet(4). Bestämmelserna i det direktivet, särskilt de som avser information till arbetstagare, samråd och samverkan med arbetstagarna samt arbetstagares utbildning, är således också fullt tillämpliga för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär, utan att det påverkar tillämpningen av strängare eller mer detaljerade bestämmelser i det här direktivet.
6. Detta direktiv bidrar konkret till att förverkliga den inre marknadens sociala dimension.
7. I Europaparlamentets och rådets direktiv 94/9/EG av den 23 mars 1994 om tillnärmning av medlemsstaternas lagstiftning om utrustning och säkerhetssystem avsedda för användning i explosionsfarliga omgivningar(5) fastställs att det på grundval av artikel 137 i fördraget skall utarbetas ett kompletterande direktiv som i synnerhet skall täcka explosionsfara till följd av användning av en viss utrustning eller till följd av typer av och metoder för installation av utrustning.
8. Explosionsskydd är särskilt viktigt för säkerheten. Genom explosioner äventyras arbetstagarnas liv och säkerhet till följd av okontrollerade flammor och tryckvågor, förekomsten av hälsofarliga reaktionsprodukter och förbrukningen av den omgivande luftens syre som arbetstagarna behöver för att kunna andas.
9. För att fastställa en sammanhängande strategi för explosionsskydd krävs att organisatoriska åtgärder kompletterar de tekniska åtgärderna på arbetsplatsen. I direktiv 89/391/EEG krävs att arbetsgivaren skall ha tillgång till en bedömning av riskerna för arbetstagarnas hälsa och säkerhet på arbetsplatsen. I detta direktiv preciseras detta krav genom att det här föreskrivs att arbetsgivaren skall utarbeta ett explosionsskyddsdokument eller ett antal dokument som uppfyller de minimikrav som fastställs i detta direktiv och som skall hållas aktuellt/a. Detta/dessa explosionsskyddsdokument inbegriper fastställande av farorna, en bedömning av riskerna och fastställande av de särskilda åtgärder som skall vidtas för att säkra arbetstagares hälsa och säkerhet, när de är utsatta för fara orsakad av explosiv atmosfär i enlighet med artikel 9 i direktiv 89/391/EEG. Explosionsskyddsdokument kan vara en del av den riskbedömning i fråga om hälsa och säkerhet i arbetet som krävs enligt artikel 9 i direktiv 89/391/EEG.
10. En bedömning av explosionsrisker kan krävas enligt annan gemenskapslagstiftning. För att undvika onödigt dubbelarbete bör arbetsgivaren, i enlighet med nationell praxis, ha möjlighet att slå ihop dokument, delar av dokument eller liknande rapporter som skall utarbetas i enlighet med annan lagstiftning till en enda säkerhetsrapport.
11. Förebyggande av att explosiva atmosfärer uppstår inbegriper även tillämpning av substitutionsprincipen.
12. Samordning bör ske när arbetstagare från flera företag befinner sig på samma arbetsplats.
13. Förebyggande åtgärder måste vid behov kompletteras med andra åtgärder som genomförs när antändning har skett. Högsta möjliga skyddsnivå uppnås genom att förena förebyggande åtgärder med andra åtgärder som begränsar de skadliga effekterna för arbetstagarna av en explosion.
14. Rådets direktiv 92/58/EEG av den 24 juni 1992 om minimikrav beträffande varselmärkning och signaler för hälsa och säkerhet i arbetet (nionde särdirektivet enligt artikel 16.1 i direktiv 89/391/EEG)(6) är fullt tillämpligt, i synnerhet beträffande områden som omedelbart gränsar till explosionsfarliga områden, där rökning, användning av vinkelslip, svetsning och andra verksamheter som medför lågor eller gnistor kan integreras med explosionsfarliga områden.
15. I direktiv 94/9/EG, delas den utrustning och de säkerhetssystem som omfattas in i utrustningsgrupper och -kategorier. I detta direktiv föreskrivs att arbetsgivaren klassificerar områden där explosiv atmosfär kan uppstå i zoner och beslutar vilka grupper och kategorier av utrustning och säkerhetssystem, som skall användas i varje zon.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
AVDELNING I
ALLMÄNNA BESTÄMMELSER
Artikel 1
Syfte och räckvidd
1. I detta direktiv, som är det femtonde särdirektivet i den mening som avses i artikel 16.1 i direktiv 89/391/EEG, fastställs minimikrav för säkerhet och hälsa för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär enligt definitionen i artikel 2.
2. Direktivet skall inte tillämpas på
a) lokaler som används direkt för och under medicinsk behandling av patienter.
b) användning av anordningar för förbränning av gasformiga bränslen enligt direktiv 90/396/EEG(7).
c) framställning, hantering, användning, förvaring och transport av explosiva substanser eller instabila kemiska substanser.
d) utvinningsindustrin som omfattas av direktiv 92/91/EEG(8) eller 92/104/EEG(9).
e) användning av land-, sjö- och lufttransportmedel på vilka tillämpliga bestämmelser i internationella avtal (till exempel ADNR, ADR, ICAO, IMO, RID) och de gemenskapsdirektiv som ger verkan åt dessa avtal tillämpas. Transportmedel som är avsedda att användas i potentiellt explosiv atmosfär skall inte vara undantagna.
3. Bestämmelserna i direktiv 89/391/EEG och de tillämpliga särdirektiven skall tillämpas fullt ut på det område som avses i punkt 1, utan att det påverkar tillämpningen av strängare och/eller mer specifika bestämmelser i det här direktivet.
Artikel 2
Definition
I det här direktivet avses med explosiv atmosfär en blandning under atmosfäriska förhållanden av luft och brännbara ämnen i form av gas, ånga, dimma eller damm, i vilken förbränningen efter antändning sprider sig till hela den oförbrända blandningen.
AVDELNING II
ARBETSGIVARENS SKYLDIGHETER
Artikel 3
Förebyggande av och skydd mot explosioner
I syfte att i enlighet med artikel 6.2 i direktiv 89/391/EEG förhindra och skydda mot explosioner skall arbetsgivaren med hänsyn till verksamhetens art vidta de tekniska och/eller organisatoriska åtgärder som är lämpliga, i prioriterad ordning, och i enlighet med de grundläggande principerna nedan, för att
- förhindra att explosiv atmosfär bildas, eller, där verksamhetens art inte medger detta,
- undvika att explosiv atmosfär antänds, och
- begränsa de skadliga effekterna av en explosion, för att säkerställa arbetstagarnas hälsa och säkerhet.
Dessa åtgärder skall vid behov kombineras och/eller kompletteras med åtgärder som förhindrar spridning av explosioner och de skall ses över regelbundet och, i alla händelser, när betydande ändringar genomförs.
Artikel 4
Bedömning av explosionsrisker
1. När arbetsgivaren utför de skyldigheter som fastställs i artiklarna 6.3 och 9.1 i direktiv 89/391/EEG skall denne bedöma de särskilda risker som uppstår genom explosiv atmosfär och åtminstone ta hänsyn till
- sannolikheten för att explosiv atmosfär uppstår, samt dess varaktighet,
- sannolikheten för att tändkällor, inklusive elektrostatiska laddningar, förekommer och att dessa aktiveras och får effekt,
- installationerna, ämnen som används, processerna och möjlig växelverkan mellan dessa,
- de förväntade verkningarnas omfattning.
Explosionsriskerna skall bedömas som en helhet.
2. Områden som genom öppningar har eller kan få förbindelse med områden där explosiv atmosfär kan uppstå skall beaktas vid bedömningen av explosionsrisker.
Artikel 5
Allmänna skyldigheter
För att säkerställa arbetstagarnas säkerhet och hälsa och i enlighet med de grundläggande principerna för riskbedömning och de principer som anges i artikel 3 skall arbetsgivaren vidta de åtgärder som är nödvändiga så att
- arbetsmiljön där explosiv atmosfär kan uppstå i sådana mängder att arbetstagares eller andras säkerhet och hälsa äventyras, arbetsmiljön är sådan att arbete kan utföras på ett säkert sätt,
- lämplig övervakning under arbetstagares närvaro säkerställs i enlighet med riskbedömningen genom användning av lämpliga tekniska medel i en arbetsmiljö där explosiv atmosfär kan uppstå i sådana mängder att arbetstagares säkerhet och hälsa äventyras.
Artikel 6
Samordningsskyldighet
Om arbetstagare från flera företag befinner sig på samma arbetsplats skall varje arbetsgivare ansvara för alla frågor som ligger under hans kontroll.
Utan att det åsidosätter det enskilda ansvar som varje arbetsgivare har i enlighet med direktiv 89/391/EEG skall den arbetsgivare som i enlighet med nationell lagstiftning och/eller praxis har ansvaret för arbetsplatsen samordna genomförandet av alla åtgärder om arbetstagarnas hälsa och säkerhet samt i sitt explosionsskyddsdokument, som avses i artikel 8, ange målsättningen för denna samordning liksom åtgärderna och förfarandena för genomförandet.
Artikel 7
Områden där explosiv atmosfär kan uppstå
1. Arbetsgivaren skall klassificera områden där explosiv atmosfär kan uppstå i zoner i enlighet med bilaga I.
2. Arbetsgivaren skall säkerställa att de minimikrav som fastställs i bilaga II tillämpas på områden som omfattas av punkt 1 ovan.
3. Områden där explosiv atmosfär kan uppstå i sådana mängder att arbetstagarnas säkerhet och hälsa äventyras skall vid behov märkas med skyltar vid deras ingångar i enlighet med bilaga III.
Artikel 8
Explosionsskyddsdokument
Vid uppfyllandet av de skyldigheter som anges i artikel 4 skall arbetsgivaren säkerställa att ett dokument, nedan kallat explosionsskyddsdokumentet, utarbetas och hålls aktuellt.
Explosionsskyddsdokument skall särskilt innehålla uppgifter om
- att explosionsriskerna har fastställts och bedömts,
- att lämpliga åtgärder kommer att vidtas för att uppnå syftet med det här direktivet,
- de områden som har klassificerats och delats in i zoner i enlighet med bilaga I,
- de områden på vilka minimikraven i bilaga II tillämpas,
- att arbetsplatsen och arbetsutrustning, inbegripet varningsanordningar, utformas, används och underhålls med vederbörlig hänsyn till säkerhet,
- att åtgärder i enlighet med rådets direktiv 89/655/EEG(10) har vidtagits så att arbetsutrustning används på ett säkert sätt.
Explosionsskyddsdokumentet skall ha utarbetats innan arbetet påbörjas och skall ses över när väsentliga ändringar, utvidgningar eller omvandlingar av arbetsplatsen, arbetsutrustningen eller arbetsorganisationen genomförs.
Arbetsgivaren får kombinera befintliga explosionsriskbedömningar, dokument eller andra jämförliga rapporter som upprättas enligt andra gemenskapsrättsakter.
Artikel 9
Särskilda krav för arbetsutrustning och arbetsplatser
1. Arbetsutrustning, som skall användas i områden där explosiv atmosfär kan uppstå och som redan används eller tillhandahålls i företaget eller i verksamheten för första gången före den 30 juni 2003, skall från och med detta datum uppfylla minimikraven i bilaga II del A, om inga andra gemenskapsdirektiv är tillämpliga eller endast delvis är tillämpliga.
2. Arbetsutrustning, som skall användas i områden där explosiv atmosfär kan uppstå och som tillhandahålls på företaget eller i verksamheten för första gången efter den 30 juni 2003 skall uppfylla de minimikrav som fastställs i bilaga II del A och del B.
3. Arbetsplatser med områden där explosiv atmosfär kan uppstå och som tas i bruk för första gången efter den 30 juni 2003 skall uppfylla minimikraven i detta direktiv.
4. Arbetsplatser med områden där explosiv atmosfär kan uppstå som redan tagits i bruk före den 30 juni 2003 skall senast tre år efter den tidpunkten uppfylla minimikraven i detta direktiv.
5. Om arbetsplatser med områden där explosiv atmosfär kan uppstå förändras, utvidgas eller byggs om efter den 30 juni 2003 skall arbetsgivaren vidta de åtgärder som är nödvändiga så att dessa ändringar, utvidgningar eller ombyggnader överensstämmer med de tillämpliga minimikraven i detta direktiv.
AVDELNING III
ÖVRIGA BESTÄMMELSER
Artikel 10
Ändringar i bilagorna
Rent tekniska ändringar i bilagorna som föranleds av
- antagandet av direktiv om teknisk harmonisering och standardisering avseende området explosionsskydd, och/eller
- den tekniska utvecklingen, ändringar i internationella regelverk eller specifikationer samt nya rön om förebyggande av och skydd mot explosioner
skall antas enligt det förfarande som fastställs i artikel 17 i direktiv 89/391/EEG.
Artikel 11
Handbok för god praxis
Kommissionen skall i en handbok för god praxis av icke bindande natur utarbeta praktiska riktlinjer. Handboken skall behandla de ämnen som anges i artiklarna 3, 4, 5, 6, 7 och 8, bilaga I och bilaga II del A.
Kommissionen skall först samråda med Rådgivande kommittén för arbetarskyddsfrågor i enlighet med rådets direktiv 74/325/EEG(11).
Vid tillämpningen av detta direktiv skall medlemsstaterna i möjligast mån beakta ovannämnda handbok när de utarbetar sin nationella politik för skydd av arbetstagares hälsa och säkerhet.
Artikel 12
Information till företag
Medlemsstaterna skall på begäran sträva efter att göra relevant information tillgänglig för arbetsgivare i enlighet med artikel 11, med särskild hänvisning till handboken för god praxis.
Artikel 13
Slutbestämmelser
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 30 juni 2003. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de redan har antagit eller antar inom det område som omfattas av detta direktiv.
3. Medlemsstaterna skall vart femte år till kommissionen inge en rapport om den praktiska tillämpningen av bestämmelserna i detta direktiv och i denna ange synpunkter som framförts av arbetsmarknadens parter. Kommissionen skall underrätta Europaparlamentet, rådet, Ekonomiska och sociala kommittén samt Rådgivande kommittén för arbetarskyddsfrågor därom.
Artikel 14
KOMMISSIONENS DIREKTIV 1999/98/EG
av den 15 december 1999
om anpassning till den tekniska utvecklingen av Europaparlamentets och rådets direktiv 96/79/EG om skydd av förare och passagerare i motorfordon vid frontalkollision
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(1), senast ändrat genom Europaparlamentets och rådets direktiv 98/91/EG(2), särskilt artikel 13.2 i detta,
med beaktande av Europaparlamentets och rådets direktiv 96/79/EG av den 16 december 1996 om skydd av förare och passagerare i motorfordon vid frontalkollision och om ändring av direktiv 70/156/EEG(3), och
av följande skäl:
1. Direktiv 96/79/EG är ett av särdirektiven i det förfarande för typgodkännande på gemenskapens nivå som inrättats genom direktiv 70/156/EEG. Bestämmelserna i direktiv 70/156/EEG om system, komponenter och tekniska enheter i fordonet är följaktligen tillämpliga på det här direktivet.
2. I enlighet med artikel 4.b i direktiv 96/79/EG skall kommissionen se över och vid behov ändra tillägg 7 till bilaga II så att hänsyn tas till den provning som är avsedd för bedömning av Hybrid III-provdockans fotled, inklusive provning av fordonen.
3. De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från den kommitté för anpassning till teknisk utveckling som inrättats i enlighet med direktiv 70/156/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga II till direktiv 96/79/EG skall ändras i enlighet till bilagan till detta direktiv.
Artikel 2
1. Från och med den 1 oktober 2000 får medlemsstaterna inte, av skäl som hänför sig till den provning som är avsedd för bedömning av Hybrid III-provdockans fotled,
- vägra EG-typgodkännande för en ny fordonstyp, eller
- förbjuda registrering, försäljning eller ibruktagande av ett fordon,
om den provning som är avsedd för bedömning av Hybrid III-provdockans fotled uppfyller kraven i direktiv 96/79/EG, i dess lydelse efter ändringar genom det här direktivet.
2. Från och med den 1 april 2001 får medlemsstaterna inte längre bevilja EG-typgodkännande för en fordonstyp i enlighet med artikel 4 i direktiv 70/156/EEG om den inte uppfyller kraven i direktiv 96/79/EG, i dess lydelse efter ändringar genom det här direktivet.
Artikel 3
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 30 september 2000. De skall genast underrätta kommissionen om detta.
När medlemsstaterna antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texten till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
INTERINSTITUTIONELLT AVTAL
av den 25 maj 1999
EUROPAPARLAMENTET, EUROPEISKA UNIONENS RÅD OCH EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR,
med hänvisning till Europaparlamentets resolution av den 7 oktober 1998 om oberoende, roll och ställning för enheten för samordning av bedrägeribekämpning (Uclaf)(1),
med hänvisning till rådets slutsatser av den 15 mars 1999, som antogs efter en fördjupad diskussion med företrädare för Europaparlamentet och kommissionen,
med beaktande av kommissionens beslut 1999/352/EG, EKSG, Euratom av den 28 april 1999 om inrättande av en europeisk byrå för bedrägeribekämpning(2),
och av följande skäl: (1) Europaparlamentets och rådets förordning (EG) nr 1073/1999(3) och rådets förordning (Euratom) nr 1074/1999(4) om utredningar som utförs av Europeiska byrån för bedrägeribekämpning innehåller bestämmelser om att byrån skall inleda och utföra administrativa utredningar inom de institutioner, organ och byråer som inrättats genom EG-fördraget och Euratomfördraget eller på grundval av dessa fördrag.
(2) Ansvaret för Europeiska byrån för bedrägeribekämpning, som inrättats av kommissionen, förutom skyddet av de ekonomiska intressena även omfattar all verksamhet som har samband med skyddet av gemenskapens intressen mot oegentligheten, som kan leda till administrativa eller straffrättsliga påföljder.
(3) Det är viktigt att öka bedrägeribekämpningens omfattning och effektivitet med hjälp av de experter som finns inom området för administrativa utredningar.
(4) Alla institutioner, organ och byråer bör i kraft av sin administrativa självständighet ge byrån i uppdrag att inom dessa utföra administrativa utredningar för att efterforska sådana omständigheter av allvarlig art som har samband med tjänsteutövningen och som skulle kunna utgöra sådana brister när det gäller att uppfylla de skyldigheter som åligger tjänstemän och anställda i gemenskaperna som avses i artiklarna 11, 12 andra och tredje styckena, 13, 14, 16 och 17 första stycket i tjänsteföreskrifterna för tjänstemän och anställningsvillkoren för övriga anställda i Europeiska gemenskaperna (nedan kallade "Tjänsteföreskrifterna"), brister som kan skada dessa gemenskapers intressen och som kan leda till disciplinära åtgärder och, i förekommande fall, straffrättsliga åtgärder, eller ett allvarligt fel i tjänsten enligt artikel 22 i tjänsteföreskrifterna eller en bristande uppfyllelse av motsvarande skyldigheter som åvilar ledamöter, chefer eller medlemmar av personalen vid gemenskapens institutioner, organ eller byråer, som inte omfattas av tjänsteföreskrifterna.
(5) Dessa utredningar skall utföras med iakttagande av tillämpliga bestämmelser i fördragen om upprättandet av Europeiska gemenskaperna, särskilt protokollet om immunitet och privilegier, texter som antagits för deras tillämpning samt tjänsteföreskrifterna.
(6) Dessa utredningar skall utföras på samma villkor inom alla institutioner, organ och byråer inom gemenskapen utan att överlämnandet av denna uppgift till byrån skall påverka institutionernas, organens och byråernas eget ansvar eller på något sätt minska de berörda personernas rättsliga skydd.
(7) De praktiska villkoren bör fastställas för hur institutionernas och organens ledamöter, byråernas chefer och tjänstemännen och de anställda inom dessa skall samarbeta för att de interna utredningarna skall kunna utföras väl, i avvaktan på att tjänsteföreskrifterna ändras,
efter samråd om att införa en gemensam ordning för detta ändamål, och
med uppmaning till övriga institutioner, organ och byråer att ansluta sig till detta avtal,
INGÅTT FÖLJANDE AVTAL:
1. Europaparlamentet, rådet och kommissionen (nedan kallade: institutionerna) beslutar att anta en gemensam ordning för åtgärder som behövs för att underlätta att de utredningar som genomförs av byrån bedrivs på ett korrekt sätt inom institutionerna. Dessa utredningar har som ändamål att
- bekämpa bedrägerier, korruption och all annan olaglig verksamhet som riktar sig mot Europeiska gemenskapernas ekonomiska intressen,
- efterforska sådana omständigheter av allvarlig art som har samband med tjänsteutövningen och som skulle kunna utgöra brister när det gäller att uppfylla de skyldigheter som åligger tjänstemän och anställda i gemenskaperna, brister som skulle kunna leda till disciplinära åtgärder och, i förekommande fall, straffrättsliga åtgärder, eller en bristande uppfyllelse av motsvarande skyldigheter, som åvilar ledamöter, chefer eller medlemmar av personalen, som inte omfattas av tjänsteföreskrifterna.
Dessa utredningar skall genomföras med iakttagande av tillämpliga bestämmelser i fördragen om upprättandet av Europeiska gemenskaperna, särskilt protokollet om immunitet och privilegier, texter som antagits för deras tillämpning samt tjänsteföreskrifterna.
Utredningarna skall också utföras i enlighet med de villkor och närmare bestämmelser som avses i Europeiska gemenskapens och Europeiska atomenergigemenskapens förordningar.
2. Institutionerna åtar sig att inrätta en sådan ordning och att göra den omedelbart tillämplig genom att anta ett internt beslut enligt den modell som bifogas detta avtal och att inte avvika från modellbeslutet annat än om särskilda förhållanden inom den egna institutionen gör detta nödvändigt av tekniska skäl.
3. Institutionerna är eniga om behovet av att till byrån för yttrande överlämna varje begäran om upphävande av immunitet mot rättsliga förfaranden för tjänstemän eller anställda i samband med eventuella fall av bedrägeri, korruption eller all annan olaglig verksamhet. Om en begäran om upphävande av immunitet gäller någon av institutionernas ledamöter skall byrån underrättas.
4. Institutionerna skall till byrån översända de bestämmelser som de har fastställt för att genomföra detta avtal.
Detta avtal får bara ändras efter uttryckligt medgivande från de undertecknande institutionerna.
De andra institutioner, organ och enheter som inrättats genom EG-fördraget och Euratomfördraget eller på grundval av dessa, uppmanas att ansluta sig till detta avtal genom att, var för sig, avge en förklaring som skall lämnas till ordförandena för de institutioner som undertecknat avtalet.
Detta avtal träder i kraft den 1 juni 1999.
RÅDETS FÖRORDNING (EG) nr 150/1999 av den 19 januari 1999 om ändring av förordning (EEG) nr 2262/84 om särskilda bestämmelser för olivolja
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i denna,
med beaktande av kommissionens förslag (1),
med beaktande av Europaparlamentets yttrande (2), och
av följande skäl: Enligt artikel 1.5 i förordning (EEG) nr 2262/84 (3) skall rådet med kvalificerad majoritet, på förslag från kommissionen, före den 1 januari 1999 fastställa formen för finansieringen av organens utgifter från och med regleringsåret 1999/2000.
Det har fattats beslut om en treårig övergångsperiod från och med regleringsåret 1998/1999 med hänvisning till reformen av den gemensamma organisationen av marknaden för olivolja. De arbetsuppgifter som vanligtvis åläggs organen måste genomföras under övergångsperioden och under det första regleringsåret efter denna period. Det är därför lämpligt att föreskriva att gemenskapen delar organens kostnader för denna period för att se till att de fungerar effektivt och kontinuerligt inom ramen för det administrativa självstyre som föreskrivs i förordning (EEG) nr 2262/84.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 1.5 i förordning (EEG) nr 2262/84 skall de två sista styckena ersättas med följande:
"Organens faktiska utgifter skall för en treårsperiod med början på regleringsåret 1999/2000 till 50 % täckas av gemenskapernas allmänna budget.
Kommissionen skall före den 1 oktober år 2001 undersöka om det är nödvändigt att gemenskapen fortsätter att dela organens utgifter och skall vid behov presentera ett förslag för rådet. Rådet skall, enligt förfarandet i artikel 43.2 i fördraget, före den 1 januari år 2002 besluta om eventuell finansiering av de berörda utgifterna".
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 568/1999 av den 16 mars 1999 om ändring av förordning (EG) nr 577/97 om vissa tillämpningsföreskrifter för rådets förordning (EG) nr 2991/94 om regler för bredbara fetter och rådets förordning (EEG) nr 1898/87 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2991/94 av den 5 december 1994 om regler för bredbara fetter (1), särskilt artikel 8 i denna,
med beaktande av rådets förordning (EEG) nr 1898/87 av den 2 juli 1987 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter (2), senast ändrad genom förordning (EG) nr 222/98 (3), särskilt artikel 4.2 i denna, och
Enligt kompletterande uppgifter som lämnats a
KOMMISSIONENS FÖRORDNING (EG) nr 676/1999 av den 26 mars 1999 om ändring för femte gången av förordning (EG) nr 785/95 om tillämpningsföreskrifter för rådets förordning (EG) nr 603/95 om den gemensamma marknaden för torkat foder
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 603/95 av den 21 februari 1995 om den gemensamma marknaden för torkat foder (1), senast ändrad genom förordning (EG) nr 1347/95 (2), särskilt artikel 18 i denna, och
av följande skäl: I artikel 2.2 a första strecksatsen i kommissionens förordning (EG) nr 785/95 av den 6 april 1995 om tillämpningsföreskrifter för rådets förordning (EG) nr 603/95 (3), senast ändrad genom förordning (EG) nr 1794/97 (4), föreskrivs att dehydratisering av färskt foder skall ske med hjälp av torkar som håller en temperatur på minst 93 °C i början av processen.
Enligt omfattande forskning och vetenskapliga studier bevaras näringsvärdet, särskilt betakarotinhalten, i en produkt av hög kvalitet om torkningen av fodret äger rum vid hög temperatur.
Marknadsläget för torkat foder karakteriseras av fallande försäljningspriser och ökad produktion och är sådant att det är nödvändigt att garantera tillgången på en slutprodukt av näringsmässigt hög kvalitet framställd under likartade konkurrensvillkor och att motivera det stödbelopp som beviljas till bearbetningskostnaderna. Detta kan uppnås genom att torkning av foder vid hög temperatur tillämpas allmänt.
På de flesta företag äger bearbetning av foder rum vid hög temperatur. Det är därför lämpligt att föreskriva att de anläggningar som fortfarande håller en temperatur på 93 °C i början av processen inom rimlig tid justeras för att vara anpassade till torkning av foder vid hög temperatur.
För de tekniska justeringar som är nödvändiga i detta syfte krävs en bekräftelse på att den behöriga myndigheten godkänt företaget.
I vissa medlemsstater används för närvarande ett litet antal bandtorkar med en temperatur på minst 110 °C vid torkningsprocessens början. Det rör sig om små installationer med låg kapacitet vars driftstemperatur inte kan höjas utan radikala tekniska justeringar. Därför bör de omfattas av undantag från minimikravet på en torkningstemperatur på 350 °C, samtidigt som det skall stå klart att ingen ny installation av denna typ får godkännas efter det att regleringsåret 1999/2000 inletts.
I artikel 15 b i ovannämnda förordning (EG) nr 785/95 föreskrivs att medlemsstaterna skall meddela kommissionen de arealer och kvantiteter som berörs av kontrakt och leveransdeklarationer. Erfarenheten har visat att denna rapportering är en källa till motsägelsefulla och otillfredsställande uppgifter. Den bör därför avskaffas.
Förvaltningskommittén för torkat foder har inte avgivet något yttrande inom den tid som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 785/95 ändras på följande sätt:
1. I artikel 2.2 a skall den första strecksatsen ersättas med följande:
Artikel 2
1. De tekniska justeringar i torkningsanläggningarna som är nödvändiga enligt bestämmelserna i artikel 1.1 skall göras utan att det påverkar kravet om att underrätta den behöriga myndigheten inom den tidsfrist som anges i artikel 4.1 a sista stycket i förordning (EG) nr 785/95.
2. Medlemsstaterna skall senast den 15 maj 1999 till kommissionen översända en förteckning över de bandtorkar som godkänts före inledningen av regleringsåret 1999/2000 och som därför får omfattas av undantaget i artikel 1.1.
Artikel 3
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 730/1999
av den 7 april 1999
om handelsnormer för morötter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom kommissionens förordning (EG) nr 2520/97(2), särskilt artikel 2.2 i denna, och
av följande skäl: I bilaga I till förordning (EG) nr 2200/96 återfinns morötter bland de produkter för vilka normer skall antas. Kommissionens förordning (EEG) nr 920/89 av den 10 april 1989 om kvalitetsnormer för morötter, citrusfrukt, äpplen och päron(3), senast ändrad genom förordning (EG) nr 2536/98(4), har genomgått ett flertal ändringar som medför att den ur juridisk synpunkt inte längre kan anses tydlig.
Det är följaktligen nödvändigt att omarbeta nämnda förordning och låta bilaga I till förordning nr 920/89 utgå. För att förbättra överskådligheten på världsmarknaden bör därför de normer för morötter beaktas som rekommenderats av den arbetsgrupp för standardisering av lättfördärvliga livsmedel samt för kvalitetsförbättring som inrättats vid Förenta nationernas ekonomiska kommission för Europa (ECE/FN).
Syftet med dessa normer är att avlägsna produkter av otillfredsställande kvalitet från marknaden, att styra produktionen på ett sådant sätt att den uppfyller konsumenternas krav samt att underlätta handelsförbindelserna på grundval av sund konkurrens och därigenom bidra till att förbättra lönsamheten.
Normerna skall tillämpas i samtliga handelsled. Vid transport över långa sträckor, lagring under en viss tid och olika typer av hantering kan det inträffa att produkterna försämras till följd av sin biologiska utveckling eller sin benägenhet att förfaras. Hänsyn bör därför tas till sådan försämring när normerna tillämpas i de handelsled som ligger efter avsändningstillfället. Eftersom produkter i klass "Extra" skall vara mycket noggrant sorterade och förpackade bör för dem avvikelser endast medges i fråga om bristande färskhet och saftspändhet.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för färsk frukt och färska grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Handelsnormerna för morötter som omfattas av KN-nummer 0706 10 00 anges i bilagan.
Dessa normer skall tillämpas i samtliga handelsled och i enlighet med villkoren i förordning (EG) nr 2200/96.
I de handelsled som ligger efter avsändningstillfället får dock produkterna i förhållande till de föreskrivna normerna
- uppvisa en viss bristande färskhet och saftspändhet, och
- uppvisa mindre förändringar till följd av sin utveckling och benägenhet att förfaras, dock inte om de klassificerats som klass "Extra".
Artikel 2
Förordning (EEG) nr 920/89 ändras på följande sätt:
1) I artikel 1 första stycket skall första strecksatsen utgå.
2) Bilaga I skall utgå.
Artikel 3
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1081/1999
av den 26 maj 1999
om öppnande och förvaltning av tullkvoter för import av tjurar, kor och kvigor av vissa alp- och bergraser som inte är slaktboskap, om upphävande av förordning (EG) nr 1012/98 och om ändring av förordning (EG) nr 1143/98
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött(1), senast ändrad genom förordning (EG) nr 1633/98(2), särskilt artikel 12.1 i denna,
med beaktande av rådets förordning (EG) nr 3066/95 av den 22 december 1995 om vissa medgivanden i form av gemenskapstullkvoter för vissa jordbruksprodukter och om autonom anpassning under en övergångsperiod av vissa jordbrukskoncessioner som föreskrivs i Europaavtalen i syfte att beakta det jordbruksavtal som ingåtts inom ramen för de multilaterala handelsförhandlingarna under Uruguayrundan(3), senast ändrad genom förordning (EG) nr 2435/98(4), särskilt artikel 8 i denna,
med beaktande av rådets förordning (EG) nr 1095/96 av den 18 juni 1996 om genomförande av medgivandena i lista CXL som fastställs sedan förhandlingarna enligt GATT artikel XXIV.6 avslutats(5), särskilt artikel 1.1 i denna, och av följande skäl:
(1) Inom ramen för Världshandelsorganisationen (WTO) har gemenskapen åtagit sig att öppna två tullkvoter med en årlig kvantitet på 5000 djur vardera med en tull på 6 % respektive 4 %. Tullkvoterna gäller tjurar, kor och kvigor av brokig Simmentalras och Schwyz- och Fribourgras som inte är slaktboskap samt kor och kvigor av grå, brun, gul och brokig Simmentalras och Pinzgauras som inte är slaktboskap. Dessa kvoter bör öppnas på flerårsbasis för perioder om tolv månader, nedan kallade importår, som inleds den 1 juli, och tilllämpningsföreskrifter bör fastställas.
(2) Garantier bör särskilt ställas för att alla berörda gemenskapsaktörer skall ges lika och fortlöpande tillträde till kvoten och för att de tullar som fatställts för dessa kvoter skall tillämpas fortlöpande på all import av djuren i fråga fram till dess att kvoten är förbrukad.
(3) Erfarenheten visar att begränsningen av importen kan ge upphov till ansökningar om importlicens i spekulativt syfte. För att de planerade åtgärderna skall fungera som avsett bör huvuddelen av de tillgängliga kvantiteterna förbehållas s.k. traditionella importörer av tjurar, kor och kvigor av vissa alp- och bergraser. I vissa fall finns det en risk för att administrativa felaktigheter som begåtts av den nationella behöriga myndigheten begränsar importörernas tillträde till denna del av kovten. Bestämmelser bör fastställas för att korrigera eventuella felaktigheter.
(4) För att inte förorsaka alltför stor stelhet i handelsförbindelserna inom sektorn bör dock ytterligare en kvantitet ställas till förfogande för sådana importörer som kan visa att de bedriver seriös verksamhet och handlar med betydande kvantiteter med tredje land. För detta ändamål och för att säkerställa en effektiv förvaltning är det lämpligt att kräva att de berörda aktörerna skall ha importerat minst 15 djur under de tolv månader som föregår importåret i fråga. Ett parti på 15 djur utgör i princip en normal last och erfarenheten har visat att försäljning eller inköp av ett enstaka parti utgör ett minimikrav för att en transaktion skall kunna betraktas som reell och ekonomiskt lönsam.
(5) För kontrollen av dessa kriterier krävs att ansökningen lämnas in i den medlemsstat där importören är registrerad i ett register för mervärdesskatt.
(6) För att undvika spekulationer bör s.k. traditionella importörer som inte längre var verksamma inom nötköttssektorn den 1 juni före importåret i fråga inte vara berättigade till kvoten.
(7) Det bör föreskrivas att importtillstånden skall fördelas efter en viss betänketid och eventuellt med tillämpning av en enhetlig procentsats för nedsättning.
(8) Det bör föreskrivas att systemet skall administreras med hjälp av importlicenser. I detta syfte bör närmare bestämmelser fastställas, i synnerhet om inlämnande av ansökningar och om de uppgifter som skall lämnas i ansökningarna och i licenserna, i förekommande fall som undantag från eller tillägg till vissa bestämmelser i kommissionens förordning (EEG) nr 3719/88 av den 16 november 1988 om gemensamma tillämpningsföreskrifter för systemet med import- och exportlicenser samt förutfastställelselicenser för jordbruksprodukter(6), senast ändrad genom förordning (EG) nr 168/1999(7), och i kommissionens förordning (EG) nr 1445/95 av den 26 juni 1995 om tillämpningsföreskrifter för systemet med import- och exportlicenser för nötköttssektorn och om uphävande av förordning (EEG) nr 2377/80(8), senast ändrad genom förordning (EG) nr 2648/98(9).
(9) I artikel 82 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(10), senast ändrad genom förordning (EG) nr 955/1999(11), fastställs att varor som övergår till fri omsättning till en nedsatt tullsats med hänvisning till deras särskilda slutanvändning skall stå under tullens övervakning. En kontroll skall utföras för att säkerställa att de importerade djuren inte slaktas under en viss period. En säkerhet bör ställas för att garantera att dessa djur inte slaktas, vilken skall täcka skillnaden mellan tullarna enligt den gemensamma tulltaxan (GTT) och de nedsatta tullar som gäller den dag då djuren i fråga övergår till fri omsättning.
(10) Kommissionens förordning (EG) nr 1012/98 av den 14 maj 1998 om öppnande och förvaltning av tullkvoter för import av tjurar, kor och kvigor av vissa alp- och bergraser som inte är slaktboskap(12), senast ändrad genom förordning (EG) nr 1143/98(13), bör upphävas.
(11) I artikel 7.2 och 7.3 i kommissionens förordning (EG) nr 1143/98 av den 2 juni 1998 om fastställande av tillämpningsföreskrifter för en tullkvot för kor och kvigor av vissa bergraser som inte är slaktboskap med ursprung i vissa tredje länder och om ändring av förordning (EG) nr 1012/98 föreskrivs, för att garantera efterlevnaden av bestämmelsen om att slakt av de importerade djuren inte är tillåten under en viss period, identifiering av de importerade djuren i enlighet med bestämmelserna i rådets förordning (EG) nr 820/97 av den 21 april 1997 om upprättande av ett system för identifiering och registrering av nötkreatur och om märkning av nötkött och nötköttsprodukter(14) liksom vissa ytterligare relevanta uppgifter. Eftersom dessa uppgifter redan är obligatoriska bör ovan nämnda två punkter utgå.
(12) För tydlighetens skull bör bestämmelserna i artiklarna 2.1 a och 8 c i förordning (EG) nr 1143/98 rättas till.
(13) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för nötkött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. För en flerårsperiod skall under perioden 1 juli-30 juni följande år, nedan kallad importåret, följande tullkvoter öppnas:
>Plats för tabell>
2. Vid tillämpningen av denna förordning skall de djur som avses i punkt 1 inte anses vara slaktdjur om de inte slaktas inom fyra månader från det att deklarationen om övergång till fri omsättning har godkänts.
Undantag kan emellertid beviljas i vederbörligen styrkta fall av force majeure.
3. Tilldelning ur tullkvoten med löpnummer 09.0003 skall beviljas på villkor att följande dokument uppvisas:
- För tjurar: Stamtavla.
- För kor och kvigor: En stamtavla eller ett intyg om registrering i stamboken som styrker rasrenheten.
Artikel 2
1. De två kvoter som avses i artikel 1.1 skall delas i två delar om 80 %, dvs. 4000 djur, respektive 20 %, dvs. 1000 djur.
a) Den första delen av varje kvot om 80 % skall fördelas mellan importörer från gemenskapen som kan styrka att de har importerat djur som omfattas av kvoter med löpnummer 09.0001 och/eller 09.0003 under de 36 månader som föregåJar importåret i fråga.
Medlemsstaterna får som referenskvantiteter emellertid godkänna importtillstånd som hänför sig till föregående importår men som inte har delats ut om detta beror på ett administrativt fel som begåtts av den nationella behöriga myndigheten.
b) Den andra delen av kvoten om 20 % förbehålls sökande som kan styrka att de under de tolv månader som föregick importåret i fråga har importerat minst 15 levande nötkreatur som omfattas av KN-nummer 0102 från tredje land.
Importörerna skall vara registrerade i ett nationellt register för mervärdesskatt.
2. På grundval av ansökningarna om importtillstånd skall fördelningen av den första delen mellan de olika importörerna ske i proportion till storleken på deras import av djur enligt punkt 1 a första stycket under de 36 månader som har föregått importåret i fråga.
3. På grundval av ansökningarna om importtillstånd skall fördelningen av den andra delen ske i proportion till de kvantiteter som de importörer som nämns i punkt 1 b har ansökt om.
Ansökan om importtillstånd
- skall avse minst 15 djur, och
- får inte avse mer än 50 djur.
Ansökningar om importtillstånd för mer än 50 djur skall automatiskt sänkas till detta antal.
4. Import får uteslutande bevisas med hjälp av tulldokumentet om övergång till fri omsättning som vederbörligen attesterats av tullmyndigheterna.
Medlemsstaterna får godta kopior av dessa dokument, som vederbörligen bestyrkts av den utfärdande myndigheten, om den sökande till den behöriga myndighetens tillfredsställelse kan visa att det varit omöjligt för honom att skaffa fram originaldokumentet.
Artikel 3
1. De aktörer som den 1 juni före importåret i fråga inte längre utövade någon verksamhet inom nötköttssektorn skall inte beaktas vid fördelningen i enlighet med artikel 2.1 a första stycket.
2. Ett företag som uppstått genom en sammanslagning av företag som vart och ett enligt artikel 2.2 var berättigat att delta, skall ha samma rättigheter som de ursprungliga företaget.
Artikel 4
1. Ansökan om importtillstånd får endast lämnas in i den medlemsstat där den sökande är registrerad i ett nationellt register för mervärdesskatt.
2. Endast en ansökan per kvot får lämnas in av en och samme aktör och den får avse endast en av delarna av en enskild tullkvot.
Om en sökande lämnar in mer än en ansökan för en enskild kvot, skall inga ansökningar från denne sökande för den aktuella kvoten godtas.
3. Vid tillämpningen av artikel 2.1 a och b skall importörer senast den 15 juni före importåret i fråga för varje löpnummer lämna in ansökningar om importtillstånd till de behöriga myndigheterna, tillsammans med det bevis som anges i artikel 2.4.
4. Efter kontroll av dokumenten skall medlemsstaterna senast den tionde arbetsdagen efter det att perioden för inlämnande av ansökningar löpt ut för varje löpnummer anmäla följande till kommissionen:
- När det gäller den ordning som avses i artikel 2.1 a första stycket, en förteckning över de importörer som uppfyller villkoren för godkännande, med uppgift om deras namn och adress samt antalet importerade djur under den period som avses i artikel 2.2.
- När det gäller den ordning som avses i artikel 2.1 b, en förteckning över de sökande, med uppgift om deras namn och adress samt de kvantiteter som de har ansökt om.
5. Samtliga sådana anmälningar, även anmälningar om att inga ansökningar tagits emot, skall göras via telefax, och utformas enligt förlagorna i bilagorna II och III i de fall då ansökningar har lämnats in.
Artikel 5
1. Kommissionen skall besluta om i vilken utsträckning ansökningar får godkännas.
2. Om de kvantiteter för vilka ansökningar enligt artikel 4.4 andra strecksatsen har lämnats in överstiger de disponibla kvantiteterna, skall kommissionen minska kvantiteterna i ansökningarna med en enhetlig procentsats.
Om den minskning som avses i första stycket resulterar i en kvantitet på mindre än 15 djur per ansökan, skall partier på 15 djur fördelas genom lottdragning av de berörda medlemsstaterna. Om den återstående kvantiteten uppgår till mindre än 15 djur, skall den kvantiteten utgöra ett enda parti.
Artikel 6
1. För att de tilldelade kvantiteterna skall få importeras, krävs det att en eller flera importlicenser uppvisas.
2. Ansökan om importlicens får endast lämnas in till den behöriga myndigheten i den medlemsstat där den sökande har ansökt om importtillstånd.
3. När kommissionen har meddelat fördelningen enligt artikel 5.1, skall importlicenserna utfärdas på begäran av den importör som erhållit importtillståndet och i dennes namn.
4. Licenserna skall vara giltiga i 90 dagar från och med utfärdandedagen enligt artikel 21.1 i förordning (EEG) nr 3719/88. Licenserna får dock endast utfärdas från och med den 1 juli varje importår och skall upphöra att gälla senast den 30 juni.
5. De utfärdade licenserna skall vara giltiga i hela gemenskapen.
6. Utan att det påverkar tillämpningen av bestämmelserna i den här förordningen skall bestämmelserna i förordningarna (EEG) nr 3719/88 och (EG) nr 1445/95 tillämpas.
7. Genom undantag från artikel 9.1 i förordning (EEG) nr 3719/88 får importlicenser, som utfärdats i enlighet med denna förordning, inte överlåtas och de kan endast ge tillgång till tullkvoter om de är utfärdade i samma namn som de deklarationer om övergång till fri omsättning som åtföljer dem.
8. Artikel 8.4 i förordning (EEG) nr 3719/88 skall inte tillämpas.
Artikel 7
1. Kontrollen av att de importerade djuren inte slaktas under en period på fyra månader från dagen för övergång till fri omsättning skall ske i överensstämmelse med bestämmelserna i artikel 82 i förordning (EEG) nr 2913/92.
2. För att garantera att skyldigheten enligt punkt 1 att inte slakta djuren efterlevs, och för att säkerställa uppbörden av obetalda tullar om denna skyldighet inte fullgörs, skall en säkerhet ställas hos de behöriga myndigheterna. Denna säkerhet skall motsvara skillnaden mellan de tullar som fastställts i den gemensamma tulltaxan och de tullar som avses i artikel 1.1 och som är tillämpliga den dag då djuren i fråga övergår till fri omsättning.
Säkerheten skall frisläppas omedelbart om bevis har lagts fram för de berörda tullmyndigheterna att djuren
a) inte har slaktats före utgången av perioden på fyra månader från dagen för deras övergång till fri omsättning,
Artikel 8
Licensansökan och licensen skall innehålla följande:
a) I fält 8, uppgift om ursprungslandet. Licensen innebär skyldighet att importera från det angivna landet.
b) I fält 16, de KN-nummer som anges i bilaga I.
c) I fält 20, en av följande uppgifter:
- Bergrassen (Verordening (EG) nr. 1081/1999), invoerjaar: ...
Artikel 9
1. De kvantiteter som inte omfattas av en ansökan om importlicens per den 15 mars under importåret skall omfattas av en sista fördelning för samma importår som förbehålls de berörda importörer som har ansökt om importlicens för alla de kvantiteter de har rätt till, utan att hänsyn tas till bestämmelserna i artikel 2.1 a och b.
2. I detta syfte skall medlemsstaterna senast den 22 mars under importåret för varje löpnummer till kommissionen anmäla de kvantiteter för vilka det inte har ansökts om importlicens.
3. Kommissionen skall snarast möjligt besluta om dessa återstående kvantiteter.
4. En ansökan om importtillstånd från en importör som avses i punkt 1 skall gälla en kvantitet på 15 djur.
Oavsett om en ansökan avser en kvantitet som överstiger denna kvantitet, skall endast den kvantiteten beaktas.
5. Endast en ansökan per kvot får lämnas in av en och samme aktör.
Om en sökande lämnar in mer än en ansökan för en enskild kvot skall inga ansökningar från denne för den berörda kvoten godtas.
6. Samtliga ansökningar om importtillstånd skall vara de behöriga myndigheterna till handa senast fem arbetsdagar efter dagen för ikraftträdandet för det kommissionsbeslut som avses i punkt 3.
7. För varje löpnummer skall medlemsstaterna senast den sjunde dagen efter det att den period för inlämnande av ansökningar som anges i punkt 6 gått till ända till kommissionen överlämna en förteckning över de sökande och vilka kvantiteter de har ansökt om.
8. Vid tillämpningen av denna artikel skall bestämmelserna i artiklarna 5-8 gälla i tillämpliga delar.
Artikel 10
förordning (EG) nr 1012/98 upphör att gälla.
Artikel 11
Förordning (EG) nr 1143/98 ändras på följande sätt:
1) Artikel 2.1 a andra stycket skall ersättas med följande: "Medlemsstaterna får emellertid som referenskvantiteter godkänna importtillstånd som hänför sig till föregående importår men som inte har delats ut om detta beror på ett administrativt fel som begåtts av den nationella behöriga myndigheten."
2) I artikel 7 skall punkterna 2 och 3 utgå.
3) Artikel 8 c skall ersättas med följande: "c) I fält 20, en av följande uppgifter:
- Bjergracer (forordning (EF) nr. 1143/98), importår: ...
- Bergraser (förordning (EG) nr 1143/98), importår: ..."
Artikel 12
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1125/1999
av den 28 maj 1999
om ändring av kommissionens förordning (EG) nr 111/1999 om tillämpningsföreskrifter för rådets förordning (EG) nr 2802/98 om ett program för leverans av jordbruksprodukter till Ryska federationen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2802/98 av den 17 december 1998 om ett program för leverans av jordbruksprodukter till Ryska federationen(1), särskilt artikel 4.2 i denna, och av följande skäl:
(1) I kommissionens förordning (EG) nr 111/1999(2) fastställs allmänna tillämpningsföreskrifter för genomförande av leveranser enligt den ordning som fastställs i förordning (EG) nr 2802/98.
(2) Mot bakgrund av de tekniska arrangemang som överenskommits mellan de ryska myndigheterna och kommissionen, efter det att förordningen trädde i kraft, bör de allmänna tillämpningsföreskrifterna ändras på ett antal punkter, särskilt när det gäller bestämmelserna för hur mottagarlandet övertar produkterna och kommissionens förfarande för kontroll av hur leveranserna genomförs.
(3) Beträffande bearbetade produkter på basis av produkter från interventionslager eller på basis av produkter som anskaffats på gemenskapsmarknaden bör bestämmelserna om intyg om överensstämmelse ändras, särskilt när det gäller hur kontrollerna organiseras, och det bör fastställas mer detaljerade bestämmelser för hur den aktör som innehar kontraktet för transport av varorna utanför gemenskapen skall överta produkterna.
(4) För att göra det enklare för aktörer att delta i anbudsförfarandena förefaller det lämpligt att lätta på vissa av de ursprungliga kraven i anbudsinfordran och att ange mer detaljerade bestämmelser för hur leveranserna skall genomföras.
(5) Det är lämpligt att föreskriva omedelbar tillämpning av de ändringar som följer av de tekniska arrangemang som överenskommits med de ryska myndigheterna beträffande bestämmelserna för produktövertag och beträffande vissa bestämmelser för kontroll i samband med produktuttag och för frisläppande av säkerheter till förmån för aktörerna.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandena från samtliga berörda förvaltningskommittéer.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 111/1999 ändras på följande sätt:
5) I artikel 5.1 f skall punkt 4 utgå.
8) I artikel 5.1 g skall punkt 4 utgå.
9) I artikel 5.1 i skall "i enlighet med den förlaga som återfinns i bilaga III" ersättas med "i enlighet med den förlaga som återfinns i bilaga IV".
14) Artikel 6.5 skall utgå.
Varorna kan lastas så snart interventionsorganet erhållit bevis för att det har ställts en leveranssäkerhet i enlighet med punkt 4."
1. För de leveranser som avser produktion av helt slipat ris eller anskaffande av griskött på gemenskapsmarknaden skall kontraktsinnehavaren erhålla ett fast belopp på 0,45 euro per ton (netto) och dag för ris och på 0,90 euro per ton (netto) och dag för griskött för att täcka alla omkostnader (parkering, försäkring, bevakning, säkerhet, osv.) som uppstår i de fall då transportören utan egen förskyllan inte kan agera inom de föreskrivna tidsramarna.
2. Vid leverans enligt artikel 2.1 a skall interventionsorganet utfärda uttagsintyget senast tre arbetsdagar efter det att samtliga varor i ett av de magasin som anges i respektive förordning om leverans tagits ut. Interventionsorganet skall stå för de omkostnader som uppstår på grund av att uttagsintyget utfärdas för sent och dessa omkostnader skall beräknas genom tillämpning av en räntesats som skall vara samma som den räntesats som anges i bilaga VII och som är tillämplig i den berörda medlemsstaten den sista dagen för inlämning av anbud, höjd med 1 1/2 punkt."
17) I artikel 9.1 skall andra stycket ersättas med följande: "För de leveranser som avser produktion av helt slipat ris eller anskaffande av griskött på gemenskapsmarknaden skall det uttagsintyg som utfärdas i enlighet med bilaga V och som undertecknas av det organ som ansvarar för utfärdandet av detsamma utgöra bevis för att produkten uppfyller de krav som fastställts för leveransen."
1. Begäran om betalning för leveransen skall inlämnas till det interventionsorgan som avses i artikel 4 inom två månader från utgången av den leveransperiod som fastställs i anbudsinfordran. Om denna bestämmelse inte iakttas, med undantag för fall av force majeure, skall beloppet minskas med 10 % för den första månadens försening. Vid ytterligare försening skall beloppet minskas med 5 % per månad.
2. Begäran om betalning för leveransen skall
a) i de fall då artikel 2.1 b tillämpas, åtföljas av
- en kopia av transportdokumenten,
- övertagandeintyg i original, i enlighet med bilaga I, utfärdat av det kontrollorgan som utsetts av kommissionen och undertecknat av den företrädare för mottagarlandet som anges i bilagan till förordningen om anbudsförfarande,
- intyg om överensstämmelse vid bestämmelseorten i enlighet med artikel 9.7,
- en kopia av exportlicensen eller exportdeklarationen, i de fall då det enligt lagstiftningen beträffande den gemensamma organisationen av marknaden inte krävs någon exportlicens,
b) i de fall då artikel 2.1 a tillämpas och utöver de intyg som anges ovan i a, åtföljas av det kontrolldokument som anges i artikel 14.2.
3. Vid leverans enligt artikel 2.1 a eller b skall leveranskostnaderna betalas för den kvantitet som anges i övertagandeintyget som skall utfärdas av det kontrollorgan som kommissionen utser och som skall viseras av de företrädare för mottagarlandet som anges i förordningen om öppnande av ett anbudsförfarande. Övertagandeintyget skall utfärdas i enlighet med bilaga I.
4. Vid anbudsförfarande enligt artikel 2.2 skall den kvantitet interventionsprodukter för vilken anbudsgivaren tilldelats kontrakt ställas till dennes förfogande när det har styrkts att det ställts säkerhet i enlighet med artikel 7.2.
5. Vid leverans enligt artikel 2.3 skall betalningen till den anbudsgivare som tilldelats kontrakt för anskaffande av produkter ske mot uppvisande av det uttagsintyg i enlighet med bilaga V som skall utfärdas av transportören och som skall viseras av kontrollorganet enligt artikel 9.1 efter det att hela partiet lastats.
6. Om övertagandet på bestämmelseorten fördröjs på grund av omständigheter som inte kan påverkas av kontraktsinnehavaren, skall mottagarlandet ersätta anbudsgivaren för dennes extrakostnader på grundval av bestyrkande handlingar.
"3. Om det vid leveransstadiet kan konstateras att förseningar har uppstått skall 0,75 euro per ton av leveranssäkerheten förverkas för varje dags försening av den del av kvantiteten som lastats eller levererats för sent. Om sådana förseningar överstiger elva dagar skall avdraget ökas till 1 euro per ton för varje ytterligare dag. Dessa bestämmelser skall tillämpas när kontraktsinnehavaren är ansvarig för förseningen av lastningen eller leveransen."
24) I artikel 13 skall följande införas som tredje stycket: "Förskottssäkerheten skall frisläppas när villkoren för betalning av leveransen i enlighet med artikel 10 har uppfyllts."
3. I de fall då det för export av en produkt krävs att exportlicensansökan uppvisas skall denna åtföljas av ett bevis för att sökanden är innehavare av ett kontrakt avseende leveranser enligt förordning (EG) nr 2802/98. Beviset skall utgöras av en kopia av det meddelande om tilldelning av leveranskontrakt som avses i artikel 6.3.
Exportlicensen skall utfärdas endast om det bevisas att den leveranssäkerhet som avses i artikel 7 har ställts. Ställandet av denna säkerhet skall anses utgöra ställandet av licenssäkerheten. Trots bestämmelserna i avdelning III avsnitt 4 i förordning (EEG) nr 3719/88 skall säkerheten frisläppas på de villkor som fastställs i artikel 12.2."
26) Bilaga II skall ersättas med bilaga A till den här förordningen.
28) Bilaga B till den här förordningen skall införas som bilaga VII.
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1245/1999
av den 16 juni 1999
om godkännande av nya fodertillsatser
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 70/524/EEG av den 23 november 1970 om fodertillsatser(1), senast ändrat genom kommissionens förordning (EG) nr 866/1999(2), särskilt artiklarna 9j och 3 i detta, och av följande skäl:
(1) Enligt direktiv 70/524/EEG får nya fodertillsatser och nya användningsområden för fodertillsatser tillåtas mot bakgrund av den vetenskapliga och tekniska utvecklingen.
(2) I flera medlemsstater har försök i stor skala gjorts med en ny fodertillsats, "natrolit-fonolit" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel". Med hänsyn till de erfarenheter som har gjorts bör denna nya fodertillsats kunna tillåtas.
(3) I vissa medlemsstater har framgångsrika försök gjorts med en annan ny fodertillsats, "Hydratiserad kalciumaluminiumsilikat av vulkaniskt ursprung" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel". Denna nya fodertillsats bör tillåtas tillfälligt.
(4) Nya fodertillsatser och nya användningsområden för fodertillsatser får tillåtas tillfälligt under förutsättning att de halter som tillåts i foder inte medför fara för miljön eller människors eller djurs hälsa och inte är till skada för konsumenterna genom att djurproduktens egenskaper förändras, att tillsatsens närvaro i foder kan kontrolleras och att närvaron av fodertillsatsen enligt tillgängliga forskningsresultat sannolikt har en gynnsam effekt på foderegenskaperna eller på djuruppfödningen.
(5) Det tillfälliga godkännandet av "natrolit-fonolit" slutade gälla redan den 21 april 1999. Av rättssäkerhetsskäl är det därför nödvändigt att denna förordning tillämpas retroaktivt.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga foderkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
"Natrolit-fonolit" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel" skall tillåtas enligt direktiv 70/524/EEG som fodertillsats E 566 på de villkor som anges i bilaga I till den här förordningen.
Artikel 2
"Hydratiserad kalciumaluminiumsilikat av vulkaniskt ursprung" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel" får tillåtas enligt direktiv 70/524/EEG som fodertillsats nr 3 på de villkor som anges i bilaga II till den här förordningen.
Artikel 3
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
RÅDETS FÖRORDNING (EG) nr 1258/1999
av den 17 maj 1999
om finansiering av den gemensamma jordbrukspolitiken
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3),
med beaktande av revisionsrättens yttrande(4), och
av följande skäl: 1. Genom förordning nr 25 om finansieringen av den gemensamma jordbrukspolitiken(5) upprättade rådet Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ), nedan kallad "fonden", som utgör en del av Europeiska gemenskapernas allmänna budget. I den förordningen fastställs de principer som skall tillämpas för finansieringen av den gemensamma jordbrukspolitiken.
2. Med hänsyn till att den inre marknaden innebär enhetliga prissystem och en gemensam jordbrukspolitik, bör gemenskapen stå för de ekonomiska följderna. I enlighet med denna princip, som fastställs i artikel 2.2 i förordning nr 25, bör fondens garantisektion finansiera bidrag vid export till tredje land, intervention i syfte att stabilisera jordbruksmarknader, åtgärder för landsbygdsutveckling, särskilda veterinäråtgärder enligt rådets beslut 90/424/EEG av den 26 juni 1990 om utgifter inom veterinärområdet(6), åtgärder för att informera om den gemensamma jordbrukspolitiken samt vissa utvärderingar i syfte att uppnå målen i artikel 33.1 i fördraget.
3. Fondens utvecklingssektion bör finansiera utgifter för vissa åtgärder för landsbygdsutveckling i regioner som utvecklas långsammare samt för gemenskapens initiativ för landsbygdsutveckling.
4. Kommissionen ansvarar för förvaltningen av fonden. Ett nära samarbete mellan medlemsstaterna och kommissionen i en kommitté för Europeiska utvecklings- och garantifonden för jordbruket föreskrivs.
5. Ansvaret för kontrollen av garantisektionens utgifter inom fonden ligger i första hand hos medlemsstaterna, som utser myndigheter och andra organ som skall verkställa utgifter. Medlemsstaterna skall fullt ut och på ett effektivt sätt ta på sig denna uppgift. Kommissionen, som är ansvarig för att verkställa gemenskapens budget, måste kontrollera de sätt på vilka dessa utbetalningar och kontroller har utförts. Kommissionen får finansiera utgifter enbart om detta sker på ett sätt som ger tillräckliga garantier för att gemenskapsbestämmelserna efterlevs. Inom ramen för ett decentraliserat system för förvaltning av gemenskapens utgifter är det av avgörande betydelse att kommissionen, som är den institution som är ansvarig för finansieringen, är berättigad till och har möjlighet att utföra alla kontroller som den anser nödvändiga, med avseende på förvaltningen av utgifterna, samt att öppenheten och det ömsesidiga biståndet mellan medlemsstaterna och kommissionen är effektiva och fullständiga.
6. I samband med granskning och godkännande av räkenskaperna kan kommissionen inom skälig tid besluta om de totala utgifter som skall införas i garantisektionen i räkenskaperna, endast om den får tillfredsställande garantier för att de nationella kontrollerna är tillräckliga och ger insyn i verksamheten, och att utbetalningsställena försäkrar sig om att de utbetalningar som de gör är lagliga och riktiga. Bestämmelser bör därför antas för ackreditering av utbetalningsställena från medlemsstaternas sida. För att säkerställa konsekvens i den standard som krävs för ackreditering i medlemsstaterna skall kommissionen dra upp riktlinjer avseende de kriterier som skall tillämpas. Det bör därför föreskrivas att enbart utbetalningar som görs av de utbetalningsställen som är ackrediterade av medlemsstaterna får verkställas. För alt säkerställa insyn i de nationella kontrollsystemen, särskilt såvitt avser förfarandet för godkännande, bemyndigande och utbetalning, bär i förekommande fall antalet myndigheter och organ som anförtros detta ansvar begränsas med hänsyn till varje medlemsstats konstitutionella bestämmelser.
7. Ett decentraliserat förvaltningssystem för gemenskapens fonder innebär, särskilt efter reformen av den gemensamma jordbrukspolitiken, att flera utbetalningsställen kan utses. När en medlemsstat ackrediterar fler än ett utbetalningsställe måste den därför utse ett enda kontaktorgan för att säkerställa konsekvens av fondernas förvaltning, upprätta kontakter mellan kommissionen och de olika ackrediterade utbetalningsställena och säkerställa att sådana uppgifter om olika utbetalningsställens transaktioner som kommissionen begär skall kunna göras tillgängliga med kort varsel.
8. Medlemsstaterna måste tillhandahålla finansiella medel i enlighet med utbetalningsställenas behov, medan kommissionen gör förskottsutbetalningar mot utbetalningsställenas verkställda utgifter. Inom ramen för åtgärder för landsbygdsutveckling bör verkliga förskottsbetalningar göras för genomförande av program. Dessa förskottsbetalningar bör behandlas enligt de finansiella mekanismer som har upprättats för förskott mot de verkställda utgifter som har betalats under en referensperiod.
9. Det är lämpligt att föreskriva två olika slag av beslut, ett som avser granskning och godkännande av räkenskaperna för fondens garantisektion, och ett som lägger fast vilka slutsatser, inbegripet finansiella rättelser, som kan dras av resultaten av granskningen huruvida utgifterna överensstämmer med gemenskapsbestämmelserna.
10. Granskningen av överensstämmelse och därpå följande beslut om ackreditering kommer således inte längre att vara knutna till verkställandet av budgeten för ett visst budgetår. Det är nödvändigt att fastställa den längsta period som slutsatserna av granskningen av överensstämmelse kan avse. Åtgärderna för landsbygdsutveckling är emellertid fleråriga, vilket gör att det inte är möjligt att tillämpa en sådan längsta period.
11. Åtgärder måste vidtas för att förhindra och ingripa mot oegentligheter och för att återkräva belopp som förlorats till följd av sådana oegentligheter eller sådan försumlighet. Det ekonomiska ansvaret för sådana oegentligheter eller sådan försumlighet måste fastställas.
12. Gemenskapens utgifter måste noga övervakas. Utöver den övervakning som medlemsstaterna utför på eget initiativ och som förblir av största vikt, bör bestämmelser fastställas så att kommissionens tjänstemän kan genomföra kontroller och ha rätt att begära hjälp från medlemsstaterna.
13. Det är nödvändigt att i största möjliga utsträckning använda informationsteknik för att få fram den information som skall sändas till kommissionen. När kommissionen utför kontroller måste den ha fullständig och omedelbar tillgång till uppgifter som rör utgifter, både i dokument och i datafiler.
14. Med hänsyn till omfattningen av gemenskapsfinansieringen måste Europaparlamentet och rådet regelbundet informeras genom finansiella rapporter.
15. För att förenkla den finansiella förvaltningen är det önskvärt att närma fondens finansieringsperiod till budgetåret såsom det anges i artikel 272.1 i fördraget. För att detta skall kunna göras måste det finnas en klar bild av vilka medel som finns tillgängliga vid utgången av budgetåret i fråga. Det bör därför föreskrivas att kommissionen får nödvändig befogenhet att anpassa fondens finansieringsperiod om tillräckliga budgetmedel finns tillgängliga.
16. Rådets förordning (EEG) nr 729/70 av den 21 april 1970 om finansiering av den gemensamma jordbrukspolitiken(7) har ändrats i betydande omfattning vid ett flertal tillfällen. Nu när nya ändringar görs av nämnda förordning är det önskvärt att bestämmelserna i fråga omarbetas för att förtydliga vissa frågor.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Den skall bestå av följande två sektioner:
- Garantisektionen.
- Utvecklingssektionen.
2. Garantisektionen skall finansiera
a) bidrag vid export till tredje land,
b) intervention i syfte att stabilisera jordbruksmarknaden,
c) åtgärder för landsbygdsutveckling utanför mål 1-program med undantag av gemenskapsinitiativet för landsbygdsutveckling,
d) gemenskapens finansiella bidrag till särskilda veterinära åtgärder, kontrollåtgärder på veterinärområdet och program för bekämpning och övervakning av djursjukdomar (veterinära åtgärder) samt till växtskyddsåtgärder,
e) åtgärder avsedda att ge information om den gemensamma jordbrukspolitiken och vissa utvärderingar av åtgärder som finansieras av fondens garantisektion.
3. Utveckingssektionen skall finansieras sådana åtgärder för landsbygdsutveckling som inte omfattas av punkt 2 c.
4. Utgifter för administration och personal som belastar medlemsstater och mottagare av stöd från fonden skall inte finansieras av fonden.
Artikel 2
1. Bidrag vid export till tredje land, beviljade i enlighet med gemenskapsbestämmelserna inom ramen för den gemensamma organisationen av jordbruksmarknaderna skall finansieras enligt artikel 1.2 a.
2. Intervention för att stabilisera jordbruksmarknaderna som görs i enlighet med gemenskapsbestämmelser inom ramen för den gemensamma organisationen av jordbruksmarknaderna skall finansieras enligt artikel 1.2 b.
3. Om det är nödvändigt skall rådet, på förslag av kommissionen, med kvalificerad majoritet fastställa föreskrifter för finansiering av de åtgärder som avses i punkterna 1 och 2.
Artikel 3
1. Åtgärder för landsbygdsutveckling utanför mål 1-programmen som vidtas enligt gemenskapsbestämmelser skall finansieras enligt artikel 1.2 c.
2. Veterinära åtgärder och växtskyddsåtgärder som vidtas enligt gemenskapsbestämmelser skall finansieras enligt artikel 1.2 d.
3. Informationsåtgärder och utvärderingsåtgärder som vidtas enligt gemenskapsbestämmelser skall finansieras enligt artikel 1.2 e.
4. Tillämpningsföreskrifter för denna artikel skall antas i enlighet med förfarandet i artikel 13.
Artikel 4
1. Varje medlemsstat skall underrätta kommissionen om följande:
a) De myndigheter och organ som den ackrediterar för att göra de betalningar som avses i artiklarna 2 och 3, nedan kallade "utbetalningsställen".
b) Om fler än ett utbetalningsställe har ackrediterats, den myndighet eller det organ, nedan kallat "samordningsorgan", som den ger i uppdrag dels att samla in och överföra de uppgifter som skall ges in till kommissionen, dels att främja en enhetlig tillämpning av gemenskapsbestämmelserna.
2. Utbetalningsställena skall vara medlemsstaternas myndigheter och organ som, såvitt avser de betalningar som skall göras inom deras områden skall ge tillräckliga garantier för att
a) ansökningarnas berättigande och överensstämmelse med gemenskapsbestämmelserna kontrolleras innan betalningarna godkänns,
b) de gjorda betalningarna redovisas korrekt och fullständigt i räkenskaperna,
c) nödvändiga handlingar ges in inom den tid och i den form som föreskrivs i gemenskapsbestämmelserna.
3. Utbetalningsställena skall inneha verifikationshandlingar avseende de gjorda utbetalningarna och handlingar som gäller genomförandet av de föreskrivna administrativa och fysiska kontrollerna. Om de relevanta handlingarna förvaras hos de organ som har till uppgift att godkänna utgifterna, skall dessa organ tillställa utbetalningsstället rapporter om antalet genomförda kontroller, dessas innehåll och de åtgärder som har vidtagits mot bakgrund av resultaten.
4. Endast utgifter som betalas av ackrediterade utbetalningsställen skall finansieras av gemenskapen.
5. Varje medlemsstat skall, med beaktande av landets konstitutionella bestämmelser och institutionella struktur, begränsa antalet ackrediterade utbetalningsställen till minsta möjliga antal för att de utgifter som avses i artiklarna 2 och 3 skall kunna betalas under tillfredsställande förvaltnings- och redovisningsförhållanden.
6. Varje medlemsstat skall till kommissionen överlämna följande upplysningar om utbetalningsställena:
a) Namn och stadgar.
b) Förvaltnings- och redovisningsförhållanden samt interna kontrollförhållanden under vilka betalningar skall göras i samband med genomförandet av gemenskapsbestämmelserna inom ramen för den gemensamma jordbrukspolitiken.
c) Ackrediteringshandlingen.
Kommissionen skall omedelbart underrättas om dessa uppgifter ändras på något sätt.
7. Om ett eller flera av villkoren för ackrediteringen inte har uppfyllts eller inte längre uppfylls av ett godkänt utbetalningsställe skall ackrediteringen återkallas, såvida inte utbetalningsstället genomför nödvändiga anpassningar inom den tid som bestäms utifrån hur allvarligt problemet är. Den berörda medlemsstaten skall underrätta kommissionen om detta.
8. Tillämpningsföreskrifterna för denna artikel skall antas i enlighet med förfarandet i artikel 13.
Artikel 5
1. De ekonomiska resurser som krävs för att täcka de utgifter som avses i artiklarna 2 och 3 skall göras tillgängliga för medlemsstaterna av kommissionen genom förskott på utgifter som verkställts under en referensperiod.
Förskottsbetalning för genomförande av program inom ramen för de åtgärder för landsbygdsutveckling som avses i artikel 3.1 får beviljas av kommissionen när dessa program godkänns och skall betraktas som utgifter som verkställts den första dagen i månaden efter beslutet om beviljandet.
2. Till dess att förskotten på verkställda utgifter har utbetalats skall medlemsstaterna tillhandahålla de medel som är nödvändiga för att täcka nämnda utgifter, alltefter de godkända utbetalningsställenas behov.
3. Tillämpningsföreskrifterna för denna artikel skall antas i enlighet med förfarandet i artikel 13.
Artikel 6
1. Medlemsstaterna skall med jämna mellanrum tillställa kommissionen följande uppgifter om de ackrediterade utbetalningsställena och samordningsorganen och de transaktioner som finansieras av fondens garantisektion:
a) En redovisning av utgifterna och en bedömning av finansieringsbehoven.
b) Årsredovisningen tillsammans med nödvändiga underlag för granskning och godkännande samt ett intyg avseende den vidarebefordrade redovisningens fullständighet, exakthet och sanningsenlighet.
2. Tillämpningsföreskrifter för denna artikel, särskilt de som gäller det redovisningsintyg som avses i punkt 1 b, skall antas enligt förfarandet i artikel 13.
Artikel 7
1. Efter att ha hört fondkommittén skall kommissionen fatta de beslut som anges i punkterna 2, 3 och 4.
2. Kommissionen skall besluta om månatliga förskott på verkställda utgifter som betalas av de ackrediterade utbetalningsställena.
Utgifterna för oktober skall hänföras till oktober om de verkställs mellan den 1 och den 15 oktober och till november om de verkställs mellan den 16 och den 31 oktober. Förskottsbetalningar skall göras till medlemsstaten senast den tredje arbetsdagen i den andra månaden efter den månad då utgifterna verkställs.
Ytterligare förskott får göras om fondkommittén underrättas vid nästa samråd.
3. Kommissionen skall före den 30 april året efter det aktuella budgetåret på grundval av de uppgifter som avses i artikel 6.1 b granska och godkänna räkenskaperna för utbetalningsställena.
Beslutet att granska och godkänna räkenskaperna skall omfatta den överlämnade redovisningens fullständighet, exakthet och sanningsenlighet. Beslutet skall inte påverkar antagandet av ett senare beslut i enlighet med punkt 4.
4. Kommissionen skall besluta om vilka utgifter som inte skall omfattas av gemenskapsfinansiering enligt artiklarna 2 och 3 om den finner att utgifterna inte har verkställts i överensstämmelse med gemenskapsbestämmelserna.
Före varje beslut om att vägra finansiering skall resultaten av kommissionens kontroller och den berörda medlemsstatens svar överlämnas skriftligen, varefter båda parter skall söka nå en överenskommelse om vilka åtgärder som skall vidtas.
Om ingen överenskommelse nås får medlemsstaten begära att ett förfarande inleds i syfte att medla mellan deras respektive ståndpunkter inom en tid av fyra månader; resultaten härav skall anges i en rapport, som skall överlämnas till och granskas av kommissionen innan ett beslut om att vägra finansiering fattas.
Kommissionen skall göra en bedömning av de belopp som skall undantas, särskilt med hänsyn till hur stor bristen på överensstämmelse är. Kommissionen skall beakta överträdelsens art och betydelse samt den ekonomiska förlust som gemenskapen lidit.
En vägran att finansiera får inte omfatta följande:
a) De utgifter som avses i artikel 2 och som verkställts före de tjugofyra månader som föregick kommissionens skriftliga meddelande till den berörda medlemsstaten om resultaten av kontrollerna.
b) De utgifter för åtgärder som avses i artikel 3 och där den slutliga betalningen verkställdes före de tjugofyra månader som föregick kommissionens skriftliga meddelande till den berörda medlemsstaten om resultaten av kontrollerna.
Bestämmelsen i femte stycket skall emellertid inte tillämpas på de ekonomiska följderna
a) av oegentligheter enligt artikel 8.2,
b) av statligt stöd eller överträdelser för vilka förfarandena som anges i artiklarna 88 och 226 i fördraget har inletts.
5. Tillämpningsföreskrifterna för denna artikel skall antas i enlighet med förfarandet i artikel 13. Dessa föreskrifter skall särskilt omfatta de förskottsbetalningar som avses i artikel 5.1 andra stycket under punkterna 2, 3 och 4 i denna artikel och förfarandena för de beslut som avses i nämnda punkterna 2, 3 och 4.
Artikel 8
1. Medlemsstaterna skall i enlighet med nationella bestämmelser i lagar och andra författningar vidta de åtgärder som är nödvändiga för att
a) försäkra sig om att transaktioner som finansieras av fonden verkligen äger rum och att de genomförs korrekt,
b) förhindra och ingripa mot oegentligheter,
c) indriva belopp som förlorats till följd av oegentligheter eller försumlighet.
Medlemsstaterna skall underrätta kommissionen om de åtgärder som vidtagits i dessa syften, särskilt i vilket stadium de förvaltningsmässiga och rättsliga förfarandena befinner sig.
2. Om en fullständigt indrivning inte kan åstadkommas skall de ekonomiska följderna av oegentligheter eller försumlighet bäras av gemenskapen, med undantag för följderna av sådana oegentligheter eller sådan försumlighet som kan tillskrivas medlemsstaternas myndigheter eller andra organ.
De indrivna beloppen skall betalas till de ackrediterade utbetalningsställena och dessa organ skall dra av de indrivna beloppen från de utgifter som fonden finansierar. Räntan på de belopp som drivits in eller som betalats för sent skall betalas in till fonden.
3. Rådet skall, på förslag av kommissionen, med kvalificerad majoritet fastställa de allmänna tillämpningsföreskrifterna för denna artikel.
Artikel 9
1. Medlemsstaterna skall till kommissionens förfogande ställa alla uppgifter som behövs för att fonden skall fungera väl och de skall även vidta alla lämpliga åtgärder för att underlätta den kontroll som kommissionen kan anse vara nödvändig inom ramen för förvaltningen av gemenskapsfinansieringen, inbegripet kontroller på plats.
Medlemsstaterna skall underrätta kommissionen om alla bestämmelser i lagar och andra författningar som de har antagit för tillämpningen av gemenskapens rättsakter avseende den gemensamma jordbrukspolitiken, i den mån dessa akter har ekonomiska följder för fonden.
2. Utan att det påverkar den kontroll som medlemsstaterna utför i enlighet med nationella bestämmelser i lagar och andra författningar och utan att det påverkar tillämpningen av bestämmelserna i artikel 248 i fördraget eller sådana kontroller som företas med stöd av artikel 279 c i fördraget skall företrädare som kommissionen utsett att genomföra kontroller på plats ha tillgång till alla böcker och andra handlingar, inbegripet uppgifter som upprättas eller lagras i elektronisk form, avseende utgifter som finansieras av fonden.
De får särskilt kontrollera
a) om förvaltningsrutinerna är förenliga med gemenskapsreglerna,
b) om de erforderliga underlagen finns och om dessa överensstämmer med de transaktioner som finansieras av fonden,
c) under vilka förhållanden transaktioner som finansieras av fonden genomförs och kontrolleras.
Kommissionen skall i god tid före kontrollen underrätta den berörda medlemsstaten eller den medlemsstat inom vars territorium kontrollen skall äga rum. Tjänstemän från den berörda medlemsstaten får delta i kontrollen.
På begäran av kommissionen och med medlemsstatens samtycke skall kontroller eller utredningar beträffande de transaktioner som avses i denna förordning utföras av den medlemsstatens behöriga myndigheter. Tjänstemän från kommissionen får också delta.
För att effektivisera kontrollen får kommissionen, med de berörda medlemsstaternas samtycke, ombesörja att myndigheter i dessa stater deltar i vissa kontroller eller utredningar.
3. Rådet skall vid behov, på förslag av kommissionen, med kvalificerad majoritet fastställa allmänna tilllämpningsföreskrifter för denna artikel:
Artikel 10
Före den 1 juli varje år skall kommissionen tillställa Europaparlamentet och rådet en finansiell rapport om förvaltningen av fonden under det föregående räkenskapsåret, särskilt dess ekonomiska ställning och utvecklingen av utgifternas storlek och utgiftsslagen samt förutsättningarna för gemenskapsfinansieringens genomförande.
Artikel 11
Kommittén för Europeiska utvecklings- och garantifonden för jordbruket (nedan kallad fondkommittén) skall bistå kommissionen med förvaltningen av fonden i enlighet med bestämmelserna i artiklarna 12-15.
Artikel 12
Fondkommittén skall bestå av företrädare för medlemsstaterna och för kommissionen. Varje medlemsstat skall i fondkommittén företrädas av högst fem tjänstemän. Ordförande för fondkommittén skall vara en företrädare för kommissionen.
Artikel 13
1. Om förfarandet i denna artikel skall tillämpas skall ordföranden, antingen på eget initiativ eller på begäran av en företrädare för en medlemsstat, hänskjuta ärendet till fondkommittén.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 205.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Medlemsstaternas röster skall vägas enligt den artikeln. Ordföranden får inte rösta.
3. a) Kommissionens beslut skall ha omedelbar verkan.
b) Om beslutet inte är förenligt med fondkommitténs yttrande skall kommissionens emellertid genast underrätta rådet. I sådana fall
- får kommissionen uppskjuta verkställandet av de beslutade åtgärderna under den tid som inte överstiger en månad från den dag då rådet underrättats.
- Rådet får inom den tidsfrist som anges i föregående strecksats fatta ett annat beslut med kvalificerad majoritet.
Artikel 14
1. Fondkommittén skall höras
a) i samtliga fall där det är föreskrivet att den skall höras,
b) angående den bedömning av fondens anslag som skall skrivas in i kommissionens upskattning för kommande budgetår och vid behov i ytterligare budgetsförslag,
c) om utkast till rapporter om fonden som skall överlämnas till rådet.
2. Fondkommittén får undersöka alla andra frågor som dess ordförande, antingen på eget initiativ eller på begäran av en företrädare för en medlemsstat, har hänskjutit till den.
Fondkommittén skall regelbundet informeras om fondens verksamheter.
Artikel 15
Ordföranden skall sammankalla fondkommittén.
Kommissionen skall ställa sekretariatstjänster till fondkommitténs förfogande.
Fondkommittén skall själv fastställa sin arbetsordning.
Artikel 16
1. Förordning (EEG) nr 729/70 skall upphävas.
2. Hänvisningar till den upphävda förordningen skall tolkas som hänvisningar till denna förordning och skall läsas i enlighet med jämförelsetabellen i bilagan.
Artikel 17
Artikel 15 tredje stycket och artikel 40 i beslut 90/424/EEG skall utgå.
Artikel 18
De åtgärder som krävs för att underlätta övergången från bestämmelserna i förordning (EEG) nr 729/70 till bestämmelserna i den här förordningen skall antas enligt förfarandet i artikel 13.
Artikel 19
Kommissionen får stryka första meningen i artikel 7.2 andra stycket enligt förfarandet i artikel 13, om de budgetmedel som beviljats fondens garantisektion och som finns tillgängliga i slutet av ett visst budgetår, gör det möjligt för fonden att finansiera de tilläggsutgifter som blir följden av strykningen för samma budgetår. Om kommissionen använder sig av denna befogenhet får den i enlighet med samma förfarande senarelägga startdatum till den 1 november för de betalningsperioder för åtgärder som påbörjas för att löpa mellan den 16 till och med den 31 oktober.
Artikel 20
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 1636/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 70/524/EEG av den 23 november 1970 om fodertillsatser(1), senast ändrat genom kommissionens förordning (EG) nr 1411/1999(2), särskilt artiklarna 9j och 3 i detta, och av följande skäl:
1. Enligt bestämmelserna i direktiv 70/524/EEG får nya fodertillsatser och nya användningsområden för fodertillsatser godkännas om detta verkar rimligt mot bakgrund av den vetenskapliga och tekniska utvecklingen.
2. Genom undantag från direktiv 70/524/EEG tillåts medlemsstaterna genom rådets direktiv 93/113/EG av den 14 december 1993 om användning och saluföring av enzymer och mikroorganismer och preparat av dessa i djurfoder(3), senast ändrat genom rådets direktiv 97/40/EG(4), att tillfälligt tillåta användning och saluföring av enzymer, mikroorganismer och preparat av dessa i foder.
3. Nya fodertillsatser eller nya användningsområden för fodertillsatser får ges ett provisoriskt godkännande om de vid den halt som tillåts i foder inte negativt påverkar människors eller djurs hälsa eller miljön, och inte heller skadar konsumenten genom att de förändrar animalieproduktens egenskaper, om deras förekomst i fodret kan kontrolleras, och om det är rimligt att anta - med hänsyn till tillgängliga resultat - att de har en positiv effekt på fodrets eller aminalieproduktionens egenskaper om de används i sådant foder.
4. Bestämmelserna i rådets direktiv 89/391/EEG av den 12 juni 1989(5) om åtgärder för att främja förbättringar av arbetstagarnas säkerhet och hälsa i arbetet och andra enskilda direktiv, särskilt rådets direktiv 90/679/EEG av den 26 november 1990(6) om skydd för arbetstagare mot risker vid exponering för biologiska agenser i arbetet, senast ändrat genom direktiv 97/65/EG(7), kan till fullo tillämpas när det gäller arbetstagare som handlar fodertillsatser.
5. En granskning av de akter som medlemsstaterna har överlämnat i enlighet med artikel 3 i direktiv 93/113/EG ger vid handen att vissa preparat av typen enzymer och mikroorganismer kan godkännas tills vidare.
6. Vetenskapliga foderkommittén har i ett yttrande fastställt att dessa preparat är ofarliga.
7. De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga foderkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De preparat av typen enzymer som förtecknas i bilaga I till denna förordning får godkännas som fodertillsatser i enlighet med direktiv 70/524/EEG på de villkor som anges i nämnda bilaga.
Artikel 2
Det preparat av typen enzymer som förtecknas i bilaga II till denna förordning får godkännas som fodertillsats i enlighet med direktiv 70/524/EEG på de villkor som anges i nämnda bilaga.
Artikel 3
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2376/1999
av den 9 november 1999
om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom kommissionens förordning (EG) nr 1835/1999(2), särskilt artikel 9 i denna, och
av följande skäl:
1. För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
2. I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
3. Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
4. Det är lämpligt att bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning fortfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3), senast ändrad genom rådets och Europaparlamentets förordning (EG) nr 955/1999(4), under en period av tre månader.
5. De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställas i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2562/1999
av den 3 december 1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 70/524/EEG av den 23 november 1970 om fodertillsatser(1), senast ändrat genom kommissionens förordning (EG) nr 2439/1999(2), särskilt artiklarna 9h.3 b och 9i.3 b i detta, och
av följande skäl:
1. På grund av den risk som dåliga plagiat av zootekniska tillsatser inom gemenskapen utgör för människors och djurs hälsa, skall enligt direktiv 70/524/EEG, ändrat genom rådets direktiv 96/51/EG(3), godkännandet av vissa grupper av tillsatser knytas till den som är ansvarig för avyttringen.
2. Efter den 31 december 1987 skall, särskilt enligt artikel 9h i direktiv 70/524/EEG, de preliminära godkännandena för tillsatser som avses i bilaga I och som hör till gruppen antibiotika och som förts över till bilaga B, kapitel II ersättas med godkännanden som knyts till den som är ansvarig för avyttringen för en tid av tio år.
3. Före den 1 april 1998 skall, särskilt enligt artikel 9i i direktiv 70/524/EEG, de preliminära godkännandena för tillsatser som avses i bilaga II och som hör till grupperna antibiotika och som förts över till bilaga B, kapitel III ersättas med godkännanden som knyts till den som är ansvarig för avyttringen.
4. För de tillsatser som förtecknas i bilagorna till den här förordningen har den som är ansvarig för den dokumentation utifrån vilken det tidigare godkännandet meddelades eller dennes efterträdare lämnat in nya ansökningar om godkännande. Ansökningarna för dessa tillsatser åtföljdes av erforderlig monografi och identitetsbeskrivning.
5. Godkännandet knyts till en person som är ansvarig för avyttringen på grundval av rent administrativa förfaranden och innebär inte någon ny utvärdering av tillsatserna. Även om godkännandena enligt denna förordning beviljas för en viss tid, kan de när som helst återkallas enligt artikel 9m och artikel 11 i direktiv 70/524/EEG. De kan särskilt återkallas mot bakgrund av följande: Vetenskapliga styrkommittén avgav den 28 maj 1999 ett yttrande om antimikrobiell resistens. Användningen av vissa antibiotika i foder håller för närvarande på att utvärderas på nytt enligt artikel 9g i direktiv 70/524/EEG. Sverige har på grundval av artikel 11 i direktiv 70/524/EEG inom sitt territorium förbjudit användningen av alla former av antibiotika som tillsats i foder. Kommissionen håller dessutom på att gå igenom de data som lämnats in och den mer allmänna frågan huruvida användningen av antibiotika som tillsats i foder uppfyller de villkor som föreskrivs i artikel 3a i direktiv 70/524/EEG för att godkännande som tillsats skall meddelas.
6. De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga foderkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De preliminära godkännandena av de tillsatser som förtecknas i bilaga I till denna förordning skall ersättas med ett godkännande som knyts till den som är ansvarig för avyttringen av tillsatserna och som anges i andra kolumnen i bilaga I.
Artikel 2
De preliminära godkännandena av de tillsatser som förtecknas i bilaga II till denna förordning skall ersättas med preliminära godkännanden som knyts till den som är ansvarig för avyttringen av tillsatserna och som anges i andra kolumnen i bilaga II.
Artikel 3
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
KOMMISSIONENS FÖRORDNING (EG) nr 2654/1999
av den 16 december 1999
om ändring av förordning (EEG) nr 2921/90 om beviljande av stöd för framställningen av kasein och kaseinater av skummjölk
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), särskilt artikel 15 i denna, och
av följande skäl:
1. Förordning (EG) nr 1255/1999 ersätter, från och med den 1 januari 2000, rådets förordning (EEG) nr 804/68(2), senast ändrad genom förordning (EG) nr 1587/96(3) och, bland andra, rådets förordning (EEG) nr 987/68 av den 15 juli 1968 om fastställande av allmänna bestämmelser om beviljande av stöd för skummjölk som förädlas till kasein eller kaseinater(4), senast ändrad genom förordning (EEG) nr 1435/90(5). För att ta hänsyn till denna nya ordning bör ändringar göras av bestämmelserna i kommissionens förordning (EEG) nr 2921/90 av den 10 oktober 1990 om beviljande av stöd för framställningen av kasein och kaseinater av skummjölk(6), senast ändrad genom förordning (EG) nr 2501/1999(7). Den förordningen bör kompletteras med definitioner av de produkter som berörs av denna stödordning och det bör preciseras till vilket organ ansökan om stöd skall lämnas. Dessa bestämmelser bör gälla från och med den 1 januari 2000.
2. Förvaltningskommittén för mjölk och mjölkprodukter har inte avgivit något yttrande inom den tid som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 1 i förordning (EEG) nr 2921/90 skall ändras på följande sätt:
a) skummjölk: mjölk från en eller flera kor eller getter, fri från tillsatser och som endast genomgått partiell skumning, så att fetthalten sjunkit till högst 0,10 %,
b) råkasein: den produkt, olöslig i vatten, som erhålls från skummjölk genom utfällning medelst syrning med bakteriekultur eller tillsats av syra, löpe eller andra mjölkkoagulerande enzymer, utan hänsyn till eventuell föregående jonbytes- eller koncentreringsbehandling,
c) kasein: den, i vatten olösliga, tvättade och torkade produkt som erhålls från råkasein eller skummjölk genom utfällning medelst syrning med bakteriekultur eller tillsats av syra, löpe eller andra mjölkkoagulerande enzymer, utan hänsyn till eventuell föregående jonbytes- eller koncentreringsbehandling,
d) kaseinater: de produkter som erhålls genom torkning av kasein eller råkasein som behandlats med neutraliserande agens."
Artikel 2
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
CENTRALGRUPPENS BESLUT
av den 22 mars 1999
om allmänna principer för ersättning till uppgiftslämnare och infiltratörer
(SCH/C (99) 25)
Infiltratörerna och uppgiftslämnarna bidrar med viktig hjälp i kampen mot den allvarliga brottsligheten över gränserna, i synnerhet narkotikabrottsligheten, eftersom dessa personer i allmänhet åtnjuter brottslingarnas förtroende och det med hjälp av dessa personer är möjligt att skaffa sig en allmän bild av verksamheten i de i små, enskilda enheter uppdelade brottsorganisationerna och kriminella strukturerna.
Arbetsgruppen för narkotikafrågor åtog sig detta ämne under det tyska ordförandeskapet och den har granskat rättsläget och rättspraxis i var och en a
KOMMISSIONENS BESLUT
av den 21 december 1999
om ändring av kommissionens beslut 93/436/EEG om särskilda villkor för import av fiskeriprodukter med ursprung i Chile
[delgivet med nr K(1999) 4749]
(Text av betydelse för EES)
(2000/61/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktionen och marknadsföringen av fiskeriprodukter(1), senast ändrat genom rådets direktiv 97/79/EG(2), särskilt artikel 11 i detta, och
2. Villkoren för import av musslor, tagghudingar, manteldjur och marina snäckor och sniglar med ursprung i Chile fastställs i kommissionens beslut 96/675/EG(5).
3. Hänvisningarna till lagstiftning i förlagan till sundhetsintyg i bilaga A till beslut 93/436/EEG innehåller vissa misstag och bör ändras.
4. De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga A till beslut 93/436/EEG skall ersättas med bilagan till det här beslutet.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 9 mars 2000
om att inte uppta monolinuron som ett verksamt ämne i bilaga I till rådets direktiv 91/414/EEG och om upphävande av tillstånd för växtskyddsmedel som innehåller detta verksamma ämne
[delgivet med nr K(2000) 656]
(Text av betydelse för EES)
(2000/234/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(1), senast ändrat genom kommissionens direktiv 97/73/EG(2),
med beaktande av kommissionens förordning (EEG) nr 3600/92 av den 11 december 1992 om närmare bestämmelser för genomförandet av den första etappen i det arbetsprogram som avses i artikel 8.2 i rådets direktiv 91/414/EEG om utsläppande av växtskyddsprodukter på marknaden(3), senast ändrad genom förordning (EG) nr 1199/97(4), särskilt artikel 7.3a led b i denna, och
av följande skäl:
(1) I kommissionens förordning (EG) nr 933/94(5), senast ändrad genom förordning (EG) nr 2230/95(6) anges verksamma ämnen i växtskyddsmedel, utses de rapporterande medlemsstaterna för genomförandet av kommissionens förordning (EEG) nr 3600/92 och fastställs anmälare för varje verksamt ämne.
(2) Monolinuron är ett av de 90 verksamma ämnen som omfattas av den första etappen av det arbetsprogram som fastställs i artikel 8.2 i rådets direktiv 91/414/EEG.
(3) I enlighet med artikel 7.1 c i förordning (EEG) nr 3600/92 ingav Förenade kungariket, som utsetts till rapporterande medlemsstat, den 30 april 1996 en rapport till kommissionen om sin utvärdering av de uppgifter som anmälarna lämnat enligt artikel 6.1 i den förordningen.
(4) Kommissionen och medlemsstaterna har granskat den ingivna rapporten inom Ständiga kommittén för växtskydd. I enlighet med bestämmelserna i artikel 7.6 i förordning (EEG) nr 3600/92 slutfördes denna granskning den 20 juli 1999 genom kommissionens granskningsrapport för monolinuron.
(5) Det framgår av de utvärderingar som gjorts att de uppgifter som lämnats inte visar att växtskyddsmedel som innehåller det verksamma ämnet i fråga uppfyller kraven enligt artikel 5.1 a, 5.1 b i direktiv 91/414/EEG.
(6) Den enda anmälaren har informerat kommissionen och den rapporterande medlemsstaten om att denne inte längre önskar delta i arbetsprogrammet för detta verksamma ämne. Viktiga delar av den information som krävs för att uppfylla kraven i direktiv 91/414/EEG kommer därför inte att överlämnas.
(7) Det är därför inte möjligt att uppta detta verksamma ämne i bilaga I till direktiv 91/414/EEG.
(8) Ett tidsbegränsat anstånd skall fastställas i enlighet med artikel 4.6 i direktiv 91/414/EEG under vilken tid kvarvarande lager får omhändertas, lagras, släppas ut på marknaden och användas.
(9) Detta beslut påverkar inte de eventuella åtgärder som kommissionen kan vidta i ett senare skede med hänsyn till detta verksamma ämne inom ramen för rådets direktiv 79/117/EEG(7).
(10) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för växtskydd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Monolinuron skall inte tas upp som ett verksamt ämne i bilaga I till direktiv 91/414/EEG.
Artikel 2
Medlemsstaterna skall garantera att
1. tillstånden för växtskyddsmedel som innehåller monolinuron upphävs inom en period på sex månader efter den dagen för anmälan av detta beslut,
2. inga tillstånd för växtskyddsmedel som innehåller monolinuron beviljas eller förnyas enligt undantaget i artikel 8.2 i direktiv 91/414/EEG från och med dagen för anmälan av detta beslut.
Artikel 3
Medlemsstaterna skall bevilja ett tidsbegränsat anstånd, under vilken tid kvarvarande lager får omhändertas, lagras, släppas ut på marknaden och användas i enlighet med artikel 4.6 i direktiv 91/414/EEG, som är så kort som möjligt och upphör inom 18 månader efter dagen för anmälan av detta beslut.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 25 juli 2000
om ändring av bilaga IV till rådets direktiv 90/539/EEG om djurhälsovillkor för handel inom gemenskapen med och för import från tredje land av fjäderfä och kläckningsägg och om ändring av beslut 96/482/EG om djurhälsovillkor och veterinärintyg för import från tredje land av fjäderfä och kläckningsägg, med undantag av strutsfåglar och ägg från strutsfåglar, inbegripet djurhälsoåtgärder som skall vidtas efter sådan import
[delgivet med nr K(2000) 2261]
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/539/EEG av den 15 oktober 1990 om djurhälsovillkor för handel inom, gemenskapen med och för import från tredje land av fjäderfä och kläckningsägg(1), senast ändrat genom rådets direktiv 1999/90/EG(2), särskilt artikel 23.1, artikel 24, artikel 26.2 samt artiklarna 27a och 34 i detta,
med beaktande av rådets direktiv 91/496/EEG av den 15 juli 1991 om fastställande av regler för hur veterinärkontroller skall organiseras för djur som importeras till gemenskapen från tredje land och om ändring av direktiven 89/662/EEG, 90/425/EEG och 90/675/EEG(3), senast ändrat genom direktiv 96/43/EG(4), särskilt artikel 10 i detta, och
av följande skäl:
(1) I kommissionens beslut 96/482/EG(5), senast ändrat genom beslut 1999/549/EG(6), fastställs djurhälsovillkor och veterinärintyg för import från tredje land av fjäderfä och kläckägg med undantag av strutsfåglar och ägg från strutsfåglar, inbegripet djurhälsoåtgärder som skall vidtas efter sådan import.
(2) Med hänsyn till de erfarenheter som gjorts vid tillämpningen av de föreskrivna åtgärderna bör villkoren för handel inom gemenskapen med dagsgamla kycklingar från kläckägg som importerats från tredje land ändras. Genom ändringen bör det bli möjligt för medlemsstaterna att sända dagsgamla kycklingar till anläggningar i en annan medlemsstat under förutsättning att kycklingarna isoleras efter import.
(3) Det är därför nödvändigt att ändra den förlaga till intyg som anges i bilaga IV till direktiv 90/539/EEG samt att ändra beslut 96/482/EG.
(4) Det är nödvändigt att den behöriga myndigheten i den avsändande medlemsstaten via Animo-systemet informerar den behöriga myndigheten på de dagsgamla kycklingarnas slutliga destinationsort om de djurhälsokrav avseende isoleringstid som skall tillämpas i dessa fall.
(5) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förlaga 2 i bilaga IV till direktiv 90/539/EEG skall ersättas med bilagan till detta beslut.
Artikel 2
Följande skall läggas till i artikel 3.1 i beslut 96/482/EG:"Om dagsgamla kycklingar inte föds upp i den medlemsstat till vilken kläckäggen importerats skall de direkt transporteras till och förvaras på den anläggning som avses i punkt 9.2 i förlaga 2 till hälsointyg i bilaga IV till rådets direktiv 90/539/EEG under åtminstone tre veckor från kläckningsdagen."
Artikel 2
Detta beslut gäller för sändningar av dagsgamla kycklingar för vilka det utfärdas intyg från och med den 1 oktober 2000.
Artikel 4
Detta beslut riktar sig till alla medlemsstater.
Kommissionens beslut
av den 26 juli 2000
enligt Europaparlamentets och rådets direktiv 95/46/EG om huruvida ett adekvat skydd säkerställs genom de principer om integritetsskydd (Safe Harbor Privacy Principles) i kombination med frågor och svar som Förenta staternas handelsministerium utfärdat
(2000/520/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter(1), särskilt artikel 25.6 i detta, och
av följande skäl:
(1) Enligt direktiv 95/46/EG skall medlemsstaterna föreskriva att överföring av personuppgifter till tredje land endast får ske om ifrågavarande tredje land säkerställer en adekvat skyddsnivå och om medlemsstatens lagar genom vilka andra bestämmelser i direktivet genomförs, efterlevs före överföringen.
(2) Kommissionen kan konstatera att ett tredje land har en adekvat skyddsnivå. I sådana fall får personuppgifter överföras från medlemsstaterna utan att det behövs några ytterligare garantier.
(3) Enligt direktiv 95/46/EG skall bedömningen av skyddsnivån ske på grundval av alla de förhållanden som har samband med en överföring eller en grupp överföringar av uppgifter och vissa omständigheter skall särskilt beaktas. Arbetsgruppen för skydd av enskilda med avseende på behandling av personuppgifter som inrättats genom det direktivet(2) har utfärdat riktlinjer för hur sådana beddömningar skall göras(3).
(4) Mot bakgrund av de olika sätten att se på frågan om uppgiftsskydd i olika tredje länder bör bedömningen av om skyddsnivån är adekvat ske, och beslut som grundar sig på artikel 25.6 i direktiv 95/46/EG verkställas, utan godtycklig eller obefogad diskriminering i förhållande till tredje land eller mellan tredje länder där liknande förhållanden råder och så att det inte utgör ett dolt handelshinder. Härvid bör hänsyn tas till gemenskapens nuvarande internationella åtaganden.
(5) Den adekvata skyddsnivån för överföring av uppgifter från gemenskapen till Förenta staterna i enlighet med detta beslut bör anses ha uppnåtts om organisationer följer Safe Harbor Privacy-principerna för skydd av personuppgifter som överförs från en medlemsstat till Förenta staterna (nedan kallade principerna) och de vägledande frågorna och svaren (nedan kallade FoS) som utfärdats av Förenta staternas regering den 21 juli 2000. Organisationerna bör dessutom offentliggöra sin politik för skydd av personuppgifter och vara underställda antingen Federal Trade Commission (FTC) enligt avsnitt 5 i Federal Trade Commission Act, som förbjuder illojala eller bedrägliga handlingar eller metoder i handeln och i verksamhet som påverkar handeln, eller någon annan tillsynsmyndighet som på ett effektivt sätt ser till att principerna, tillämpade i överensstämmelse med FoS, efterlevs.
(6) Områden och/eller databehandling som inte lyder under någon av de myndigheter i Förenta staterna som anges i bilaga VII till detta beslut bör inte omfattas av beslutet.
(7) För att se till att detta beslut tillämpas korrekt är det nödvändigt att de organisationer som ansluter sig till principerna och FoS kan erkännas av berörda parter, t.ex. de registrerade, exportörer av uppgifter och dataskyddsmyndigheter. I detta syfte bör Förenta staternas handelsministerium, eller det organ som ministeriet bestämmer, förbinda sig att föra och göra tillgänglig för allmänheten en förteckning över de organisationer som förpliktat sig att följa principerna i överensstämmelse med FoS och som lyder under åtminstone en av de myndigheter som nämns i bilaga VII till detta beslut.
(8) För att värna om öppenhet och för att bevara förmågan hos de behöriga myndigheterna i medlemsstaterna att garantera skydd av enskilda med avseende på behandlingen av deras personuppgifter är det nödvändigt att i detta beslut specificera vilka omständigheter som i undantagsfall bör medföra att vissa dataflöden avbryts, trots att skyddsnivån befunnits vara adekvat.
(9) Systemet med safe harbor sådant det utformats enligt principerna och FoS kan behöva ses över i ljuset av erfarenheter från utveckling på integritetsskyddets område under förhållanden då tekniken ständigt gör det lättare att överföra och behandla personuppgifter och i ljuset av rapporter om genomförande av berörda tillsynsmyndigheter.
(10) Arbetsgruppen för skydd av enskilda med avseende på behandling av personuppgifter som inrättats genom artikel 29 i direktiv 95/46/EG har avgivit yttranden om den skyddsnivå som erbjuds av safe harbor-principerna i Förenta staterna, och vid utarbetandet av föreliggande beslut har hänsyn tagits till dessa yttranden(4).
(11) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som inrättats genom artikel 31 i direktiv 95/46/EG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Med avseende på artikel 25.2 i direktiv 95/46/EG skall i fråga om all verksamhet som omfattas av det direktivet, safe harbor-principerna om integritetsskydd (nedan kallade principerna), se bilaga I till detta beslut, tillämpade i enlighet med den vägledning som ges i de frågor och svar (nedan kallade FoS) som utfärdats av Förenta staternas handelsministerium den 21 juli 2000, se bilaga II till detta beslut, anses utgöra en adekvat skyddsnivå för personuppgifter som överförs från gemenskapen till organisationer som är etablerade i Förenta staterna med beaktande av följande dokument som utfärdats av Förenta staternas handelsministerium:
a) En översikt över genomförandet av safe harbor, bilaga III.
b) Ett memorandum om ersättning vid kränkning av enskildas integritet och uttryckliga behörigheter i Förenta staternas lagstiftning, bilaga IV.
c) En skrivelse från Federal Trade Commission, bilaga V.
d) En skrivelse från Förenta staternas transportministerium, bilaga VI.
2. I samband med varje överföring av uppgifter skall följande villkor vara uppfyllda:
a) Den organisation som tar emot uppgifterna har otvetydigt och offentligt förpliktat sig att följa principerna såsom de tillämpas i enlighet med FoS, och
b) denna organisation omfattas av de lagstadgade befogenheter som tillkommer någon av de myndigheter i Förenta staterna som anges i bilaga VII till detta beslut och som är bemyndigade att handlägga klagomål och ge upprättelse vid användning av illojala och bedrägliga metoder och att utverka skadestånd åt enskilda, oberoende av deras bosättningsland eller nationalitet, om principerna inte följs i överensstämmelse med FoS.
3. De villkor som anges i punkt 2 skall anses vara uppfyllda för varje organisation som genom självcertifiering förbinder sig att följa principerna i överensstämmelse med FoS från den dag då organisationen underrättar Förenta staternas handelsministerium, eller det organ som ministeriet bestämmer, om offentliggörandet av den förpliktelse som avses i punkt 2 a och om namnet på den myndighet som avses i punkt 2 b.
Artikel 2
Detta beslut gäller endast frågan om den skyddsnivå är adekvat som enligt principerna och FoS erbjuds i Förenta staterna, i förhållande till de krav som ställs i artikel 25.1 i direktiv 95/46/EG, och det påverkar inte tillämpningen av andra bestämmelser i det direktivet som gäller behandling av personuppgifter inom medlemsstaterna, särskilt artikel 4 i direktivet.
Artikel 3
1. Utan att det påverkar de befogenheter behöriga myndigheter i medlemsstaterna har att vidta åtgärder för att säkra efterlevnaden av nationella bestämmelser som antagits enligt andra bestämmelser i direktiv 95/46/EG än artikel 25, får dessa myndigheter utöva sin befogenhet att tillfälligt förbjuda överföringen av uppgifter till en organisation som genom självcertifiering förbundit sig att följa principerna i överensstämmelse med FoS, i syfte att skydda enskilda med avseende på behandling av deras personuppgifter i de fall då
a) den myndighet i Förenta staterna som avses i bilaga VII till detta beslut eller en sådan oberoende instans för handläggning av klagomål som avses under a i avsnittet om kontroll av efterlevnaden i bilaga I till detta beslut, har funnit att organisationen agerar i strid med principerna tillämpade i överensstämmelse med FoS, eller
b) det är i hög grad sannolikt att principerna överträds, det finns välgrundad anledning att tro att den berörda instansen för handläggning av klagomål inte vidtar och inte i rätt tid kommer att vidta de åtgärder som behövs för att lösa problemet, en fortsatt överföring av uppgifterna skulle innebära en överhängande risk för allvarlig skada för registrerade, och de behöriga myndigheterna i medlemsstaten har gjort vad som under rådande omständigheter rimligvis kan krävas för att anmärka mot organisationen och ge den tillfälle att gå i svaromål.
Förbudet skall hävas så snart det säkerställts att organisationen följer principerna i överensstämmelse med FoS och de behöriga myndigheterna i Europeiska unionen har underrättats härom.
2. Medlemsstaterna skall utan dröjsmål underrätta kommissionen om åtgärder som vidtagits med stöd av punkt 1.
3. Medlemsstaterna och kommissionen skall även underrätta varandra om varje fall där en myndighet, som är ansvarig för att principerna tillämpade i överensstämmelse med FoS följs i Förenta staterna, inte kunnat säkerställa detta.
4. Om den information som inhämtats i enlighet med punkterna 1, 2 och 3 visar att någon av de myndigheter som har ansvar för att principerna tillämpade i överensstämmelse med FoS följs i Förenta staterna inte fullgör denna uppgift på ett effektivt sätt, skall kommissionen underrätta Förenta staternas handelsministerium om detta och vid behov lägga fram förslag till bestämmelser i enlighet med det förfarande som föreskrivs i artikel 31 i direktivet i syfte att helt eller tills vidare upphäva detta beslut eller begränsa dess tillämpningsområde.
Artikel 4
2. Kommissionen skall om så behövs föreslå åtgärder i enlighet med det förfarande som föreskrivs i artikel 31 i direktivet.
Artikel 5
Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att följa detta beslut senast nittio dagar efter det att beslutet har delgivits medlemsstaterna.
Artikel 6
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 6 september 2000
om ett principiellt erkännande av fullständigheten hos den dokumentation som inlämnats för detaljerad granskning inför ett eventuellt införande av RH-7281 (zoxamid) och B-41; E-187 (milbemectin), BAS500F (pyraclostrobin) och AEF130360 (foramsulfuron) i bilaga I till rådets direktiv 91/414/EEG om utsläppande av växtskyddsmedel på marknaden
[delgivet med nr K(2000) 2285]
(2000/540/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(1), senast ändrat genom kommissionens direktiv 2000/10/EG(2), särskilt artikel 6.3 i detta, och
av följande skäl:
(1) I direktiv 91/414/EEG (nedan kallat direktivet) föreskrivs att en gemenskapsförteckning skall upprättas över verksamma ämnen som får användas i växtskyddsmedel.
(2) Företaget Rohm & Haas France SA lämnade den 2 juni 1999 in en akt med dokumentation för det verksamma ämnet RH-7281 (zoxamid) till myndigheterna i Förenade kungariket för införande av detta verksamma ämne i bilaga I till direktivet.
(3) Företaget Sankyo Company Limited lämnade den 6 mars 2000 in en akt med dokumentation för det verksamma ämnet B-41; E-187 (milbemectin) till de nederländska myndigheterna.
(4) Företaget BASF AG lämnade den 28 februari 2000 in en akt med dokumentation för det verksamma ämnet BAS500F (pyraclostrobin) till de tyska myndigheterna.
(5) Företaget Aventis GmbH lämnade den 30 mars 2000 in en akt med dokumentation för det verksamma ämnet AEF130360 (foramsulfuron) till de tyska myndigheterna.
(6) Myndigheterna i fråga underrättade kommissionen om resultaten av en första undersökning av huruvida dokumentationen var fullständig vad gäller kraven på uppgifter och upplysningar enligt bilaga II och, vad beträffar åtminstone ett växtskyddsmedel som innehåller det verksamma ämnet i fråga, enligt bilaga III till direktivet. I enlighet med artikel 6.2 överlämnade de ansökande företagen därefter akterna till kommissionen och övriga medlemsstater.
(7) Akterna för RH-7281 (zoxamid), B-41; E-187 (milbemectin), BAS500F (pyraclostrobin) och AEF130360 (foramsulfuron) remitterades till Ständiga kommittén för växtskydd den 31 maj 2000.
(8) Enligt artikel 6.3 i direktivet krävs en bekräftelse på gemenskapsnivå av att varje akt med dokumentation uppfyller kraven på faktauppgifter och upplysningar enligt bilaga II och, vad beträffar åtminstone ett växtskyddsmedel som innehåller det verksamma ämnet i fråga, enligt bilaga III till direktivet.
(9) En sådan bekräftelse är nödvändig för att en detaljerad granskning av dokumentationen skall kunna äga rum. Den skall också göra det möjligt för medlemsstaterna att tills vidare godkänna växtskyddsmedel som innehåller det verksamma ämnet i fråga, med beaktande av de villkor som anges i artikel 8.1 i direktivet, särskilt villkoret om att en detaljerad utvärdering av de verksamma ämnena och av växtskyddsmedlen skall göras i enlighet med direktivets bestämmelser.
(10) Ett sådant beslut hindrar inte att ytterligare faktauppgifter och upplysningar kan komma att begäras in från de ansökande företagen för att klargöra vissa punkter i den dokumentation som lagts fram. Då den rapporterande medlemsstaten begär in sådana upplysningar som är nödvändiga för att klargöra innehållet i dokumentationen skall detta inte påverka tidsfristen för inlämnande av den rapport som avses i skäl 12.
(11) Medlemsstaterna och kommissionen har enats om att Förenade kungariket skall fortsätta att noggrant granska dokumentationen om RH-7281 (zoxamid), att Nederländerna skall fortsätta att noggrant granska dokumentationen om B-41; E-187 (milbemectin) och att Tyskland skall fortsätta att noggrant granska dokumentationen om BAS500F (pyraclostrobin) och AEF130360 (foramsulfuron).
(12) Förenade kungariket, Nederländerna och Tyskland skall rapportera resultaten av sina undersökningar till kommissionen, och samtidigt ge rekommendationer om huruvida införande bör beviljas eller inte, samt även ange eventuella villkor för införande senast inom ett år efter det att detta beslut har offentliggjorts.
(13) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för växtskydd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Med hänsyn till de föreslagna användningsområdena uppfyller följande akter med dokumentation i princip de krav beträffande uppgifter och upplysningar som anges i bilaga II och, vad beträffar minst ett växtskyddsmedel som innehåller det verksamma ämnet i fråga, i bilaga III till direktivet:
1. Den dokumentation som lämnats in av Rohm & Haas France SA till kommissionen och medlemsstaterna beträffande införandet av RH-7281 (zoxamid) som ett verksamt ämne i bilaga I till direktiv 91/414/EEG, och som överlämnades till Ständiga kommittén för växtskydd den 31 maj 2000.
2. Den dokumentation som lämnats in av Sankyo Company Limited till kommissionen och medlemsstaterna beträffande införandet av B-41; E-187 (milbemectin) som ett verksamt ämne i bilaga I till direktiv 91/414/EEG, och som överlämnades till Ständiga kommittén för växtskydd den 31 maj 2000.
3. Den dokumentation som lämnats in av BASF AG till kommissionen och medlemsstaterna beträffande införandet av BAS500F (pyraclostrobin) som ett verksamt ämne i bilaga I till direktiv 91/414/EEG, och som överlämnades till Ständiga kommittén för växtskydd den 31 maj 2000.
4. Den dokumentation som lämnats in a
Europaparlamentets och rådets direktiv 2000/13/EG
av den 20 mars 2000
om tillnärmning av medlemsstaternas lagstiftning om märkning och presentation av livsmedel samt om reklam för livsmedel
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 95 i detta,
med beaktande av kommissionens förslag,
med beaktande av Ekonomiska och sociala kommitténs yttrande(1),
i enlighet med det förfarande som anges i artikel 251 i fördraget(2) och
av följande skäl:
(1) Rådet direktiv 79/112/EEG av den 18 december 1978 om tillnärmning av medlemsstaternas lagstiftning om märkning och presentation av livsmedel samt om reklam för livsmedel(3) har undergått flera och omfattande ändringar(4). För att skapa klarhet och av rationella skäl bör därför en kodificering företas av nämnda direktiv.
(2) Skillnader mellan medlemsstaternas lagar och andra författningar om märkning av livsmedel kan hämma den fria rörligheten av dessa varor och kan leda till ojämlika konkurrensvillkor.
(3) Det är därför nödvändigt att närma dessa lagstiftningar till varandra för att bidra till att den inre marknaden fungerar smidigare.
(4) Syftet med detta direktiv bör vara att anta allmänna gemenskapsregler som skall gälla horisontellt för alla livsmedel som släpps ut på marknaden.
(5) Specialregler som tillämpas vertikalt endast på vissa livsmedel bör fastställas inom ramen för de bestämmelser som behandlar dessa varor.
(6) Det huvudsakliga syftet med regler om märkning av livsmedel bör vara behovet att informera och skydda konsumenten.
(7) Detta behov innebär att medlemsstaterna, med hänsyn tagen till bestämmelserna i fördraget, skall kunna ställa språkliga krav.
(8) Detaljerad märkning för att ange produktens exakta art och beskaffenhet gör det möjligt för konsumenten att göra sitt val med full sakkännedom och är det lämpligaste eftersom det medför minsta möjliga hinder för den fria handeln.
(9) En förteckning bör därför göras upp över alla uppgifter som i princip bör framgå av märkningen på alla livsmedel.
(10) Med hänsyn till att detta direktiv är horisontellt var det från början inte möjligt att bland de obligatoriska märkningsanvisningarna ta med samtliga uppgifter som gäller för varje livsmedel och som måste framgå av den förteckning som i princip gäller för samtliga livsmedel; i ett senare steg bör gemenskapsbestämmelser antas som kompletterar de bestämmelser som redan finns.
(11) Medlemsstaterna bör vidare, om det saknas specialregler inom gemenskapen, behålla rätten att fastställa vissa nationella bestämmelser som komplement till de allmänna bestämmelserna i detta direktiv, dock bör dessa bestämmelser vara underkastade en gemenskapsprocedur.
(12) En sådan procedur måste utgöras av ett gemenskapsbeslut, när en medlemsstat önskar att införa ny lagstiftning.
(13) Bestämmelser måste också skapas för att ge gemenskapens lagstiftare möjlighet att, i undantagsfall, avvika från vissa förpliktelser som har fastställts generellt.
(14) Reglerna för märkning bör också förbjuda användning av information som skulle kunna vilseleda köparen eller som tillskriver livsmedel hälsobringande egenskaper; detta förbud bör för att vara verksamt gälla också presentation av och reklam för livsmedel.
(15) I syfte att underlätta handeln mellan medlemsstaterna får det i handelsleden före försäljningen till konsumenter tillåtas att endast den viktigaste informationen framgår av den yttre förpackningen och att vissa obligatoriska uppgifter som måste finnas på ett färdigförpackat livsmedel behöver framgå endast av handelsdokument som rör detta.
(16) Medlemsstaterna bör behålla rätten att, beroende på lokala förhållanden och praktiska omständigheter, fastställa regler för märkning av livsmedel som säljs i lös vikt; informationen bör i sådana fall likväl göras tillgänglig för konsumenten.
(17) För att förenkla och påskynda förfarandet bör kommissionen anförtros uppgiften att besluta om verkställighetsåtgärder av teknisk natur.
(18) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(5).
(19) Detta direktiv får inte påverka medlemsstaternas förpliktelser vad gäller de tidsgränser för genomförande av direktiven som anges i bilaga IV del B.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Detta direktiv gäller även livsmedel avsedda för restauranger, sjukhus; personalrestauranger och andra liknande storkök (i det följande benämnda storkök).
3. I detta direktiv avses med
a) märkning: varje ord, uppgift, varumärke, märkesnamn, illustration eller symbol i samband med livsmedel som anbringas på förpackning, dokument, meddelande, etikett, ring eller hylsa som medföljer eller avser sådant livsmedel,
b) färdigförpackat livsmedel: varje enskild vara som i oförändrat skick är avsedd att tillhandahållas konsumenter och storkök och som består av ett livsmedel och den förpackning i vilket det placerades innan det erbjöds till försäljning, oavsett om förpackningen omsluter livsmedlet helt eller endast delvis, men förutsatt att förpackningen omsluter livsmedlet på sådant sätt att innehållet inte kan ändras utan att förpackningen öppnas eller ändras.
Artikel 2
1. Märkningen och dess närmare utformning får inte
a) vara sådan att den på ett avgörande sätt skulle kunna vilseleda köparen, i synnerhet
i) om vad som är utmärkande för livsmedlet, särskilt dess slag, identitet, egenskaper, sammansättning, kvantitet, hållbarhet, ursprung eller härkomst, framställnings- eller produktionsmetod,
ii) genom att tillskriva livsmedlet verkningar eller egenskaper som det inte har,
iii) genom att antyda att livsmedlet har speciella egenskaper, då i själva verket alla liknande livsmedel har sådana egenskaper,
b) såvida något annat inte följer av gemenskapsbestämmelser för naturliga mineralvatten och specialdestinerade livsmedel, tillskriva livsmedel egenskaper som förebygger, behandlar eller botar någon sjukdom hos människor eller antyda sådana egenskaper.
2. Rådet skall på det sätt som anges i artikel 95 i fördraget, upprätta en icke uttömmande förteckning över sådana påståenden som avses i punkt 1 och vilkas användning i alla händelser måste förbjudas eller begränsas.
3. De förbud och begränsningar som avses i punkterna 1 och 2 skall gälla också
a) presentationen av livsmedel, särskilt med avseende på deras form, utseende eller förpackning, de förpackningsmaterial som används och det sätt på vilket livsmedlen arrangeras samt den miljö i vilken de exponeras,
b) reklam.
Artikel 3
1. Om något annat inte följer av artiklarna 4-17, är endast följande uppgifter obligatoriska vid märkning av livsmedel:
1. Det namn under vilket varan säljs.
2. Ingrediensförteckning.
3. Mängden av särskilda ingredienser eller kategorier av ingredienser i enlighet med bestämmelserna i artikel 7.
4. Nettokvantitet i fråga om färdigförpackade livsmedel.
5. Datum för minsta hållbarhetstid eller, när det gäller livsmedel som ur mikrobiologisk synpunkt är lättfördärvliga, datum för sista förbrukningsdag.
6. Speciella förvarings- eller användningsanvisningar.
7. Förpackarens eller tillverkarens namn eller firma samt adress eller uppgift om säljare som är etablerad inom gemenskapen.
Medlemsstaterna skall dock ha rätt att i fråga om smör som framställts inom deras territorium, kräva uppgift endast om tillverkaren, förpackaren eller säljaren.
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt andra stycket.
8. Uppgift om den plats där livsmedlet är producerat eller varifrån det kommer i fall då underlåtenhet att lämna sådana uppgifter kan vilseleda konsumenten i fråga om livsmedlets rätta ursprung eller härkomst.
9. Bruksanvisning, om det utan en sådan skulle vara omöjligt att använda livsmedlet på rätt sätt.
10. För drycker som innehåller mer än 1,2 volymprocent alkohol, den verkliga alkoholhalten uttryckt i volym.
2. Utan hinder av punkt 1 får medlemsstaterna behålla nationella bestämmelser som föreskriver att tillverkaren eller förpackaren skall anges, såvitt avser deras nationella livsmedelsproduktion.
3. Bestämmelserna i denna artikel skall inte påverka tillämpningen av mer precisa eller långtgående bestämmmelser om mått och vikt.
Artikel 4
1. Gemenskapsbestämmelser som gäller endast för vissa livsmedel och inte livsmedel i allmänhet får i särskilda fall avvika från de krav som fastställs i artikel 3.1 punkterna 2 och 5, under förutsättning att detta inte leder till att köparen blir bristfälligt informerad.
3. De gemenskapsbestämmelser som avses i punkterna 1 och 2 skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
Artikel 5
1. Det namn under vilket ett livsmedel säljs skall vara det namn som förbehållits livsmedlet i gemenskapens bestämmelser för livsmedlet.
a) Om gemenskapen saknar bestämmelser skall försäljningsnamnet vara det namn som föreskrivs i lag eller andra författningar som gäller i den medlemsstat i vilken varan säljs till konsumenter eller till institutioner och storkök.
Om försäljningsnamn saknas skall det namn under vilket varan säljs vara det namn som är vedertaget i den medlemsstat i vilken den säljs till konsumenter eller institutioner och storkök, eller en beskrivning av livsmedlet och om det behövs av dess användning, vilket skall vara tillräckligt klargörande för att informera köparen om livsmedlets verkliga art och göra det möjligt för köparen att särskilja det från andra varor som det skulle kunna förväxlas med.
b) Det skall också vara tillåtet att i den medlemsstat där livsmedlet saluförs använda det namn under vilken produkten tillverkas och saluförs i den medlemsstat där tillverkningen sker.
I fall där övriga bestämmelser i detta direktiv, särskilt de i artikel 3, inte är tillräckliga för att säkerställa att konsumenterna i den medlemsstat där produkten saluförs har kännedom om produktens verkliga art och kan särskilja det från produkter som det skulle kunna förväxlas med, skall försäljningsnamnet emellertid kompletteras med ytterligare beskrivande information bredvid namnet.
c) I undantagsfall får försäljningsnamnet i den medlemstat där tillverkningen sker inte användas i den medlemsstat där saluföringen sker, när den produkt som betecknas i fråga om sammansättning eller framställning skiljer sig så mycket från den produkt som är känd under det namnet att bestämmelserna i punkt b inte är tillräckliga för att säkerställa att konsumenterna i den medlemsstat där varan saluförs ges korrekt information.
2. Inget varumärke, märkesnamn eller fantasinamn får användas i stället för det namn under vilket varan säljs.
3. Det namn under vilket varan säljs skall omfatta eller åtföljas av uppgifter om livsmedlets fysiska tillstånd eller den särskilda behandling som livsmedlet fått (t.ex. pulvrisering, frystorkning, djupfrysning, koncentrering, rökning) i samtliga fall då avsaknaden av sådan information skulle kunna skapa förvirring hos köparen.
Alla livsmedel som har behandlats med joniserande strålning skall förses med någon av följande uppgifter:
- på spanska:
"irradiado" eller "tratado con radiación ionizante"
- på danska:
"bestrålet/..." eller "strålekonserveret" eller "behandlet med ioniserende stråling" eller "konserveret med ioniserende stråling"
- på tyska:
"bestrahlt" eller "mit ionisierenden Strahlen behandelt".
- på engelska:
"irradiated" eller "treated with ionizing radiation"
- på franska:
"traité par rayonnements ionisants" eller "traité par ionisation."
- på italienska:
"irradiato" eller "trattato con radiazioni ionizzanti"
- på nederländska:
"doorstraald" eller "door bestraling behandeld" eller "met ioniserende stralen behandeld"
- på portugisiska:
"irradiado" eller "tratado por irradiação" eller "tratado por radiação ionizante".
- på finska:
"säteilytetty" eller "käsitelty ionisoivalla säteilyllä"
- på svenska:
"bestrålad" eller "behandlad med joniserande strålning."
Artikel 6
1. Ingredienser skall anges i enlighet med denna artikel och bilagorna I, II och III.
2. Ingredienser behöver inte anges beträffande
a) - färsk frukt och färska grönsaker, inklusive potatis, som inte skalats, delats i bitar elelr behandlats på liknande sätt,
- kolsyrat vatten, om det framgår av försäljningsnammet att vattnet har kolsyrats,
- mikrobiellt framställd ättika som utvunnits ur en enda basprodukt coh som inte fillsatts någon annan ingrediens,
b) - ost,
- smör,
- kulturmjölk och syrad grädde,
förutsatt att ingen ingrediens har tillsatts utom mjölkprodukter, enzymer och kulturer av mikroorganismer som är nödvändiga för framställningen, eller det salt som behövs för framställning av annan ost än färskost och smältost,
c) varor som består av en enda ingrediens
- om försäljningsnamnet är identiskt med nammet på ingrediensen, eller
- om ingrediensen klart framgår av försäljningsnamnet utan risk för förväxling.
3. I fråga om drycker som innehåller mer än 1,2 volymprocent alkohol skall rådet på förslag av kommissionen före den 22 december 1982, bestämma reglerna för hur ingredienser skall anges.
4. a) Med ingrediens menas varje ämne, inklusive tillsatser, som använts i tillverkningen eller beredningen av ett livsmedel och som finns kvar i den färdiga produkten, om än i annan form.
b) Om en ingrediens i ett livsmedel består av flera ingredienser, skall dessa anses som ingredienser i det aktuella livsmedlet.
c) Som ingredienser anses inte
i) beståndsdelarna av en ingrediens som under framställningsprocessen tillfälligt avskiljts men senare åter tillförts livsmedlet i proportioner som inte överskrider de ursprungliga,
ii) tillsatser
- vilkas förekomst i ett visst livsmedel uteslutande beror på att de ingått i en eller flera ingredienser i det aktuella livsmedlet, förutsatt att tillsatserna inte har någon teknisk funktion i den färdiga varan,
- som används som processhjälpmedel,
iii) ämnen som används i de mängder som är absolut nödvändiga som lösningsmedel för tillsatser eller aromämnen.
d) Enligt der förfarande som fastställs i artikel 20.2 kan det i vissa fall avgöras huruvida villkoren i c ii och iii är uppfyllda.
5. Ingrediensförteckningen skall omfatta samtliga ingredienser i livsmedlet i fallande storleksordning efter den vikt som ingrediensen hade vid framställningstidpunkten. Den skall föregås av en lämplig rubrik som innehåller ordet "ingredienser".
Undantag:
- Tillsatt vatten och flyktiga ämnen skall anges i storleksordning efter vikt i den färdiga varan; den mängd vatten som tillsatts som ingrediens i ett livsmedel skall beräknas genom att den färdiga varans totala mängd minskas med den totala mängden av övriga använda ingredienser. Denna mängd behöver inte beaktas om den inte överstiger 5 % av den färdiga varans vikt.
- Ingredienser som använts i koncentrerad eller torkad form och som under framställningen rekonstitueras får anges i storleksordning efter den vikt som ingredienserna hade innan de koncentrerades eller torkades.
- Ingredienserna i koncentrerade eller torkade livsmedel som är avsedda att rekonstitueras genom tillsats av vatten får anges efter proportion i den rekonstituerade varan, förutsatt att ingrediensförteckningen åtföljs av uttrycket "ingredienser i den rekonstituerade varan" eller "ingredienser i den konsumtionsfärdiga varan" eller liknande uttryck.
- Ingredienserna i frukt eller grönsaksblandningar, i vilka ingen särskild frukt eller grönsak påtagligt dominerar med hänsyn till vikt får anges i annan ordning, förutsatt att denna ingrediensförteckning åtföljs av uttrycket "i varierande proportion" eller liknande uttryck.
- Ingredienserna i krydd- eller örtblandningar, i vilka ingen krydda eller ört påtagligt dominerar med hänsyn till vikt får anges i annan ordning, förutsatt att ingrediensförteckningen följs av uttrycket "i varierande proportion" eller liknande uttryck.
6. Ingredienser skall vid behov anges med sina särskilda beteckningar i enlighet med de regler som fastställts i artikel 5.
Undantag:
- Ingredienser som tillhör någon av de i bilaga 1 uppräknade kategorierna och som är beståndsdelar i ett annat livsmedel, behöver anges endast med namnet på denna kategori.
Förteckningen över kategorier i bilaga I kan ändras i enlighet med förfarandet i artikel 20.2.
Beteckningen "stärkelse" i bilaga I måste dock alltid kompletteras med en angivelse av vilken specifik växt den framställts ur, då denna ingrediens kan innehålla gluten.
- Ingredienser som tillhör någon av de i bilaga II uppräknade kategorierna skall alltid anges med namnet på denna kategori åtföljt av deras särskilda beteckning eller E-nummer. Om en ingrediens tillhör mer än en av kategorierna skall den kategori anges som är lämpligast med hänsyn till ingrediensens huvudsakliga funktion i det aktuella livsmedlet.
Ändringar av nämnda bilaga som grundas på framsteg när det gäller vetenskapligt eller tekniskt kunnande skall antas i enlighet med förfarandet i artikel 20.2.
Beteckningen "modifierad stärkelse" i bilaga II måste dock alltid kompletteras med en angivelse av vilken specifik växt den framställs ur, då denna ingrediens kan innehålla gluten.
- Aromer skall benämnas enligt bilaga III.
- De särskilda gemenskapsbestämmelserna om angivelse av behandling av en ingrediens med joniserande strålning skall antas senare i enlighet med artikel 95 i fördraget.
7. Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser, får fastställa att det namn, som ett visst livsmedel säljs under, skall åtföljas av uppgift om en eller flera särskilda ingredienser.
Det förfarande som fastställs i artikel 19 skall tillämpas på varje sådan nationell bestämmelse.
De gemenskapsbestämmelser som avses i denna punkt skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
8. I det fall som avses i punkt 4 b får en sammansatt ingrediens uttryckt i total vikt ingå i ingrediensförteckningen under sin egen beteckning, om denna fastställts enligt lag eller sedvana, förutsatt att den omedelbart följs av en uppräkning av de ingredienser som ingår i den sammansatta ingrediensen.
En sådan förteckning skall dock inte vara obligatorisk i följande fall:
a) Om den sammansatta ingrediensen utgör mindre än 25 % av den färdiga varan. Detta undantag skall dock inte gälla i fråga om tillsatser som faller under bestämmelserna i punkt 4 c.
b) Om den sammansatta ingrediensen är ett livsmedel för vilket någon ingrediensförteckning inte krävs enligt gemenskapsregler.
9. Utan hinder av punkt 5 behöver innehållet av vatten inte anges särskilt
a) om vattnet används under framställningsprocessen enbart för att rekonstituera en ingrediens som använts i koncentrerad eller torkad form,
b) om detta utgör en lag som normalt inte konsumeras.
Artikel 7
1. Mängden av en ingrediens eller av en kategori av ingredienser som används vid tillverkningen eller beredningen av ett livsmedel skall anges i enlighet med denna artikel.
2. Den angivelse som avses i punkt 1 skall vara obligatorisk,
a) om den berörda ingrediensen eller kategorin av ingredienser ingår i försäljningsnamnet eller vanligtvis förknippas med det namnet av konsumenterna, eller
b) om den berörda ingrediensen eller kategorin av ingredienser skriftligen, genom en illustration eller grafiskt, framhävs i märkningen, eller
c) om den berörda ingrediensen eller kategorin av ingredienser är nödvändig för att känneteckna livsmedlet och särskilja det från produkter som det skulle kunna förväxlas med på grund av sitt namn och utseende, eller
d) i de fall som fastställs i enlighet med det förfarande som anges i artikel 20.2.
3. Punkt 2 skall inte tillämpas
a) på en ingrediens eller kategori av ingredienser
- vars avrunna nettovikt anges i enlighet med artikel 8.4,
- vars mängd, på grund av gemenskapsbestämmelser, redan måste anges i märknignen,
- som används i små mängder i aromgivande syfte, eller
- som trots att den ingår i försäljningsnamnet inte kommer att styra konsumenternas val i den medlemsstat där saluföringen sker, då variationen i mängd inte är avgörande för att känneteckna livsmedlet eller är sådan att den särskiljer livsmedlet från liknande varor; enligt förfarandet i artikel 20.2 skall det i tveksamma fall avgöras om villkoren i denna strecksats är uppfyllda,
b) om särskilda gemenskapsbestämmelser exakt föreskriver mängden av en ingrediens eller kategori av ingredienser utan att föreskriva att detta skall anges i märkningen,
c) i de fall som avses i artikel 6.5 fjärde och femte strecksatserna,
d) i de fall som fastställs i enlighet med det förfarande som anges i artikel 20.2
4. Den angivna mängden, uttryckt i procent, skall motsvara mängden av ingrediensen eller ingredienserna vid den tidpunkt då de användes. Gemenskapsbestämmelser får emellertid tillåta avvikelser från denna princip för vissa livsmedel. Sådanna bestämmelser skall antas i enlighet med det förfarande som anges i artikel 20.2.
5. Den angivelse som avses i punkt 1 skall antingen ingå i det namn under vilket livsmedlet säljs eller anges omedelbart därintill eller också anges i ingrediensförteckningen i anslutning till ingrediensen eller kategorin av ingredienser i fråga.
6. Denna artikel skall tillämpas utan att det påverkar tilllämpningen av gemenskapens regler om näringsvärdesdeklaration.
Artikel 8
1. Nettoinnehållet i färdigförpackade livsmedel skall anges
- i volymenheter i fråga om vätskor,
- i viktenheter i fråga om andra varor,
varvid liter, centiliter, milliliter, kilogram eller gram skall användas allt efter omständigheterna.
Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser, som gäller för vissa livsmedel, får avvika från denna regel.
Det förfarande som fastställs i artikel 19 skall tillämpas på varje sådan nationell bestämmelse.
2. a) Om gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser innehåller föreskrifter om att ett innehåll skall anges på ett visst sätt (t.ex. nominell kvantitet, minimikvantitet, genomsnittskvantitet) skall denna kvantitet anses som nettoinnehåll enligt detta direktiv.
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemstaterna om varje åtgärd som vidtagits enligt denna punkt.
b) Gemenskapsbestämmelser eller, som sådana saknas, nationella bestämmelser får för vissa livsmedel, som delas in i kategorier efter mängd, innehålla föreskrifter om att mängd skall anges på annat sätt.
Det förfarande som fastställs i artikel 19 skall tillämpas på varje sådan nationell bestämmelse.
c) Om en färdigförpackad vara består av två eller flera separata färdigförpackningar som innehåller samma mängd av samma vara, skall nettoinnehållet anges genom uppgift om nettoinnehållet för varje separat förpackning och det totala antalet sådana förpackningar. Dessa uppgifter är dock inte obligatoriska, om det totala antalet separata förpackningar är klart synligt och lätt kan räknas utifrån, och om minst en uppgift om nettoinnehållet i varje enskild förpackning är klart synlig från utsidan.
d) Om en fördigförpackad vara består av två eller flera separata förpackningar, som vid försäljning inte betraktas som enheter, skall nettoinnehållet anges genom uppgift om det totala nettoinnehållet och det totala antalet separata förpackningar. När det gäller vissa livsmedel behöver gemenskapsbestämmelser, eller om sådana saknas, nationella bestämmelser inte innehålla föreskrifter om att det totala antalet separata förpackningar skall anges.
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24 skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt denna punkt.
3. När det gäller livsmedel som normalt säljs styckevis behöver medlemsstaterna inte kräva uppgift om nettoinnehållet under forutsättning att antalet artiklar är klart synliga och lätt räknas utifrån eller, om detta inte är möjligt, framgår av märkningen.
Utan att det påverkar den anmälningskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt denna punkt.
4. Om ett livsmedel i fast form ligger i en lag, skall även livsmedlets avrunna vikt anges i märkningen.
I denna punkt avses med en "lag" följande varor, eventuellt i blandningar och även i fryst eller djupfryst tillstånd, förutsatt att vätskan bara är ett komplement till den aktuella beredningens viktiga beståndsdelar och således inte en för köpet avgörande faktor: vatten, saltlösningar, saltlake; livsmedelssyror lösta i vatten, ättika; sockerlag, vattenlösningar med andra sötningsmedel; i fråga om frukt eller grönsaker, frukt- eller grönsaksjuicer.
Denna uppräkning kan kompletteras i enlighet med det förfarande som fastställs i artikel 20.2.
Metoder för att kontrollera avrunnen vikt skall bestämmas i enlighet med det förfarande som fastställs i artikel 20.2.
5. Det skall inte vara obligatoriskt att ange nettoinnehållet för livsmedel
a) som minskar avsevärt i volym eller vikt och som säljs styckevis eller vägs i köparens nävraro,
b) vars nettoinnehåll är mindre än 5 g eller 5 ml; dock skall denna bestämmelse inte gälla för kryddor och örter.
Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser som gäller för vissa livsmedel får i undantagsfall fastställa gränsvärden som är högre än 5 g eller 5 ml, under förutsättning att detta inte leder till att köparen får bristfällig information.
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt denna punkt.
6. De gemenskapsbestämmelser som avses i punkterna 1 andra stycket, 2 b, 2 d och 5 andra stycket skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
Artikel 9
1. Datum för minsta hållbarhetstid för ett livsmedel skall vara den dag fram till vilken livsmedlet vid rätt förvaring har kvar sina särskilda egenskaper.
Det skall anges i enlighet med bestämelserna i punkterna 2-5.
2. Datumet skall föregås av orden
- "Bäst före..." när datumet omfattar uppgift om dagen,
- "Bäst före utgången av... " i övriga fall.
3. De ord som anges i punkt 2 skall följas av
- antingen själva datumet, eller
- en hänvisning till var på märkningen datumet finns angivet.
Om det behövs, skall dessa uppgifter följas av de förvaringsanvisningar som man måste rätta sig efter för att varan skall hålla sig under den angivna perioden.
4. Datumet skall bestå av dag, månad och år i okodad kronologisk form.
Dock är det i fråga om livsmedel
- med kortare hållbarhetstid än tre månader tillräckligt att ange dag och månad,
- med längre hållbarhetstid än tre månader men kortare än 18 månader tillräckligt att ange månad och år,
- med längre hållbarhetstid än 18 månader tillräckligt att ange året.
Sättet för att ange datum kan regleras närmare i enlighet med det förfarande som fastställs i artikel 20.2.
5. Om inte annat följer av gemenskapsbestämmelser som fastställer andra typer av datummärkning, skall uppgift om hållbarhetsdatum inte krävas för:
- Färsk frukt och färska grönsaker, inklusive potatis, som inte skalats, delats i bitar eller behandlats på liknande sätt. Detta undantag skall inte tillämpas på groddar och liknande produkter såsom skott av baljväxter.
- Viner, starkviner, mousserande viner, kryddade starkviner och liknande produkter framställda av andra frukter än druvor samt drycker som faller under KN-numren 22060091, 2206 00 93 och 2206 00 99 och som har framställts av druvor eller druvmust.
- Drycker som innerhåller minst 10 volymprocent alkohol.
- Läskedrycker, fruktjuice, fruktnektar och alkoholhaltiga drycker i separata kärl på mer än fem liter och avsedda för storkök.
- Bageri- eller konditorivaror som med hänsyn till sitt innehåll normalt konsumeras inom 24 timmar efter tillverkningen.
- Ättika.
- Koksalt.
- Tuggummi och liknande produkter.
- Portionsförpackningar av glass.
Artikel 10
1. I fråga om livsmedel som från mikrobiologisk synpunkt är lättfördärvliga och som därför efter en kort period kan antas utgära en omedelbar fara för människors hälsa, skall datum för minsta hållbarhetstid ersättas med uppgift om sista förbrukningsdag.
"sista förbrukningsdag".
Orden skall följas av
- antingen själva datumet, eller
- en hänvisning till var på märkningen datumet finns angivet.
Dessa uppgifter skall följas av en beskrivning av de förvaringsanvisningar som man måste rätta sig efter.
3. Datumet skall bestå av dag, månad och eventuellt år i denna ordning och i okodad form.
4. I vissa fall kan det genom det förfarande som fastställs i artikel 20.2 avgöras huruvida villkoren i punkt 1 är uppfyllda.
Artikel 11
1. Bruksanvisningen till ett livsmedel skall vara utformad så att livsmedlet kan användas på ett ändamålsenligt sätt.
2. Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser får i fråga om vissa livsmedel närmare ange hur bruksanvisningarna bör vara utformade.
Det förfarande som fastställs i artikel 19 skall tillämpas på sådana nationella bestämmelser.
De gemenskapsbestämmelser som avses i denna punkt skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
Artikel 12
De bestämmelser som gäller angivande av alkoholhalten uttryckt i volym skall i fråga om varor som faller under tariffrubrikerna nr 22.04 och 22.05 fastställas i särskilda gemenskapsbestämmelser som gäller för dessa varor.
För andra drycker som innehåller mer än 1,2 volymprocent alkohol skall dessa bestämmelser fastställas i enlighet med det förfarande som föreskrivs i artikel 20.2.
Artikel 13
1. a) I fråga om färdigpackade livsmedel skall de uppgifter som anges i artikel 3 och artikel 4.2 finnas på förpackningen eller på en etikett som är fästad vid denna.
b) Utan hinder av punkt a och utan att det påverkar tilllämpningen av gemenskapsbestämmelser om nominella mängder, är det, om färdigförpackade livsmedel är
- avsedda för konsumenter men saluförs i ett handelsled före försäljningen till konsumenten och under förutsättning att försäljning till storkök inte sker i detta handelsled,
c) I de fall som avses i b skall de uppgifter som avses i artikel 3.1.1, 3.1.5 och 3.1.7 och, i tilllämpliga fall, de som avses i artikel 10 också finas på den yttre förpackning, i vilken livsmedlen presenteras när de saluförs.
2. De uppgifter som anges i artikel 3 och artikel 4.2 skall vara lätta att förstå och markeras på väl synlig plats på sådant sätt att de är lätta att se, klart läsbara och outplånliga.
De skall inte på något sätt döljas, skymmas eller avbrytas av annan text eller av någon illustration.
3. De uppgifter som räknas upp i artikel 3.1.1, 3.1.4, 3.1.5 och 3.1.10 skall förekomma i samma synfält.
Detta krav får utvidgas till att omfatta även de uppgifter som avses i artikel 4.2.
4. För regurglas som har märkning som är outplånlig och därför saknar etikett, ring eller krage samt för förpackningar eller kärl med en största yta mindre än 10 cm2, behöver endast de uppgifter anges om avss i artikel 3.1.1, 3.1.4 och 3.1.5.
I detta fall skall punkt 3 inte gälla.
5. Irland, Nederländerna och Förenade kungariket får medge undantag från artikel 3.1 och punkt 3 i denna artikel när det är fråga om mjölk och mjölkprodukter i returglas.
De skall underrätta kommissionen om varje åtgärd som vidtagits i enlighet med punkt 5.
Artikel 14
För livsmedel som saluhålls till konsumenter eller till storkök utan att vara färdigförpackade, eller för livsmedel som förpackas på försäljningsstället på konsumentens begäran eller är färdigförpackade för direkt försäljning, skall medlemsstaterna anta närmare bestämmelser för hur de uppgifter som omfattas av artikel 3 och artikel 4.2 skall anges.
De får besluta att samtliga eller en del av dessa uppgifter inte behöver lämnas, förutsatt att köparen ända får tillfredsställande information.
Artikel 15
Detta direktiv skall inte inverka på bestämmelser i nationell lagstiftning, vilka i avsaknad av gemenskapsbestämmelser innebär mindre stränga krav för märkning av livsmedel som presenteras i presentförpackningar som statyetter eller souvenirer.
Artikel 16
1. Medlemsstaterna skall säkerställa att det inom deras territorier är förbjudet att saluföra livsmedel för vilka uppgifterna enligt artikel 3 och artikel 4.2 inte ges på ett språk som med lätthet förstås av konsumenten, såvida inte konsumenten faktiskt informeras genom andra åtgärder som fastställs i enlighet med det förfarande som anges i artikel 20.2 beträffande en eller flera uppgifter i märkningen.
2. Inom sitt eget territorium får den medlemsstat där saluföringen sker i enlighet med fördragets regler föreskriva att dessa uppgifter i märkningen skall ges på ett eller flera av gemenskapens officiella språk.
3. Bestämmelserna i punkterna 1 och 2 skall inte förhindra att uppgifterna i märkningen ges på flera språk.
Artikel 17
I fråga om reglerna för hur uppgifter i artikel 3 och artikel 4.2 skall anges, skall medlemsstaterna inte fastställa krav som är mer detaljerade än de som framgår av artiklarna 3-13.
Artikel 18
1. Medlemsstater får inte förbjuda handel med livsmedel som följer reglerna i detta direktiv genom att tillämpa nationella icke harmoniserade bestämmelser för märkning och presentation av vissa livsmedel eller av livsmedel i allmänhet.
2. Punkt 1 gäller inte nationella icke harmoniserade bestämmelser som motiveras av att man vill
- skydda människors hälsa,
- förebygga oredlighet, såvida inte sådana bestämmelser kan befaras hindra tillämpningen av de definitioner och regler som fastställs genom detta direktiv,
- skydda industriella och kommersiella äganderätter, uppgifter om ursprung och registrerade ursprungbeteckningar samt att förebygga illojal konkurrens.
Artikel 19
När det hänvisas till denna artikel skall följande förfarande användas, om en medlemsstat skull bedöma det som nödvändigt att anta ny lagstiftning:
Den skall anmäla de planerade åtgärderna och skälen för dessa till kommissionen och de andra medlemsstaterna. Kommissionen skall samråda med medlemsstaterna inom Ständiga livsmedelskommittén, inrättad genom rådets beslut 69/414/EG(6), om den anser att sådant samråd behövs eller om någon medlemsstat begär det.
Medlemsstaterna får vidta åtgärderna tidigast tre månader efter anmälan och under förutsättning att kommissionen inte motsatt sig det.
Om så skulle vara fallet, skall kommissionen före utgången av denna period inleda det förfarande som fastställs i artikel 20.2 för att avgöra huruvida de planerade åtgärdena kan genomföras, om det är nödvändigt med lämpliga ändringar.
Artikel 20
1. Kommissionen skall biträdas av en kommitté (nedan kallad kommittén).
2. När det hänvisas till denna punkt, skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 21
Om det visar sig nödvändigt att vidta tillfälliga åtgärder för att underlätta tillämpningen av detta direktiv, skall de antas i enlighet med det förfarande som fastställs i artikel 20.2
Artikel 22
Detta direktiv skall inte inverka på sådana gemenskapsbestämmelser om märkning och presentation av vissa livsmedel som redan antagits den 22 december 1978.
Varje ändring som är nödvändig för att harmonisera sådana bestämmelser med de regler som fastställs i detta direktiv skall beslutas i enlighet med det förfarande som är tilllämpligt för varje sådan bestämmelse.
Artikel 23
Detta direktiv skall inte gälla varor avsedda för export utanför gemenskapen.
Artikel 24
Medlemsstaterna skall se till att kommissionen får del av texten till alla väsentliga bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 25
Detta direktiv skall gälla också för Frankrikes utomeuropeiska department.
Artikel 26
1. Direktiv 79/112/EEG i dess lydelse enligt direktiven i bilaga IV del A skall upphöra att gälla utan att det påverkar medlemsstaternas förpliktelsre vad gäller de tidsfrister för genomförande som anges i bilaga IV del B.
2. Hänvisningar till det upphävda direktivet skall tolkas som hänvisningar till detta direktiv och skall läsas i enlighet med jämförelsetabellen i bilaga V.
Artikel 27
Kommissionens direktiv 2000/63/EG
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(1) Det är nödvändigt att fastställa renhetskriterier för alla de andra tillsatser än färgämnen och sötningsmedel som anges i Europaparlamentets och rådets direktiv 95/2/EG av den 20 februari 1995 om andra livsmedelstillsatser än färgämnen och sötningsmedel(3), senast ändrat genom direktiv 98/72/EG(4).
(2) I kommissionens direktiv 96/77/EG av den 2 december 1996 om särskilda renhetskriterier för andra livsmedelstillsatser än färgämnen och sötningsmedel(5), ändrat genom direktiv 98/86/EG(6), fastställs renhetskriterier för ett antal livsmedelstillsatser. Detta direktiv bör nu kompletteras med renhetskriterier för de återstående livsmedelstillsatserna i direktiv 95/2/EG.
(3) Med hänsyn till den tekniska utvecklingen är det nödvändigt att ändra de renhetskriterier för butylhydroxianisol (BHA) som anges i direktiv 96/77/EG. Det är därför nödvändigt att anpassa detta direktiv.
(4) Det är nödvändigt att beakta de specifikationer och analysmetoder för tillsatser som anges i den Codex Alimentarius som utarbetats av FAO/WHO:s gemensamma expertkommitté för livsmedelstillsatser (JECFA).
(5) Om livsmedelstillsatser bereds genom produktionsmetoder eller från utgångsmaterial som avsevärt skiljer sig från dem som utvärderats av Vetenskapliga livsmedelskommittén, eller från dem som anges i detta direktiv, bör Vetenskapliga livsmedelskommittén göra en säkerhetsutvärdering av dessa tillsatser, med särskild tonvikt på renhetskriterierna.
(6) De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga livsmedelskommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 96/77/EG ändras på följande sätt:
1) I bilagan skall texten avseende E 320 - butylhydroxianisol (BHA) ersättas med bilaga I till detta direktiv.
2) Bilaga II till detta direktiv skall läggas till i bilagan.
Artikel 2
1) Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 mars 2001. De skall genast underrätta kommissionen om detta.
2) När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
3) Produkter som släpps ut på marknaden eller som märks före den 31 mars 2001 och som inte uppfyller kraven i detta direktiv får saluföras till dess att lagren är tömda.
Artikel 3
Europaparlamentets och rådets direktiv 2000/69/EG
av den 16 november 2000
om gränsvärden för bensen och koloxid i luften
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175.1 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) På grundval av principerna i artikel 174 i fördraget syftar Europeiska gemenskapens program för politik och åtgärder för miljön och en hållbar utveckling (femte miljöhandlingsprogrammet)(4), kompletterat genom Europaparlamentets och rådets beslut nr 2179/98/EG(5) om en översyn av programmet, särskilt till ändringar i lagstiftningen om luftföroreningar. I programmet rekommenderas att det upprättas långsiktiga mål för luftkvaliteten. Enligt artikel 174 i fördraget skall försiktighetsprincipen tillämpas när det gäller skydd av miljön och av människors hälsa.
(2) Enligt artikel 152 i fördraget skall hälsoskyddskraven ingå som ett led i gemenskapens övriga politik. I artikel 3.1 p i fördraget föreskrivs också att gemenskapens verksamhet skall bidra till att uppnå en hög hälsoskyddsnivå.
(3) I enlighet med artikel 4.5 i rådets direktiv 96/62/EG av den 27 september 1996 om utvärdering och säkerställande av luftkvaliteten(6) skall rådet anta de bestämmelser som avses i punkt 1 samt i punkterna 3 och 4 i den artikeln.
(4) Enligt artikel 8 i direktiv 96/62/EG skall det upprättas handlingsplaner för de zoner där koncentrationen av luftförorenande ämnen överskrider gränsvärdena plus tillämpliga tillfälliga toleransmarginaler för att säkerställa att gränsvärdena uppnås inom de fastställda tidsfristerna.
(5) Enligt direktiv 96/62/EG skall numeriska värden för gränsvärdena bygga på resultaten från det arbete som utförs av internationella forskargrupper verksamma inom området. Kommissionen bör ta hänsyn till de senaste rönen från forskning om berörda områden inom epidemiologi och miljö och de senaste framstegen inom metrologin när de faktorer som gränsvärdena bygger på tas upp till förnyad undersökning.
(6) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(7).
(7) Ändringar som är nödvändiga för anpassning till framsteg som görs på det vetenskapliga och tekniska området får endast gälla kriterier och metoder för att bedöma koncentrationerna av bensen och koloxid eller regler för överlämnandet av information till kommissionen och får inte leda till att gränsvärdena direkt eller indirekt ändras.
(8) De gränsvärden som fastställs i detta direktiv är minimikrav. I enlighet med artikel 176 i fördraget får en medlemsstat behålla eller införa strängare skyddsåtgärder. Strängare gränsvärden kan i synnerhet införas för att skydda hälsan hos särskilt sårbara kategorier av befolkningen såsom barn och patienter på sjukhus. En medlemsstat kan kräva att gränsvärdena uppnås före de datum som fastställs i detta direktiv.
(9) Bensen är ett för människor genotoxiskt carcinogen, och det är inte möjligt att fastställa något tröskelvärde under vilket det inte föreligger någon hälsorisk.
(10) När emellertid gränsvärdena för bensen enligt detta direktiv är svåra att uppnå beroende på platsspecifika spridningskarakteristika eller relevanta klimatförhållanden, och om tillämpningen av åtgärderna skulle förorsaka allvarliga socio-ekonomiska problem, kan en medlemsstat be kommissionen om en tidsbegränsad förlängning för en enstaka gång under särskilda förhållanden.
(11) För att underlätta översynen av detta direktiv under år 2004 bör kommissionen och medlemsstaterna överväga att uppmuntra forskning om effekterna av bensen och koloxid. I detta sammanhang bör det förutom till utomhusluft också tas hänsyn till luftföroreningar i inomhusluft.
(12) Standardiserade och tillförlitliga mätmetoder och gemensamma kriterier för placeringen av mätstationer är av stor betydelse för bedömningen av luftkvaliteten om man vill uppnå jämförbara uppgifter över hela gemenskapen.
(13) Information om koncentrationer av bensen och koloxid bör översändas till kommissionen som grundval för regelbundna rapporter.
(14) Aktuella uppgifter om koncentrationer av bensen och koloxid i luften bör finnas lätt tillgängliga för allmänheten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Mål
Syftet med detta direktiv är att
a) fastställa gränsvärden för koncentrationer av bensen och koloxid i luften, så att skadliga effekter på människors hälsa och på miljön i dess helhet kan undvikas, förebyggas eller minskas,
b) utvärdera koncentrationerna av bensen och koloxid i luften på grundval av gemensamma metoder och kriterier,
c) inhämta tillförlitliga uppgifter om koncentrationer av bensen och koloxid i luften, och säkerställa att dessa uppgifter görs tillgängliga för allmänheten,
d) upprätthålla luftkvaliteten, när den är god, och i övriga fall förbättra den med hänsyn till dess halt av bensen och koloxid.
Artikel 2
Definitioner
Definitionerna i artikel 2 i direktiv 96/62/EG skall tillämpas.
I detta direktiv avses med
a) övre utvärderingströskel: den nivå som avses i bilaga III under vilken en kombination av mätningar och modelleringsmetoder kan användas för att utvärdera luftkvaliteten, i enlighet med artikel 6.3 i direktiv 96/62/EG,
b) nedre utvärderingströskel: den nivå som avses i bilaga III under vilken enbart modelleringsmetoder eller objektiva skattningsmetoder kan användas för att utvärdera luftkvaliteten, i enlighet med artikel 6.4 i direktiv 96/62/EG,
c) fasta mätningar: mätningar som utförs i enlighet med artikel 6.5 i direktiv 96/62/EG.
Artikel 3
Bensen
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att koncentrationen av bensen i luften, som utvärderats i enlighet med artikel 5, inte överskrider det gränsvärde som anges i bilaga I med hänsyn till de datum som där anges.
Den toleransmarginal som anges i bilaga I skall tillämpas i enlighet med artikel 8 i direktiv 96/62/EG.
2. När det gränsvärde som anges i bilaga I är svåra att uppnå beroende på platsspecifika spridningskarakteristika eller relevanta klimatförhållanden, t.ex. låg vindhastighet och/eller förhållanden som främjar avdunstning, och om tillämpningen av åtgärderna skulle förorsaka allvarliga socio-ekonomiska problem, kan en medlemsstat be kommissionen om en tidsbegränsad förlängning. Kommissionen kan, i enlighet med det förfarande som anges i artikel 12.2 i direktiv 96/62/EG på begäran av en medlemsstat och utan att det påverkar tillämpningen av artikel 8.3 i detta direktiv, bevilja en enstaka förlängning för en period på upp till fem år om den berörda medlemsstaten
- fastställer de zoner och/eller den tätbebyggelse som berörs,
- tillhandahåller erforderlig motivering för en sådan förlängning,
- visar att alla rimliga åtgärder har vidtagits för att sänka koncentrationerna av de berörda föroreningarna och för att begränsa det område i vilket gränsvärdet överskrids, och
- anger den framtida utvecklingens huvuddrag med avseende på de åtgärder som den kommer att vidta i enlighet med artikel 8.3 i direktiv 96/62/EG.
Det gränsvärde för bensen som tillåts under den tidsbegränsade förlängningen får emellertid inte överskrida 10 μg/m3.
Artikel 4
Koloxid
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att koncentrationen av koloxid i luften, som utvärderats i enlighet med artikel 5, inte överskrider gränsvärdet som anges i bilaga II med hänsyn till de datum som där anges.
Den toleransmarginal som anges i bilaga II skall tillämpas i enlighet med artikel 8 i direktiv 96/62/EG.
Artikel 5
Utvärdering av koncentrationer
1. De övre och nedre utvärderingströsklarna för bensen och koloxid skall vara de tröskelvärden som anges i avsnitt I i bilaga III.
Minst vart femte år skall klassificeringen av varje zon eller tätbebyggelse för de syften som avses i artikel 6 i direktiv 96/62/EG ses över i enlighet med det förfarande som fastställs i avsnitt II i bilaga III till detta direktiv. Klassificeringen skall ses över tidigare om betydande ändringar ägt rum i fråga om verksamhet som påverkar koncentrationerna av bensen eller koloxid i luften.
2. Kriterierna för att bestämma var provtagningsplatserna för mätning av bensen- och koloxid i luften skall placeras är de som anges i bilaga IV. Minsta antalet provtagningsplatser för fasta mätningar av koncentrationer av de berörda föroreningarna fastställs i bilaga V, och de skall installeras i alla zoner eller tätbebyggelser där mätningar krävs om fasta mätningar är den enda källan för uppgifter om koncentrationer i dessa.
3. För zoner och tätbebyggelser där uppgifter från fasta mätstationer kompletteras med uppgifter från andra källor, t.ex. utsläppsinventeringar, indikativa mätmetoder och luftkvalitetsmodellering, skall antalet fasta mätstationer som skall upprättas och den rumsliga upplösningen för övriga metoder vara tillräckliga för att göra det möjligt att fastställa koncentrationerna av luftföroreningar i enlighet med avsnitt I i bilaga IV och avsnitt I i bilaga VI.
4. För zoner och tätbebyggelser där inga mätningar krävs får modelleringsmetoder eller objektiva skattningsmetoder tillämpas.
5. Referensmetoderna för analys och provtagning av bensen och koloxid anges i avsnitten I och II i bilaga VII. I avsnitt III i bilaga VII kommer referensmetoder för luftkvalitetsmodellering att anges när sådana tekniker finns tillgängliga.
6. Medlemsstaterna skall underrätta kommissionen om de metoder som används för den preliminära utvärderingen av luftkvaliteten enligt artikel 11.1 d i direktiv 96/62/EG senast den dag som anges i artikel 10 i detta direktiv.
7. De ändringar som behövs för att anpassa bestämmelserna i denna artikel samt i bilagorna III-VII till den vetenskapliga och tekniska utvecklingen skall antas i enlighet med det förfarande som avses i artikel 6.2, men de får inte leda till direkta eller indirekta ändringar av gränsvärdena.
Artikel 6
Kommitté
1. Kommissionen skall biträdas av den kommitté som avses i artikel 12.2 i direktiv 96/62/EG, nedan kallad kommittén.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 7
Information till allmänheten
1. Medlemsstaterna skall se till att aktuell information om koncentrationerna av bensen och koloxid i luften rutinmässigt görs tillgänglig för allmänheten, liksom för berörda organisationer, såsom miljöorganisationer, konsumentorganisationer, organisationer som företräder känsliga befolkningsgruppers intressen och andra berörda hälso- och sjukvårdsorgan, till exempel via radio och TV, tidningar, informationstavlor och datanättjänster, teletext, telefon eller fax.
Informationen om koncentrationerna av bensen i luften skall, i form av ett genomsnittsvärde för de tolv senaste månaderna, uppdateras minst var tredje månad och, där det är praktiskt genomförbart, en gång i månaden. Information om koncentrationerna av koloxid i luften skall, i form av ett högsta genomsnittsvärde för åtta timmar i följd, uppdateras minst en gång per dag och där det är praktiskt genomförbart en gång per timme.
Den information som avses i andra stycket skall åtminstone innehålla uppgifter om överskridanden av gränsvärdena för koncentrationerna under de genomsnittsperioder som anges i bilagorna I och II. Den skall även omfatta en kort utvärdering med avseende på gränsvärdena och relevant information om hälsoeffekter.
2. När medlemsstaterna gör planer och program i enlighet med bestämmelserna i artikel 8.3 i direktiv 96/62/EG tillgängliga för allmänheten skall de också göra dem tillgängliga för de organisationer som avses i punkt 1 i denna artikel. Detta gäller också den dokumentation som erfordras enligt bilaga VI.II.
3. Information till allmänheten och organisationer i enlighet med punkterna 1 och 2 skall vara tydlig, begriplig och lättillgänglig.
Artikel 8
Rapport och översyn
1. Senast den 31 december 2004 skall kommissionen till Europaparlamentet och rådet överlämna en rapport som är grundad på de erfarenheter som gjorts vid tillämpningen av detta direktiv, och särskilt på resultaten av den senaste vetenskapliga forskningen om effekterna på människors hälsa, varvid särskild hänsyn skall tas till känsliga befolkningsgrupper, och på ekosystemen av exponering för bensen och koloxid, samt på den tekniska utvecklingen, inbegripet framsteg i fråga om mätmetoder och andra sätt att utvärdera bensen- och koloxidkoncentrationer i luften.
2. Den rapport som avses i punkt 1 skall när det gäller bensen och koloxid särskilt ta hänsyn till följande:
a) Den nuvarande luftkvaliteten och tendenserna fram till år 2010 och därefter.
b) Möjligheterna till ytterligare minskningar av förorenande utsläpp från alla relevanta källor, med beaktande av teknisk genomförbarhet och kostnadseffektivitet.
c) Förhållandet mellan föroreningar och möjligheter till kombinerade strategier för att uppnå gemenskapens mål i fråga om luftkvalitet och liknande mål.
d) Nuvarande och framtida krav i fråga om information till allmänheten och utbyte av information mellan medlemsstater och kommissionen.
e) De erfarenheter som gjorts i medlemsstaterna vid tillämpningen av detta direktiv, i synnerhet de förhållanden, enligt föreskrifterna i bilaga IV, under vilka mätningarna utförts.
3. För att upprätthålla en hög skyddsnivå för människors hälsa och för miljön skall rapporten som avses i punkt 1 vid behov kompletteras med förslag till ändringar av detta direktiv som kan inbegripa ytterligare förlängningar av tidsfristen för att uppnå gränsvärdet för bensen enligt bilaga I vilka kan komma att beviljas i enlighet med artikel 3.2.
Artikel 9
Påföljder
Medlemsstaterna skall besluta om de påföljder som skall tillämpas vid överträdelser av de nationella bestämmelser som antas i enlighet med detta direktiv. Dessa påföljder skall vara effektiva, proportionella och avskräckande.
Artikel 10
Genomförande
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 13 december 2002. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 11
Ikraftträdande
Kommissionens förordning (EG) nr 645/2000
av den 28 mars 2000
om fastställande av de tillämpningsföreskrifter som krävs för ett korrekt bruk av vissa bestämmelser i artikel 7 i rådets direktiv 86/362/EEG och artikel 4 i rådets direktiv 90/642/EEG om arrangemang för övervakning av gränsvärdena för bekämpningsmedelsrester i och på spannmål och produkter av vegetabiliskt ursprung inklusive frukt och grönsaker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 86/362/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på spannmål(1), senast ändrat genom kommissionens direktiv 1999/71/EG(2), särskilt artikel 7 i detta,
med beaktande av rådets direktiv 90/642/EEG av den 27 november 1990 om fastställande av gränsvärden för bekämpningsmedelsrester i och på produkter av vegetabiliskt ursprung inklusive frukt och grönsaker(3), senast ändrat genom direktiv 1999/71/EG, särskilt artikel 4 i detta, och
av följande skäl:
(1) I artikel 7 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG fastställs grundläggande bestämmelser för kontroll av bekämpningsmedelsrester i och på spannmål respektive frukt och grönsaker.
(2) Erfarenheterna från utformning och tillämpning av kommissionens rekommendationer har visat att flerårig planering, med möjlighet till årliga justeringar, torde vara det effektivaste sättet att upprätta Europeiska gemenskapens samordnade kontrollprogram.
(3) I artikel 7 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG föreskrivs det att nödvändiga bestämmelser skall ses över och antas, till exempel om offentliggörande i rapporter från Europeiska gemenskapen av sammanställningar av kontrollen i medlemsstaterna, och att det skall beslutas om åtgärder på gemenskapsnivån vid rapporterade överträdelser av gränsvärdena. Erfarenheterna har bekräftat att de laboratorier som gör analyser med avseende på bekämpningsmedelsrester måste uppfylla höga kvalitetskrav för att deras resultat skall vara tillförlitliga. Laboratoriernas deltagande i regelbundna kvalifikationsprövningar och tillämpning av gemensamnaa riktlinjer för kvalitetskontroll kan användas för att verifiera att de uppfyller ackrediteringskraven enligt artikel 3 i rådets direktiv 93/99/EEG av den 29 oktober 1993(4) om ytterligare åtgärder för offentlig kontroll av livsmedel.
(4) Eftersom kommissionen vid sammanställning av de uppgifter som lämnas av medlemsstaterna som underlag till de rapporter Europeiska gemenskapen skall offentliggöra måste kunna lita på uppgifternas kvalitet, noggrannhet och jämförbarhet bör kommissionen bidra ekonomiskt till åtgärder som medverkar till att kontrollprogrammen uppfyller högsta möjliga kvalitetskrav. Särskilt de regelbundna kvalifikationsprövningarna samt översynen och utformningen av riktlinjer för kvalitetskontroll i samband med regelbundna expertmöten bör stödjas.
(5) Kommissionen bör bidra ekonomiskt till åtgärder som stärker andra aspekter av samarbetet beträffande kontroll av bekämpningsmedelsrester på gemenskapsnivå. Särskilt bör sådan verksamhet stödjas som på sikt främjar utvecklingen av ett system på gemenskapsnivå som gör det möjligt att på grundval av data från kontrollprogrammen beräkna det dagliga intaget av bekämpningsmedelsrester via kosten.
(6) I kommissionens meddelande KOM(97) 183 om konsumenters hälsa och livsmedelssäkerhet beskrivs kontroll- och inspektionsverksamheten på livsmedels-, veterinär- och växtskyddsområdet. Denna bör innefatta kontrollen med avseende på bekämpningsmedelsrester i och på spannmål, frukt och grönsaker.
(7) Vid de kontroller som genomfördes 1996 och 1997 påvisades överträdelser av de gränsvärden som fastställs i direktiv 90/642/EEG i dess ändrade form.
(8) Både i direktiv 90/642/EEG i dess ändrade form och i direktiv 86/362/EEG i dess ändrade form ges förutsättningar för att det skall kunna vidtas åtgärder på gemenskapsnivå vid rapporterade överträdelser och att de tillämpningsföreskrifter skall antas som krävs för att kontrollen skall fungera väl.
(9) En sammanfattande översikt av kontrollsystemen i alla medlemsstater krävs för att förbättra kontrollen av bekämpningsmedelsrester i gemenskapen och medverka till att den fungerar på avsett sätt.
(10) De tillämpningsföreskrifter bör fastställas som krävs för ett korrekt bruk av kontrollbestämmelserna. I dessa föreskrifter bör det tydligt anges vilka åtgärder och förfaranden kommissionen får stödja ekonomiskt inom ramen för tillgängliga budgetanslag.
(11) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för växtskydd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Kommissionens rekommendationer enligt bestämmelserna i artikel 7.2 b i direktiv 86/362/EEG och artikel 4.2 b i direktiv 90/642/EEG får omfatta perioder på mellan ett och fem år.
2. För att fleråriga kontrollprogram skall kunna administreras effektivt får kommissionen lämna årliga bekräftelser och kompletteringar till förslag till rekommendationer. Dessa skall, i enlighet med artikel 7.2 b i direktiv 86/362/EEG och artikel 4.2 b i direktiv 90/642/EEG, överlämnas till Ständiga kommittén för växtskydd.
Artikel 2
Kommissionen skall underlätta tillämpningen av bestämmelserna i artikel 7.2 och 7.3 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG på följande sätt:
1. Samordna medlemsstaternas verksamhet beträffande kraven för att skapa, registrera, hantera och överföra information om kontroll och kontrollprogram, i tillämpliga fall med hjälp av riktlinjer från Ständiga kommittén för växtskydd, särskilt riktlinjerna för kvalitetskontrollförfaranden vid analys av bekämpningsmedelsrester(5) och vägledningsdokumentet till medlemsstaterna om kommissionens rekommendation om gemenskapens samordnade kontrollprogram(6).
2. Inom ramen för de tillgängliga budgetanslagen i Europeiska gemenskapens budget ge ekonomiskt stöd till
a) regelbundet anordnade kvalifikationsprövningar, i princip vartannat år, av alla laboratorier som utför analyser, i syfte att säkerställa kvalitet, noggrannhet och jämförbarhet av de uppgifter som medlemsstaterna lämnar till kommissionen och övriga medlemsstater årligen och som insamlas och sammanställs av kommissionen för offentliggörande i enlighet med artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG,
b) utveckling av kvalitetskontrollförfaranden för analys av bekämpningsmedelsrester, i form av anvisningar från Ständiga kommittén för växtskydd, och till regelbunden översyn på expertmöten, i princip vartannat år, av tillämpningen av sådana förfaranden på de laboratorier i medlemsstaterna som utför analyser med avseende på bekämpningsmedelsrester, i syfte att säkerställa kvalitet, noggrannhet och jämförbarhet av de uppgifter som medlemsstaterna lämnar till kommissionen och övriga medlemsstater årligen och som insamlas och sammanställs av kommissionen för offentliggörande i enlighet med artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG,
c) till årlig organisation av undersökningar, samråd och andra förberedelser som krävs för att kommissionen skall kunna arbeta i riktning mot ett system som gör det möjligt att på grundval av uppgifter från kontrollprogrammen beräkna det faktiska intaget av bekämpningsmedelsrester via kosten, i enlighet med andra stycket i artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG, och
d) till organisation av andra åtgärder på gemenskapsnivå, definierade av kommissionen och Ständiga kommittén för växtskydd, som krävs för en korrekt tillämpning av artikel 7.2 och 7.3 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG.
Artikel 3
1. Kommissionen skall genom ett beslut som fattas enligt förfarandena i artikel 12 i direktiv 86/362/EEG och artikel 10 i direktiv 90/642/EEG utse den eller de mottagare av ekonomiskt stöd som avses i artikel 2.2.
2. I det kommissionsbeslut som avses i punkt 1 skall särskilt anges
- namnet på mottagaren eller mottagarna av det ekonomiska stödet från gemenskapen,
- den totala kostnaden för den åtgärd som skall genomföras och åtagandena från de parter som deltar i genomförandet, inbegripet Europeiska gemenskapen,
- en sammanfattande beskrivning av åtgärden,
- en tidsplan för slutförandet av åtgärden.
Artikel 4
Medlemsstaterna skall säkerställa att de analysresultat som årligen översänds till kommissionen och till övriga medlemsstater i enlighet med bestämmelserna i artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG har erhållits från laboratorier som
- uppfyller kraven i artikel 3 i direktiv 93/99/EEG och
- på alla sätt har strävat efter att tillämpa de kvalitetskontroll-förfaranden för analys av bekämpningsmedelsrester som avses i artikel 2.2 b i denna förordning.
Medlemsstaterna skall dessutom säkerställa att endast laboratorier som har deltagit i en tidigare eller skall delta i nästa omgång av gemenskapens relevanta kvalifikationsprövningar enligt artikel 2.2 a i denna förordning deltar i gemenskapens samordnade program.
Artikel 5
1. Kommissionen skall utse särskilda tjänstemän med lämpliga kvalifikationer för att i medlemsstaterna tillsammans med nationella myndigheter följa genomförandet av nationella respektive gemenskapens kontrollprogram för bekämpningsmedelsrester i och på livsmedel av vegetabiliskt ursprung. Detta inbegriper provtagning och kvaliteten på relevanta laboratoriers arbete.
2. Tjänstemännen skall besöka de nationella myndigheterna i varje medlemsstat, som skall samarbeta med kommissionens utsedda tjänstemän och ge dem all nödvändig assistans i deras arbete. Besöksprogrammen skall organiseras och genomföras i samarbete med den berörda medlemsstaten. De nationella myndigheterna skall under alla omständigheter fortsätta att ansvara för att kontrollåtgärderna genomförs.
3. Kommissionen skall avtala om dessa besök med nationella tjänstemän inom en lämplig tidsrymd. Förutom experter från den medlemsstat som besöks får kommissionens experter vid kontrollbesöken åtföljas av en eller flera experter från en eller flera av de övriga medlemsstaterna. Under besöken skall experten eller experterna som utsetts av kommissionen från någon medlemsstat följa kommissionens administrativa föreskrifter.
4. Efter varje besök skall kommissionen sammanställa en skriftlig rapport. Den besökta medlemsstaten skall ges möjlighet att lämna synpunkter på rapporten.
5. Kommissionen skall regelbundet genom skriftliga rapporter inom Ständiga kommittén för växtskydd underrätta alla medlemsstater om resultatet av kontrollbesöken i varje medlemsstat. Kommissionen skall underrätta Europaparlamentet. Kommissionen skall också regelbundet offentliggöra rapporterna.
6. Bestämmelserna i denna artikel skall ses över senast den 31 oktober 2001.
Artikel 6
Denna förordning träder i kraft den 1 april 2000.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets förordning (EG) nr 657/2000
av den 27 mars 2000
om förstärkt dialog med fiskerisektorn och de grupper som berörs av den gemensamma fiskeripolitiken
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande, och
(2) Mot bakgrund av uppdragen för den rådgivande kommittén för fiske och vattenbruk (nedan kallad den rådgivande kommittén), vilken förnyades genom kommissionens beslut 1999/478/EG(1), kan målen dialog och öppenhet främjas genom nya åtgärder, som syftar dels till att bättre organisera den rådgivande kommitténs möten, dels till att sprida information till de berörda grupperna om insatser och resultat.
(3) De europeiska branschorganisationerna bör därför få hjälp med att förbereda den rådgivande kommitténs möten i syfte att främja analyser av alla insatser inom den gemensamma fiskeripolitiken och av effekten av dess åtgärder, att stödja olika initiativ från sektorn och att om möjligt söka finna gemensamma ståndpunkter beträffande kommissionens utkast till förslag.
(4) För att förbättra villkoren för beslutsfattandet bör också sektorn mycket tidigt informeras om planerade initiativ, och samtliga berörda grupper bör få förklaringar till olika åtgärders syften och förutsättningar inom ramen för den gemensamma fiskeripolitiken.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Kommissionen skall, enligt de villkor som föreskrivs i bilagan, svara för utgifter avseende
- de europeiska branschorganisationernas möten för att förbereda mötena i den rådgivande kommittén,
- förklaring av syften och åtgärder som avser den gemensamma fiskeripolitiken, särskilt förslag från kommissionen, och spridande av relevant information på detta område till fiskerisektorn och andra berörda grupper under upprätthållande av regelbundna kontakter med de berörda organisationerna och grupperna.
Även expertmöten som kommissionen organiserar för att stödja insatser som omfattas av första stycket, andra strecksatsen, kan finansieras.
Artikel 2
Kommissionen kan göra de kontroller den finner vara nödvändiga för att säkerställa efterlevnaden av villkoren för och fullgörandet av de uppgifter som denna förordning ger de europeiska branschorganisationerna, vilka bistår de ombud som kommissionen utser för detta ändamål.
Artikel 3
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Rådets förordning (EG) nr 813/2000
av den 17 april 2000
om komplettering av bilagan till kommissionens förordning (EG) nr 1107/96 om registrering av geografiska beteckningar och ursprungsbeteckningar enligt förfarandet i artikel 17 i förordning (EEG) nr 2081/92
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av kommissionens förslag,
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel(1), särskilt artikel 17.2 i denna, och
av följande skäl:
(1) För vissa beteckningar som medlemsstaterna har meddelat i enlighet med artikel 17 i förordning (EEG) nr 2081/92 har det begärts kompletterande uppgifter för att säkerställa att dessa beteckningar uppfyller kraven i artiklarna 2 och 4 i nämnda förordning. Efter granskning av dessa kompletterande uppgifter har det visat sig att dessa beteckningar stämmer överens med nämnda artiklar. De bör därför registreras och läggas till i bilagan till kommissionens förordning (EG) nr 1107/96(2).
(2) Den i artikel 15 i förordning (EEG) nr 2081/92 angivna kommittén har inte avgivit ett positivt yttrande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till kommissionens förordning (EG) nr 1107/96 skall kompletteras med beteckningarna i bilagan till denna förordning.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1685/2000
av den 28 juli 2000
om närmare bestämmelser för genomförandet av rådets förordning (EG) nr 1260/1999 avseende stödberättigande utgifter i samband med insatser som medfinansieras av strukturfonderna
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1260/1999 av den 21 juni 1999 om allmänna bestämmelser för strukturfonderna(1), särskilt artikel 30.3 och artikel 53.2 i denna,
efter att samråd har skett med den kommitté som avses i artikel 147 i fördraget, Kommittén för jordbruksstruktur och landsbygdsutveckling och Kommittén för fiskets och vattenbrukets struktur, och
av följande skäl:
(1) I artikel 1.3 i rådets förordning (EG) nr 1257/1999 av den 17 maj 1999 om stöd från Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) till utveckling av landsbygden och om ändring och upphävande av vissa förordningar(2) anges att åtgärder för utveckling av landsbygden som är integrerade med åtgärder som främjar utvecklingen och den strukturella anpassningen i regioner vars utveckling släpar efter (mål 1) eller som åtföljer åtgärder till stöd för ekonomisk och social omställning i områden med strukturella svårigheter (mål 2) i de berörda områdena, skall beakta strukturfondernas särskilda syften med gemenskapens stöd i enlighet med villkoren i förordning (EG) nr 1260/1999. I artikel 2 i förordning (EG) nr 1257/1999 anges vilka typer av åtgärder som kan komma i fråga för stöd till utveckling av landsbygden.
(2) I artikel 2 i Europaparlamentets och rådets förordning (EG) nr 1783/1999 av den 12 juli 1999 om Europeiska regionala utvecklingsfonden(3) anges vilken typ av åtgärder som ERUF kan delta i finansieringen av.
(3) I artikel 3 i Europaparlamentet och rådets förordning (EG) nr 1784/1999 av den 12 juli 1999 om Europeiska socialfonden(4) anges vilken typ av åtgärder som ESF kan stödja.
(4) I artikel 2 i rådets förordning (EG) nr 1263/1999 av den 21 juni 1999 om Fonden för fiskets utveckling(5) anges vilken typ av åtgärder som kan genomföras med finansiellt stöd från FFU. I rådets förordning (EG) nr 2792/1999(6) fastställs närmare föreskrifter och villkor för strukturåtgärderna inom fiskerisektorn.
(5) Enligt artikel 30.3 i förordning (EG) nr 1260/1999 skall nationella regler för stödberättigande utgifter tillämpas om inte kommissionen anser det nödvändigt att anta regler på gemenskapsnivå. För vissa typer av insatser eller projekt anser kommissionen att det är nödvändigt att anta gemensamma regler om stödberättigande utgifter så att en enhetlig och rättvis tillämpning av strukturfonderna kan garanteras över hela gemenskapen. När en regel om någon särskild typ av verksamhet antas, föregriper detta inte frågan enligt vilken av de ovan nämnda fonderna medfinansieringen kan ske. Antagandet av dessa regler bör i vissa fall som bör anges, inte hindra medlemsstaterna från att tillämpa strängare nationella bestämmelser. Reglerna bör vara tillämpliga på alla utgifter som uppstått mellan de tidpunkter som anges i artikel 30.2 i förordning (EG) nr 1260/1999.
(6) Enligt artikel 36.1 i förordning (EG) nr 1257/1999 skall förordning (EG) nr 1260/1999 och de bestämmelser som antagits för genomförandet av den förordningen, om inte något annat följer av förordning (EG) nr 1257/1999, tillämpas på landsbygdsutvecklingsåtgärder i områden som omfattas av mål 2 som finansieras av garantisektionen inom EUGFJ. Reglerna i den här förordningen skall därför tillämpas på sådana åtgärder som omfattas av programmen för de regioner som omfattas av mål 2, såvida inte något annat följer av förordning (EG) nr 1257/1999 och kommissionens förordning (EG) nr 1750/1999(7) om tillämpningsföreskrifter till förordning (EG) nr 1257/1999.
(7) Artiklarna 87 och 88 i fördraget är tillämpliga på verksamhet som medfinansieras av strukturfonderna. Ett kommissionsbeslut om att godkänna en stödform innebär inte någon förhandsbedömning av statsstödsreglerna och befriar inte medlemsstaten från sina skyldigheter enligt dessa artiklar.
(8) De åtgärder som föreskrivs i den här förordningen är förenliga med yttrandet från Kommittén för utveckling och omställning av regioner.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Reglerna i bilagan till den här förordningen skall tillämpas vid bestämmandet av om utgifter kan anses stödberättigande enligt de stödformer som definieras i artikel 9 e i förordning (EG) nr 1260/1999.
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets förordning (EG) nr 2038/2000
av den 28 september 2000
om ändring av förordning (EG) nr 2037/2000 om ämnen som bryter ned ozonskiktet vad gäller dosaerosoler och läkemedelspumpar
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175.1 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(1),
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(2), och
av följande skäl:
(1) Enligt Europaparlamentets och rådets förordning (EG) nr 2037/2000 av den 29 juni 2000 om ämnen som bryter ned ozonskiktet(3) är export av dosaerosoler till utvecklingsländer och export av läkemedelspumpar som innehåller klorfluorkarboner förbjuden. Exporten av dessa hälsovårdsprodukter som får användas på gemenskapens marknad bör dock inte begränsas.
(2) Förordning (EG) nr 2037/2000 bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande punkt skall läggas till i artikel 11.1 i förordning (EG) nr 2037/2000:
"f) dosaerosoler som innehåller klorfluorkarboner och doseringsmekanismer som innehåller klorfluorkarboner för hermetiskt tillslutna apparater avsedda att implanteras i människokroppen för att avge uppmätta läkemedelsdoser, vilka enligt artikel 4.1 kan erhålla ett tillfälligt undantag enligt det förfarande som avses i artikel 18.2."
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Rådets förordning (EG) nr 2578/2000
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3759/92 av den 17 december 1992 om den gemensamma organisationen av marknaden för fiskeri- och vattenbruksprodukter(1), särskilt artikel 2.3 i denna,
med beaktande av kommissionens förslag, och
(2) Därför bör gemensamma och harmoniserade handelsnormer fastställas för hela gemenskapsmarknaden för dessa arter genom ändring av rådets förordning (EG) nr 2406/96(3).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 2406/96 ändras på följande sätt:
1. I artikel 3 skall
a) följande strecksatser läggas till listan i punkt 1 a:
"- Mulle (Mullus barbatus, Mullus surmuletus)
- Havsruda (Spondyliosoma cantharus) och"
b) följande punkt införas i punkt 1:
"d) Stor kammussla och andra ryggradslösa vattendjur enligt KN-nummer 0307:
- Stor kammussla (Pecten maximus)
- Vanlig valthornssnäcka (Buccinum undatum)".
2. Artikel 4.3 första stycket skall ersättas med följande text:"3. Krabba, stor kammussla och vanlig valthornssnäcka enligt artikel 3 skall inte klassificeras enligt särskilda färskhetsnormer."
3. Artikel 7.1 skall ersättas med följande text:
"1. Produkter enligt artikel 3 skall bedömas efter vikt eller antal per kilo. Hästräkor och krabbor skall dock delas in i storlekskategorier på grundval av skalets omfång. Stora kammusslor och vanliga valthornssnäckor skall delas in i storlekskategorier på grundval av snäckans omfång."
4. I bilaga II skall tabellen i bilagan till den här förordningen avseende de storlekskategorier för mulle, havsruda, stor kammussla och vanlig valthornssnäcka införas efter befintlig tabell.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets förordning (EG) nr 2700/2000
av den 16 november 2000
om ändring av rådets förordning (EEG) nr 2913/92 om inrättandet av en tullkodex för gemenskapen
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 26, 95 och 133 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) I rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(4) anges det i artikel 253.4 att rådet före den 1 januari 1998 på grundval av en rapport från kommissionen, som kan åtföljas av eventuella förslag, skall se över tullkodexen för att göra nödvändiga anpassningar, med särskild hänsyn till genomförandet av den inre marknaden.
(2) Varje översyn av kodexen bör, utan att det införs några hinder för den internationella handeln, utgöra ett tillfälle att inrätta instrument och förfaranden som gör det möjligt att förebygga bedrägeri, med tanke på att förebyggande av bedrägeri är ett av de bästa sätten att skydda skattebetalarnas pengar enligt rådets slutsatser av den 19 maj 1998.
(3) Hänsyn bör tas till rådets resolution av den 25 oktober 1996 om förenkling och rationalisering av gemenskapens tullföreskrifter och tullförfaranden(5).
(4) De olika myndigheternas befogenheter att fastställa växelkurser efter införandet av euron har ännu inte fastställts.
(5) Det bör föreskrivas att en tulldeklaration som har upprättats med databehandlingsteknik inte behöver åtföljas av vissa dokument.
(6) Förfarandena för aktiv förädling, bearbetning under tullkontroll och temporär import bör göras lättare att använda genom att reglerna på området görs flexiblare.
(7) Det bör i enlighet med kommittéförfarandet fastställas ytterligare fall där taxeringen inom ramen för förfarandet för passiv förädling beräknas på grundval av kostnaderna för processen.
(8) Det kan vara lämpligt att i vissa frizoner tillåta att tullformaliteter fullgörs och myndigheternas tullkontroller utförs i enlighet med tullagerförfarandet.
(9) Under vissa omständigheter bör gynnsam behandling i tullhänseende med anledning av varors beskaffenhet eller deras användning för särskilda ändamål samt differenstaxering inom ramen för förfarandet för passiv förädling även tillämpas när en tullskuld har uppkommit av andra skäl än övergång till fri omsättning.
(10) I bestämmelserna om platsen för en tullskulds uppkomst bör särskilda regler införas för de fall där beloppet i fråga understiger en viss nivå.
(11) Det är, när det gäller förmånsbehandling, nödvändigt att definiera vad som avses med begreppen misstag som begåtts av tullmyndigheter och god tro hos gäldenären. Gäldenären bör inte bära ansvaret för att systemet fungerar dåligt på grund av ett misstag som har begåtts av myndigheter i tredje land. Sådana myndigheters utfärdande av ett oriktigt ursprungsintyg bör emellertid inte anses som ett misstag om ursprungsintyget har utfärdats på grundval av en ansökan som innehåller oriktiga uppgifter. Oriktigheten i de uppgifter som exportören lämnat i sin ansökan bör bedömas på grundval av alla de faktiska förhållanden som ansökningen innehåller. En gäldenär kan åberopa god tro när han kan visa att han handlat med tillbörlig aktsamhet, utom då ett yttrande om att det finns välgrundade tvivel har offentliggjorts i Europeiska gemenskapernas officiella tidning.
(12) Gemenskapens ekonomiska intressen och gäldenärens rättigheter bör skyddas mot alltför utdragna rättsliga förfaranden.
(13) I de fall där skulden har uppkommit på grund av att en vara har undandragits från tullkontroll och där det finns fler än en gäldenär bör uppskov med betalningen av tullskulden kunna beviljas för att göra det möjligt för tullmyndigheterna att inleda ett uppbördsförfarande gentemot en bestämd gäldenär före de andra gäldenärerna.
(14) De åtgärder som krävs för att genomföra förordning (EEG) nr 2913/92 bör fastställas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(6).
(15) Förordning (EEG) nr 2913/92 bör ändras i enlighet härmed.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 2913/92 ändras på följande sätt:
1. I artikel 4 skall punkt 24 ersättas med följande:
"24. kommittéförfarande: det förfarande som avses dels i artiklarna 247 och 247a, dels i artiklarna 248 och 248a."
2. I artikel 35 skall första stycket ersättas med följande:"Om faktorer som används för att fastställa tullvärdet på varor uttrycks i en annan valuta än den som används i den medlemsstat där värderingen görs, skall den växelkurs tillämpas som vederbörligen har offentliggjorts av de på detta område behöriga myndigheterna."
3. I artikel 77 skall den nuvarande texten betecknas punkt 1 och följande punkt skall läggas till:
"2. För tulldeklarationer som upprättas med hjälp av databehandlingsteknik får tullmyndigheterna tillåta att de åtföljande dokument som avses i artikel 62.2 inte bifogas deklarationen. I detta fall skall dokumenten hållas tillgängliga för tullmyndigheterna."
4. I artikel 115 skall punkt 4 ersättas med följande:
"4. Åtgärder avsedda att förbjuda tillämpningen av punkt 1, att underställa tillämpningen vissa villkor eller att underlätta tillämpningen kan antas enligt kommittéförfarandet."
5. I artikel 117 c skall följande mening läggas till:"De fall där de ekonomiska villkoren skall anses vara uppfyllda får fastställas enligt kommittéförfarandet."
6. Artikel 124 skall ersättas med följande:
"Artikel 124
1. Restitutionssystemet får användas för alla varor. Det får dock inte användas i de fall där, vid tidpunkten för mottagandet av deklarationen om övergång till fri omsättning
- importvarorna omfattas av kvantitativa importrestriktioner,
- importvarorna omfattas av en tullförmån inom ramen för kvotsystemet,
- importvarorna omfattas av krav på att import- eller exportintyg skall uppvisas enligt den gemensamma jordbrukspolitiken, eller
- ett exportbidrag eller en exportavgift har fastställts för förädlingsprodukterna.
2. Dessutom kan ingen återbetalning av importtullar enligt restitutionssystemet ske om förädlingsprodukterna vid mottagandet av deklarationen om export omfattas av krav på uppvisande av import- eller exportintyg enligt den gemensamma jordbrukspolitiken eller om det har fastställts ett exportbidrag eller en exportavgift för dessa produkter.
3. Undantag från bestämmelserna i punkterna 1 och 2 får fastställas enligt kommittéförfarandet."
7. Artikel 131 skall ersättas med följande:
"Artikel 131
De fall i vilka förfarandet för bearbetning under tullkontroll får användas och de särskilda villkoren för användningen skall fastställas enligt kommittéförfarandet."
8. I artikel 133 e skall följande mening läggas till:"De fall där de ekonomiska villkoren skall anses vara uppfyllda får fastställas enligt kommittéförfarandet."
9. Artikel 142 skall ersättas med följande:
"Artikel 142
1. Tillämpning av förfarandet för temporär import med partiell befrielse från importtullar skall beviljas för varor som inte omfattas av de bestämmelser som fastställts enligt artikel 141 eller som omfattas av dessa bestämmelser, men inte uppfyller alla de villkor som anges i dem för beviljande av temporär import med fullständig befrielse.
2. Listan på de varor för vilka förfarandet för temporär import med partiell befrielse från importtullar inte får användas, samt de villkor under vilka förfarandet får användas, skall fastställas enligt kommittéförfarandet."
10. I artikel 153 skall följande stycke läggas till:"Utan hinder av artikel 151 får det enligt kommittéförfarandet fastställas i vilka fall och på vilka särskilda villkor som det vid övergång till fri omsättning av varor efter passiv förädling kan medges att kostnaden för förädlingsprocessen används som grund för taxeringen vid tillämpningen av Europeiska gemenskapernas tulltaxa."
11. I artikel 167 skall punkt 3 ersättas med följande:
"3. Med undantag för de frizoner som utses i enlighet med artikel 168a skall frizonerna vara inhägnade. Medlemsstaterna skall fastställa infarts- och utfartsplatserna för varje frizon eller frilager."
12. I artikel 168 skall punkt 1 ersättas med följande:
"1. Med undantag för de frizoner som utses i enlighet med artikel 168a skall frizonernas och frilagrens gränser samt deras infarter och utfarter övervakas av tullmyndigheterna."
13. Följande artikel skall införas mellan artikel 168 och punkt B (Uppläggning av varor i frizoner eller frilager):
"Artikel 168a
1. Tullmyndigheterna får utse frizoner inom vilka tullkontroller och tullformaliteter skall utföras i enlighet med tullagerförfarandet och inom vilka bestämmelserna om tullskuld skall tillämpas i enlighet med tullagerförfarandet.
Artiklarna 170, 176 och 180 skall inte tillämpas på de frizoner som utsetts på detta vis.
2. De frizoner som avses i artiklarna 37, 38 och 205 omfattar inte frizoner enligt punkt 1."
14. Artikel 212a skall ersättas med följande:
"Artikel 212a
När det i tullagstiftningen föreskrivs en gynnsam behandling i tullhänseende för varor med anledning av deras beskaffenhet eller deras användning för särskilda ändamål, eller fullständig eller partiell befrielse från import- eller exporttullar med stöd av artiklarna 21, 82, 145 eller 184-187, skall den gynnsamma behandlingen eller befrielsen även tillämpas då en tullskuld har uppkommit i enlighet med artiklarna 202-205, 210 eller 211, om den berörda partens uppträdande inte låter förmoda bedrägligt förfarande eller påtaglig försummelse och om denne kan styrka att de övriga villkoren för tillämpning av den gynnsamma behandlingen eller befrielsen är uppfyllda."
15. I artikel 215 skall följande punkt läggas till:
"4. Om en tullmyndighet konstaterar att en tullskuld har uppkommit i en annan medlemsstat, i enlighet med artikel 202, skall tullskulden, om skuldbeloppet är lägre än 5000 euro, anses ha uppkommit i den medlemsstat där den konstaterades."
16. I artikel 220.2 skall punkt b ersättas med följande:
"b) Det tullbelopp som enligt lag skall erläggas har inte bokförts på grund av ett misstag från tullmyndigheternas sida och gäldenären kunde inte rimligen ha upptäckt detta, eftersom denne för sin del handlat i god tro och följt bestämmelserna i den gällande lagstiftningen i fråga om tulldeklarationen.
Om en vara erhåller förmånsbehandling på grundval av ett system för administrativt samarbete mellan tullmyndigheter som omfattar myndigheter i tredje land, skall ett ursprungsintyg som utfärdats av dessa myndigheter, om det skulle visa sig vara felaktigt, betraktas som ett misstag som inte rimligen kunde ha upptäckts på det sätt som avses i första stycket.
Utfärdande av ett felaktigt ursprungsintyg skall emellertid inte anses utgöra ett misstag när det grundar sig på felaktiga uppgifter från exportören, utom t.ex. i sådana fall då det är uppenbart att de utfärdande myndigheterna var eller borde ha varit medvetna om att varorna inte uppfyllde villkoren för förmånsbehandling.
Gäldenären kan åberopa god tro om han kan visa att han under den period då den berörda kommersiella verksamheten pågick visade vederbörlig aktsamhet för att förvissa sig om att samtliga villkor för förmånsbehandling var uppfyllda.
Gäldenären kan dock inte åberopa god tro när kommissionen i Europeiska gemenskapernas officiella tidning har offentliggjort ett yttrande om att det finns välgrundade tvivel om huruvida det land som omfattas av förmånsordningen tillämpar denna korrekt."
17. I artikel 221 skall punkt 3 ersättas med följande punkter:
"3. Underrättelse till gäldenären får inte ske senare än tre år efter den dag då tullskulden uppkom. Denna tidsfrist upphör att löpa från det att ett överklagande enligt artikel 243 inges till och med det att överklagandeförfarandet avslutas.
4. När tullskulden har uppkommit på grund av en handling som när den utfördes skulle ha kunnat ge upphov till straffrättsliga påföljder, får på de villkor som anges i de gällande bestämmelserna, underrättelsen till gäldenären lämnas efter det att treårsfristen enligt punkt 3 har löpt ut."
18. I artikel 222 skall punkt 2 ersättas med följande:
"2. Det kan också enligt kommittéförfarandet fastställas i vilka fall och på vilka villkor gäldenären kan beviljas uppskov med att betala tullarna, nämligen
- när en ansökan om eftergift framställs i enlighet med artiklarna 236, 238 eller 239, eller
- när varor tas i beslag för att därefter förverkas i enlighet med artikel 233c andra strecksatsen eller artikel 233d, eller
- när tullskulden uppkom i enlighet med artikel 203 och det finns flera gäldenärer."
19. Artiklarna 247, 248 och 249 skall ersättas med följande artiklar:
"Artikel 247
De åtgärder som krävs för att genomföra denna kodex, inklusive för tillämpningen av den förordning som avses i artikel 184, med undantag av avdelning VIII och om inte annat följer av artiklarna 9 och 10 i rådets förordning (EEG) nr 2658/87(7) och av artikel 248 i denna förordning, skall antas i enlighet med det föreskrivande förfarande som avses i artikel 247a.2 och med iakttagande av gemenskapens internationella åtaganden.
Artikel 247a
1. Kommissionen skall biträdas av en tullkodexkommitté (nedan kallad kommittén).
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 248
De åtgärder som krävs för att genomföra artiklarna 11, 12 och 21 skall antas i enlighet med den förvaltningskommitté som avses i artikel 248a.2.
Artikel 248a
1. Kommissionen skall biträdas av en tullkodexkommitté (nedan kallad kommittén).
2. När det hänvisas till denna punkt skall artiklarna 4 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 4.3 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 249
Kommittén får behandla alla de frågor om tullagstiftningen som tas upp av ordföranden, antingen på dennes initiativ eller på begäran av företrädaren för en medlemsstat."
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 2785/2000
av den 19 december 2000
om ändring av förordning (EG) nr 296/96 om de uppgifter som medlemsstaterna skall sända in för månatlig bokföring av de utgifter som finansieras genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) samt fastställande av vissa tillämpningsföreskrifter för rådets förordning (EG) nr 1259/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1258/1999 av den 17 maj 1999 om finansiering av den gemensamma jordbrukspolitiken(1), särskilt artiklarna 4.8, 5.3 och 7.5 i denna, och
av följande skäl:
(1) Enligt rådets beslut 2000/427/EG av den 19 juni 2000, i enlighet med artikel 122.2 i fördraget om införande av den gemensamma valutan i Grekland den 1 januari 2001(2), uppfyller Grekland de nödvändiga villkoren för att införa den gemensamma valutan.
(2) I rådets förordning (EG) nr 974/98 av den 3 maj 1998 om införande av euron(3), ändrad genom förordning (EG) nr 2596/2000(4), föreskrivs i artikel 2 andra meningen att Greklands valuta från och med den 1 januari 2001 skall vara euron.
(3) I artikel 4.1a a i kommissionens förordning (EG) nr 296/96 av den 16 februari 1996 om de uppgifter som medlemsstaterna skall sända in för månatlig bokföring av de utgifter som finansieras genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) samt fastställande av vissa tillämpningsföreskrifter för rådets förordning (EG) nr 1259/1999(5), senast ändrad genom förordning (EG) nr 2761/1999(6), föreskrivs att förskotten för utgifter, bokförda under EUGFJ:s garantisektion, skall upprättas och utbetalas i euro till deltagande medlemsstater. Förskotten som skall utbetalas i början av januari 2001 avser utgifter som verkställts under perioden 16.10.2000-30.11.2000. I Greklands fall bör dessa förskott för sista gången utbetalas i nationell valuta.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från EUGFJ-kommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 296/96 ändras på följande sätt:
1. I artikel 3.8 b skall följande läggas till:"I Greklands fall skall regeln tillämpas fr.o.m. den 1 januari 2001."
2. I artikel 4.1a c skall följande läggas till:"För utgifter som Grekland verkställt under perioden 16.10.2000-30.11.2000 skall förskotten utbetalas i nationell valutaenhet eller i nationell valuta."
Artikel 2
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2858/2000
av den 27 december 2000
om ändring av förordning (EG) nr 2125/95 om öppnande och förvaltning av tullkvoter för svampkonserver
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordningar (EG) nr 2290/2000(1), (EG) nr 2435/2000(2) och (EG) nr 2851/2000(3) om vissa medgivanden i form av gemenskapstullkvoter för vissa jordbruksprodukter och om anpassning, som en autonom övergångsåtgärd, av vissa jordbruksmedgivanden enligt Europaavtalet med, respektive, republikerna Bulgarien, Rumänien och Polen, särskilt artikel 1.3 i dessa, och
av följande skäl:
(1) I kommissionens förordning (EG) nr 2125/95(4), senast ändrad genom förordning (EG) nr 2493/98(5), fastställs tullkvoterna för svampkonserver från Polen, Rumänien och Bulgarien i bilagorna II, V respektive VI enligt rådets förordning (EG) nr 3066/95 av den 22 december 1995 om införande av vissa koncessioner i form av gemenskapstullkvoter för vissa jordbruksprodukter och om autonom anpassning under en övergångsperiod av vissa jordbrukskoncessioner som föreskrivs i Europaavtalen i syfte att beakta det jordbruksavtal som ingåtts inom ramen för de multilaterala handelsförhandlingarna under Uruguayrundan(6), senast ändrad genom förordning (EG) nr 2435/98(7).
(2) Förordning (EG) nr 3066/95 har upphävts genom förordning (EG) nr 2851/2000 och ersatts av förordningarna (EG) nr 2290/2000, (EG) nr 2435/2000 och (EG) nr 2851/2000 för respektive Bulgarien, Rumänien och Polen. Ovannämnda tullmedgivanden för svampkonserver bibehålls utan ändringar - genom förordning (EG) nr 2290/2000 och (EG) nr 2435/2000 för produkter med ursprung i Bulgarien och Rumänien, å ena sidan, och beviljas utan kvantitativa begränsningar genom förordning (EG) nr 2851/2000, för produkter med ursprung i Polen, å andra sidan. Det är därför lämpligt att ändra förordning (EG) nr 2125/95 genom att stryka alla hänvisningar till Polen, med undantag av hänvisningen till artikel 5 beträffande licensansökningar som lämnas in av traditionella importörer, för att anpassa den till dessa nya bestämmelser.
(3) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för bearbetade produkter av frukt och grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 2125/95 ändras på följande sätt:
1. Tullkvoterna för svampkonserver av Agaricus-arter enligt KN-numren 0711 90 40, 2003 10 20 och 2003 10 30, som förtecknas i bilaga I, öppnas i enlighet med de tillämpningsföreskrifter som anges i denna förordning.
Kommissionens beslut
av den 19 december 2000
om ändring av kapitel 14 i bilaga I till rådets direktiv 92/118/EEG om djurhälso- och hygienkrav för handel inom gemenskapen med produkter, som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A.I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG
[delgivet med nr K(2000) 3866]
(Text av betydelse för EES)
(2001/7/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 92/118/EEG om djurhälso- och hygienkrav för handel inom gemenskapen med produkter, som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A.I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG(1), senast ändrat genom kommissionens beslut 1999/724/EG(2), särskilt artikel 15 i detta, och
av följande skäl:
(1) Vissa översättningsskillnader mellan den tyska texten och de övriga språkversionerna bör utjämnas när det gäller gränsöverskridande handel med obearbetad gödsel. Med tanke på möjliga sjukdomsrisker är det också lämpligt att införa bättre kontroll av sådana förflyttningar.
(2) Det är nödvändigt att vid förflyttningar över gränser ta hänsyn till sjukdomssituationen i medlemsstaterna.
(3) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilaga I till rådets direktiv 92/118/EEG skall punkt 1 a i kapitel 14 del I A ersättas med följande:
"1. a) Handel med obearbetad gödsel av andra arter än fjäderfä och hästdjur skall vara förbjuden, med undantag för gödsel som:
kommer från ett område eller en anläggning där det inte finns restriktioner beträffande någon allvarlig transmissibel sjukdom
och
är avsedd att spridas under kontroll av behöriga myndigheter på mark som utgör en del av eller tillhör samma anläggning som, vare sig åtskild eller ej, ligger på båda sidor om gränsen mellan medlemstater och inom ett avstånd på cirka 20 km. För att en anläggning skall kunna godkännas måste dess ägare föra register över sådana förflyttningar över gränser. Den behöriga myndigheten skall föra register över sådana godkända anläggningar."
Artikel 2
Detta beslut träder i kraft den 1 januari 2001.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 24 januari 2001
om fastställande av en mall för förteckningarna över de enheter som godkänts av medlemsstaterna när det gäller handeln inom gemenskapen med levande djur, sperma och embryon, samt om bestämmelser avseende överlämnande av dessa förteckningar till kommissionen
[delgivet med nr K(2001) 143]
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 64/432/EEG av den 26 juni 1964 om djurhälsoproblem som påverkar handeln med nötkreatur och svin inom gemenskapen(1), senast ändrat genom direktiv 2000/20/EG(2), särskilt artikel 11.6 i detta,
med beaktande av rådets direktiv 88/407/EEG av den 14 juni 1988 om djurhälsokrav som är tillämpliga vid handel inom gemenskapen med och import av djupfryst sperma från tamdjur av nötkreatur(3), senast ändrat genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 5.2 i detta,
med beaktande av rådets direktiv 89/556/EEG av den 25 september 1989 om djurhälsovillkor för handel inom gemenskapen med och import från tredje land av embryon från tamdjur av nötkreatur(4), senast ändrat genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 5.3 i detta,
med beaktande av rådets direktiv 90/426/EEG av den 26 juni 1990 om djurhälsovillkor vid förflyttning och import av hästdjur från tredje land(5), senast ändrat genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 7 i detta,
med beaktande av rådets direktiv 90/429/EEG av de 26 juni 1990 om djurhälsokrav som är tillämpliga vid handel inom gemenskapen med och import av sperma från tamdjur av svin(6), senast ändrat genom beslut 1999/608/EG(7), särskilt artikel 5.3 i detta,
med beaktande av rådets direktiv 91/68/EEG av den 28 januari 1991 om djurhälsovillkor för handeln med får och getter inom gemenskapen(8), senast ändrat genom beslut 94/953/EG(9), särskilt artikel 2.9 i detta, och
av följande skäl:
(1) Det är tillåtet att bedriva handel inom gemenskapen med nötkreatur, svin, får, getter och hästdjur från sådana uppsamlingscentraler som godkänts av de behöriga myndigheterna i de medlemsstater där de är belägna.
(2) Det är tillåtet att bedriva handel inom gemenskapen med sperma från tama arter av nötkreatur och svin från sådana centraler som godkänts av de behöriga myndigheterna i de medlemsstater där de är belägna.
(3) Det är tillåtet att bedriva handel inom gemenskapen med embryon och ägg från arter av nötkreatur om dessa embryon och ägg har samlats in, bearbetats och lagrats av embroysamlingsgrupper som godkänts av de behöriga myndigheterna i de medlemsstater där de är verksamma.
(4) Varje enskild medlemsstat bör till kommissionen och övriga medlemsstater sända förteckningar över de uppsamlingscentraler, seminstationer och embryosamlingsgrupper i det egna landet som medlemsstaten har godkänt.
(5) För att underlätta åtkomsten till uppdaterade förteckningar för gemenskapen är det nödvändigt att harmonisera såväl mallen för dessa förteckningar som det sätt på vilket de skickas.
(6) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förteckningarna över de enheter som anges i bilaga I skall skickas till kommissionen i något av följande format: Word 97 (eller tidigare versioner), Excel 97 (eller tidigare versioner) eller pdf; filerna skall skickas till följande e-postadress: Inforvet@cec.eu.int.
Förteckningarna skall vara utformande enligt mallarna i bilaga II.
Inom ramen för Ständiga veterinärkommitténs arbete skall kommissionen underrätta medlemsstaterna om alla eventuella ändringar av ovanstående format eller av den adress till vilken filerna skall skickas.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 16 januari 2001
om ändring av avfallsförteckningen i beslut 2000/532/EG
[delgivet med nr K(2001) 108]
(Text av betydelse för EES)
(2001/118/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 75/442/EEG av den 15 juli 1975 om avfall(1), senast ändrat genom kommissionens beslut 96/350/EG(2), särskilt artikel 1 a i detta,
med beaktande av rådets direktiv 91/689/EEG av den 12 december 1991 om farligt avfall(3), ändrat genom direktiv 94/31/EG(4), särskilt artikel 1.4 andra strecksatsen i detta, och
av följande skäl:
(1) Kommissionens beslut 2000/532/EG(5) av den 3 maj 2000 om ersättning av beslut 94/3/EG om en förteckning över avfall i enlighet med artikel 1 a i rådets direktiv 75/442/EEG om avfall, och rådets beslut 94/904/EG om upprättande av en förteckning över farligt avfall i enlighet med artikel 1.4 i rådets direktiv 91/689/EEG om farligt avfall bör ändras mot bakgrund av de anmälningar som inkommit från medlemsstaterna i enlighet med artikel 1.4 andra strecksatsen i direktiv 91/689/EEG.
(2) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som upprättats i enlighet med artikel 18 i direktiv 75/442/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Beslut 2000/532/EG ändras på följande sätt:
1. Artikel 2 skall ersättas med följande:
"Artikel 2
Avfall som klassificeras som farligt anses uppvisa en eller flera av de egenskaper som avses i bilaga 3 till direktiv 91/689/EEG och, vad beträffar H3-H8, H10(6) och H11 i denna bilaga, en eller flera av följande egenskaper:
- flampunkt <= 55 °C,
- ett eller flera ämnen som klassificeras(7) som mycket giftiga vid en total koncentration >= 0,1 %,
- ett eller flera ämnen som klassificeras som giftiga vid en total koncentration >= 3 %,
- ett eller flera ämnen som klassificeras som hälsoskadliga vid en total koncentration >= 25 %,
- ett eller flera frätande ämnen som klassificeras som R35 vid en total koncentration >= 1 %,
- ett eller flera frätande ämnen som klassificeras som R34 vid en total koncentration >= 5 %,
- ett eller flera irriterande ämnen som klassificeras som R41 vid en total koncentration >= 10 %,
- ett eller flera irriterande ämnen som klassificeras som R36, R37 eller R38 vid en total koncentration >= 20 %,
- ett ämne som är känt för att vara cancerframkallande (kategori 1 eller 2) vid en koncentration >= 0,1 %,
- ett ämne som är känt för att vara cancerframkallande (kategori 3) vid en koncentration >= 1 %,
- ett ämne som är skadligt för fortplantningen (kategori 1 eller 2) och som klassificeras som R60 eller R61 vid en koncentration >= 0,5 %,
- ett ämne som är skadligt för fortplantningen (kategori 3) och som klassificeras som R62 eller R63 vid en koncentration >= 5 %,
- ett mutagent ämne (kategori 1 eller 2) som klassificeras som R46 vid en koncentration >= 0,1 %,
- ett mutagent ämne (kategori 3) som klassificeras som R40 vid en koncentration >= 1 %."
2. Bilagan skall ersättas med texten i bilagan till detta beslut.
Artikel 2
Det här beslutet skall tillämpas från och med den 1 januari 2002.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 22 februari 2001
om fastställande av provtagningsplaner och diagnostiska metoder för påvisande och bekräftelse av vissa fisksjukdomar och om upphävande av beslut 92/532/EEG
[delgivet med nr K(2001) 426]
(Text av betydelse för EES)
(2001/183/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/67/EEG av den 28 januari 1991 om djurhälsovillkor för utsläppande på marknaden av djur och produkter från vattenbruk(1), senast ändrat genom direktiv 98/45/EG(2), särskilt artikel 15 i detta, och
av följande skäl:
(1) Provtagningsplanerna och de diagnostiska metoderna för påvisande och bekräftelse av vissa fisksjukdomar fastställs i kommissionens beslut 92/532/EEG(3), senast ändrat genom kommissionens beslut 96/240/EG(4).
(2) Sedan beslut 92/532/EEG fattades har både tekniska och vetenskapliga framsteg skett, och direktiv 91/67/EEG har ändrats. Detta innebär att provtagningsplaner och diagnostiska metoder måste moderniseras.
(3) Ändringarna gäller undersökning och identifiering av virus som orsakar viral hemorragisk septikemi (VHS) och smittsam hematopoetisk nekros (IHN) samt anpassning till ändringarna av direktiv 91/67/EEG.
(4) Gemenskapens referenslaboratorium för fisksjukdomar, som inrättades genom rådets direktiv 93/53/EEG(5), har rådfrågats.
(5) De provtagningsplaner och diagnostiska metoder för påvisande och bekräftelse av vissa fisksjukdomar som infördes genom beslut 92/532/EEG måste för klarhetens skull upphävas.
(6) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Provtagningsplaner och diagnostiska metoder för påvisande och bekräftelse av viral hemorragisk septikemi (VHS) och infektiös hematopoetisk nekros (IHN) fastställs i bilagan.
Artikel 2
Detta beslut upphäver beslut 92/532/EEG.
Artikel 3
Detta beslut riktar sig till alla medlemsstater.
Rådets beslut
av den 23 juli 2001
om ändring av beslut 90/424/EEG om utgifter inom veterinärområdet
(2001/572/EG)
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets beslut 90/424/EEG av den 26 juni 1990 om utgifter inom veterinärområdet(1), särskilt artikel 24.1 och 24.2 i detta,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) I beslut 90/424/EEG fastställs att det är möjligt att ge finansiellt stöd från gemenskapen för bekämpning och övervakning av de sjukdomar som förtecknas i en bilaga till det beslutet.
(2) Förteckningen kan kompletteras eller ändras med hänsyn till hur hälsosituationen utvecklas i gemenskapen.
(3) Infektiös laxanemi är en ny sjukdom som första gången förekom i gemenskapen 1998 och som kan orsaka betydande förluster för laxodlingsnäringen.
(4) Det är viktigt att infektiös laxanemi bekämpas i syfte att förhindra dess spridning till andra områden.
(5) Bluetongue är en insektsburen virussjukdom hos får, getter, nötkreatur och andra idisslare.
(6) Bluetongue har konsekvenser på internationell nivå för förflyttning av levande djur av känsliga arter eftersom bluetongue finns upptagen på förteckning A från Internationella byrån för epizootiska sjukdomar.
(7) År 1998 kom bluetongue in på gemenskapens område från utlandet och spreds via infekterade vektorer.
(8) Vissa områden inom gemenskapen måste, på grund av klimatförhållanden, betraktas som högriskområden för bluetongue.
(9) I beslut 90/424/EEG föreskrivs nödåtgärder som förorsakas av förekomst av bluetongue. Det krävs även ett finansiellt stöd från gemenskapen för övervakning och vissa bekämpningsåtgärder, bland annat vaccinering i högriskområden för bluetongue eller i områden där sjukdomen är endemisk.
(10) Med hänsyn till ovanstående bör infektiös laxanemi och bluetongue läggas till i den ovan nämnda förteckningen, så att finansiellt stöd från gemenskapen kan erhållas för genomförande av programmen för utrotning och övervakning av dessa sjukdomar. Särskilda kriterier för bluetongue bör antas för att göra det möjligt att verkställa den finansiella åtgärd som avses i artikel 24.1.
(11) För att det finansiella stödet från gemenskapen skall kunna ges, måste de relevanta bestämmelser följas som anges i beslut 90/424/EEG och, när det gäller infektiös laxanemi, i rådets direktiv 93/53/EEG av den 24 juni 1993 om gemenskapens minimiåtgärder för bekämpning av vissa fisksjukdomar(2).
(12) Rådets förordning (EG) nr 2792/1999 av den 17 december 1999 om föreskrifter och villkor för gemenskapens strukturstöd inom fiskerisektorn(3), särskilt artikel 15.3 g i denna, utgör den rättsliga grunden för säkerställande av finansiellt stöd när det gäller infektiös laxanemi. Bestämmelserna i avdelning III i rådets förordning (EG) nr 1260/1999 av den 21 juni 1999 om allmänna bestämmelser för strukturfonderna(4) skall därför tillämpas genom undantag från bestämmelserna i artikel 24.5, 24.6, andra meningen, 24.8 och 24.9 i beslut 90/424/EEG.
(13) Beslut 90/424/EEG bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilagan till beslut 90/424/EEG skall följande strecksatser läggas till i Grupp 1: "- Infektiös laxanemi(5)
- Bluetongue i högriskområden eller områden där sjukdomen är endemisk(6)".
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Rådets beslut
av den 23 juli 2001
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT,
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/689/EEG av den 12 december 1991 om farligt avfall(1), särskilt artikel 1.4 i detta,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) En gemenskapsförteckning över avfall upprättades genom kommissionens beslut 2000/532/EG av den 3 maj 2000 om ersättning av beslut 94/3/EG om en förteckning över avfall i enlighet med artikel 1 a i rådets direktiv 75/442/EEG om avfall, och rådets beslut 94/904/EG om upprättande av en förteckning över farligt avfall i enlighet med artikel 1.4 i rådets direktiv 91/689/EEG om farligt avfall(2).
(2) Enligt artikel 1.4 i direktiv 91/689/EEG skall medlemsstaterna till kommissionen anmäla allt avfall som inte är upptaget i förteckningen över farligt avfall, och som de anser företer någon eller några av de egenskaper som anges i bilaga 3 till direktivet. Flera medlemsstater har anmält avfall som innehåller klorsilaner, avfall som innehåller silikoner och byggmaterial som innehåller asbest och begärt att förteckning över farligt avfall skall anpassas.
(3) För tydlighetens skull bör det uttryckligen anges att uteslutande fett- och oljeblandningar från oljeavskiljare som endast innehåller ätliga oljor och fetter får betraktas som icke-farliga.
(4) Beslut 2000/532/EG bör följaktligen ändras.
(5) De åtgärder som föreskrivs i detta beslut är inte förenliga med yttrandet från den kommitté som upprättats i enlighet med artikel 18 i direktiv 75/442/EEG av den 15 juli 1975 om avfall(3). De måste därför, i enlighet med artikel 18 fjärde stycket i direktiv 75/442/EEG, antas av rådet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till beslut 2000/532/EG skall ändras i enlighet med bilagan till det här beslutet.
Artikel 2
Detta beslut skall tillämpas från och med den 1 januari 2002.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 6 augusti 2001
om uppdatering av beslut 2000/112/EG om fördelning av beredskapslager av antigener mellan antigenbanker
[delgivet med nr K(2001) 2472]
(Text av betydelse för EES)
(2001/660/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets beslut 90/424/EEG av den 26 juni 1990 om utgifter inom veterinärområdet(1), senast ändrat genom beslut 2001/12/EG(2), särskilt artikel 14 i detta,
med beaktande av rådets beslut 91/666/EEG av den 11 december 1991 om att inom gemenskapen upprätta beredskapslager av vacciner mot mul- och klövsjuka(3), senast ändrat genom kommissionens beslut 2001/181/EG(4), särskilt artiklarna 7 i detta, och
av följande skäl:
(1) I enlighet med beslut 91/666/EEG ingår inköp av antigener som ett led i gemenskapens åtgärder för att upprätta beredskapslager av vacciner mot mul- och klövsjuka.
(2) I bilaga I till beslut 91/666/EEG anges närmare vilka mängder och subtyper av antigener till mul- och klövsjukeviruset som skall lagras i gemenskapens beredskapslager.
(3) Genom kommissionens beslut 93/590/EG(5), senast ändrat genom beslut 2000/112/EG(6), fastställs bestämmelser för inköp av mul- och klövsjukevirusantigen A5, A22 och O1.
(4) Genom kommissionens beslut 97/348/EG(7), senast ändrat genom beslut 2000/112/EG, fastställs bestämmelser för inköp av mul- och klövsjukevirusantigen A22-Iraq, C1 och ASIA1.
(5) Genom kommissionens beslut 2000/77/EG(8), fastställs bestämmelser för inköp av ett antal mängder av mul- och klövsjukevirusantigen A Iran 96, A Iran 99, A Malaysia 97, SAT 1, SAT 2 (stammar från östra respektive södra Afrika) och SAT 3.
(6) Genom kommissionens beslut 2000/569/EG(9), fastställs bestämmelser för inköp av ytterligare mängder av mul- och klövsjukevirusantigen A22-Iraq, O1-Manisa, ASIA 1-Shamir, A Malaysia 97, SAT 1, SAT 2 (stammar från östra respektive södra Afrika) och SAT 3.
(7) Efter skriftliga uppgifter från leverantören om tilldelning och fördelning till de godkända anläggningarna av antigen som inköpts enligt beslut 2000/569/EG är det också lämpligt att uppdatera bilagan till beslut 2000/112/EG med närmare uppgifter om antigenreservernas fördelning mellan de antigenbanker som upprättats inom ramen för gemenskapens åtgärder för att skapa beredskapslager av vacciner mot mul- och klövsjuka och att ändra kommissionens beslut 93/590/EG och 97/348/EG.
(8) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till beslut 2000/112/EG skall ersättas med bilagan till detta beslut.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Rådets rambeslut
av den 28 maj 2001
om bekämpning av bedrägeri och förfalskning som rör andra betalningsmedel än kontanter
(2001/413/RIF)
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA RAMBESLUT
med beaktande av Fördraget om Europeiska unionen, särskilt artikel 34.2 b i detta,
med beaktande av kommissionens initiativ(1),
med beaktande av Europaparlamentets yttrande(2), och
av följande skäl:
(1) Bedrägerier och förfalskningar som rör andra betalningsmedel än kontanter sker ofta på internationell nivå.
(2) Det arbete som olika internationella organisationer (t.ex. Europarådet, G8-gruppen, OECD, Interpol och FN) utför är betydelsefullt, men det behöver kompletteras med åtgärder från Europeiska unionens sida.
(3) Rådet anser att vissa former av bedrägeri som rör andra betalningsmedel än kontanter är så allvarliga och utvecklas på ett sådant sätt att det krävs övergripande lösningar. Rekommendation nr 18 i handlingsplanen för bekämpande av den organiserade brottsligheten(3), godkänd av Europeiska rådet i Amsterdam den 16-17 juni 1997, samt punkt 46 i rådets och kommissionens handlingsplan för att på bästa sätt genomföra bestämmelserna i Amsterdamfördraget om upprättande av ett område med frihet, säkerhet och rättvisa(4), godkänd av Europeiska rådet i Wien den 11-12 december 1998, innebär att åtgärder måste vidtas på detta område.
(4) Eftersom målen för detta rambeslut, nämligen att säkerställa att bedrägeri och förfalskning som rör alla andra betalningsmedel än kontanter anses vara straffbara gärningar som omfattas av effektiva, proportionella och avskräckande påföljder i alla medlemsstater, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna med hänsyn till dessa brotts internationella karaktär utan därför bättre kan uppnås på gemenskapsnivå, får gemenskapen anta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i Fördraget om upprättandet av Europeiska gemenskapen. I enlighet med proportionalitetsprincipen så som den kommer till uttryck i den artikeln går detta rambeslut inte utöver vad som är nödvändigt för att uppnå de målen.
(5) Detta rambeslut bör bidra till kampen mot bedrägeri och förfalskning som rör andra betalningsmedel än kontanter tillsammans med andra rättsakter som rådet redan har antagit, t.ex. gemensam åtgärd 98/428/RIF(5) om inrättande av ett europeiskt rättsligt nätverk, gemensam åtgärd 98/733/RIF(6) om att göra deltagande i en kriminell organisation i Europeiska unionens medlemsstater till ett brott, gemensam åtgärd 98/699/RIF(7) om penningtvätt, identifiering, spårande, spärrande, beslag och förverkande av hjälpmedel och vinning av brott samt beslut av den 29 april 1999 om utökande av Europols mandat till att omfatta bekämpning av penningförfalskning och förfalskning av betalningsmedel(8).
(6) Kommissionen överlämnade till rådet den 1 juli 1998 meddelandet "En ram för åtgärder för att bekämpa bedrägeri och förfalskning som rör andra betalningsmedel än kontanter", i vilket det förespråkas en EU-politik som omfattar både förebyggande och repressiva aspekter av problemet.
(7) Meddelandet innehåller ett utkast till gemensam åtgärd som är en del av denna övergripande strategi och utgör utgångspunkten för detta rambeslut.
(8) Det är nödvändigt att en beskrivning av de olika typer av beteenden som bör kriminaliseras i samband med bedrägeri och förfalskning som rör andra betalningsmedel än kontanter omfattar all den verksamhet som i detta avseende utgör hotet från den organiserade brottsligheten.
(9) Det är nödvändigt att dessa typer av beteenden anses vara straffbara gärningar i samtliga medlemsstater och att effektiva, proportionella och avskräckande påföljder införs för fysiska och juridiska personer som har begått eller är ansvariga för sådana brott.
(10) Avsikten med att ge straffrättsligt skydd åt i första hand betalningsinstrument med en särskild form av skydd mot efterbildning eller missbruk är att operatörerna skall uppmuntras att förse de betalningsinstrument de ger ut med detta skydd och att instrumentet därmed förses med en förebyggande faktor.
(11) Det är nödvändigt att medlemsstaterna ger varandra största möjliga ömsesidiga bistånd och samråder med varandra när fler än en medlemsstat är behöriga i fråga om samma brott.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Definitioner
I detta rambeslut avses med
a) betalningsinstrument: ett fysiskt instrument annat än lagliga betalningsmedel (legal tender) (sedlar och mynt) som genom sin särskilda karaktär, enskilt eller tillsammans med ett annat (betalnings)instrument, gör det möjligt för innehavaren eller användaren att föra över pengar eller ett penningvärde, t.ex. kreditkort, eurocheckkort, andra av finansinstitut utgivna kort, resecheckar, eurocheckar, andra checkar och växlar som är skyddade mot efterbildning eller bedräglig användning, t.ex. genom sin utformning, kod eller undertecknande,
b) juridisk person: varje enhet som har denna ställning enligt tillämplig lagstiftning, med undantag av stater eller andra offentliga organ vid utövandet av de befogenheter som de har i egenskap av statsmakter samt internationella offentliga organisationer.
Artikel 2
Brott i samband med betalningsinstrument
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att följande handlingar är straffbara när de är uppsåtliga, åtminstone när det gäller kreditkort, eurocheckkort, andra kort utgivna av finansinstitut, resecheckar, eurocheckar, andra checkar och växlar:
a) Stöld eller annat olovligt tillgrepp av ett betalningsinstrument.
b) Hel- eller delförfalskning av ett betalningsinstrument med syfte att använda det för bedrägeri.
c) Mottagande, förskaffande, transport, försäljning eller överlämnande till en annan person eller innehav av ett betalningsinstrument som stulits eller olovligen tillgripits eller som är helt eller delvis förfalskat med syfte att använda det för bedrägeri.
d) Bedräglig användning av ett betalningsinstrument som stulits eller olovligen tillgripits eller som är helt eller delvis förfalskat.
Artikel 3
Datorrelaterade brott
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att följande handlingar är straffbara när de är uppsåtliga:
- att utan rätt mata in, ändra, radera, eller undertrycka datoriserade uppgifter, särskilt identifieringsuppgifter, eller
- att utan rätt ingripa i ett dataprograms eller datasystems funktion.
Artikel 4
Brottslighet i samband med särskilt anpassad utrustning
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att följande handlingar är straffbara när de är uppsåtliga:
Bedräglig tillverkning, mottagande, anskaffande, försäljning eller överlämnande till annan person eller innehav av
- redskap, föremål, datorprogram och alla andra instrument som är särskilt avsedda för att föröva något av de brott som avses i artikel 2 b,
- datorprogram som är avsedda för att begå något av de brott som avses i artikel 3.
Artikel 5
Deltagande, anstiftan och försök
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att deltagande i och anstiftan till sådana handlingar som avses i artiklarna 2-4 eller försök till sådana handlingar som avses i artikel 2 a, 2 b, 2 d och artikel 3 är straffbara.
Artikel 6
Påföljder
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att de handlingar som avses i artiklarna 2-5 är belagda med straffrättsliga påföljder som är effektiva, proportionella och avskräckande och som, åtminstone i allvarliga fall, omfattar påföljder som är frihetsberövande och kan medföra utlämning.
Artikel 7
Juridiska personers ansvar
1. Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att juridiska personer kan ställas till ansvar för sådana handlingar som avses i artikel 2 b-d och artiklarna 3-4 och som till deras förmån begås av varje person som agerar antingen enskilt eller som en del av den juridiska personens organisation och har en ledande ställning inom den juridiska personen, grundad på
- befogenhet att företräda den juridiska personen, eller
- befogenhet att fatta beslut på den juridiska personens vägnar, eller
- befogenhet att utöva kontroll inom den juridiska personen,
samt för medhjälp eller anstiftan till ett sådant brott.
2. Utom i de fall som avses i punkt 1 skall varje medlemsstat vidta nödvändiga åtgärder för att säkerställa att en juridisk person kan ställas till ansvar när brister i övervakning eller kontroll som skall utföras av en sådan person som avses i punkt 1 har gjort det möjligt för en person, som är underställd den juridiska personen, att begå ett sådant brott som avses i artikel 2 b-d och artiklarna 3-4.
3. Den juridiska personens ansvar enligt punkterna 1 och 2 utesluter inte lagföring av fysiska personer som är gärningsmän, anstiftare eller medhjälpare till de handlingar som avses i artikel 2 b-d och artiklarna 3-4.
Artikel 8
Påföljder för juridiska personer
1. Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att en juridisk person som har ställts till ansvar i enlighet med artikel 7.1 kan bli föremål för effektiva, proportionella och avskräckande påföljder, som skall innefatta bötesstraff eller administrativa avgifter och som kan innefatta andra påföljder, t.ex.
a) fråntagande av rätt till offentliga förmåner eller stöd,
b) tillfälligt eller permanent näringsförbud,
c) rättslig övervakning,
d) rättsligt beslut om avveckling av verksamheten.
2. Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att en juridisk person som har ställts till ansvar i enlighet med artikel 7.2 kan bli föremål för effektiva, proportionella och avskräckande påföljder eller åtgärder.
Artikel 9
Behörighet
1. Varje medlemsstat skall vidta nödvändiga åtgärder för att fastställa sin behörighet rörande brott enligt artiklarna 2, 3, 4 och 5 när brott har begåtts
a) helt eller delvis på medlemsstatens territorium,
b) av en av dess medborgare, dock med förbehåll för att den medlemsstatens lagstiftning kan kräva att gärningen är straffbar även i det land där den begicks, eller
c) till förmån för en juridisk person som har sitt säte inom medlemsstatens territorium.
2. Om inte annat följer av artikel 10, kan en medlemsstat besluta att inte tillämpa behörighetsregeln eller att endast i särskilda fall eller under särskilda omständigheter tillämpa regeln i
- punkt 1 b,
- punkt 1 c.
3. Medlemsstaterna skall vederbörligen underrätta rådets generalsekretariat om de beslutar att tillämpa punkt 2, om så är lämpligt med angivande av de särskilda fall eller omständigheter då beslutet gäller.
Artikel 10
Utlämning och åtal
1. a) Varje medlemsstat som enligt sin lag inte utlämnar sina egna medborgare skall vidta nödvändiga åtgärder för att fastställa sin behörighet rörande brott enligt artiklarna 2, 3, 4 och 5 när de begås av en av dess egna medborgare utanför dess territorium.
b) Varje medlemsstat skall, när en av dess medborgare anklagas för att i en annan medlemsstat ha begått ett brott som innefattar de handlingar som beskrivs i artiklarna 2, 3, 4 och 5 och om den inte utlämnar denna person till den andra medlemsstaten enbart på grund av dennes nationalitet, lägga fram fallet för sina behöriga myndigheter i syfte att om så är lämpligt väcka åtal. För att möjliggöra att åtal väcks skall akter, information och bevisföremål som rör brottet överlämnas enligt förfarandena i artikel 6.2 i Europeiska utlämningskonventionen av den 13 december 1957. Den ansökande medlemsstaten skall informeras om det åtal som väcks och om dess resultat.
2. I denna artikel skall begreppet medborgare i en medlemsstat tolkas i enlighet med en eventuell förklaring som denna stat avgivit enligt artikel 6.1 b och c i Europeiska utlämningskonventionen.
Artikel 11
Samarbete mellan medlemsstaterna
1. Medlemsstaterna skall i enlighet med tillämpliga konventioner, multilaterala eller bilaterala avtal eller arrangemang i så hög grad som möjligt bistå varandra när det gäller förfaranden som rör brott enligt detta rambeslut.
2. Om flera medlemsstater är behöriga i fråga om brott som avses i detta rambeslut skall dessa stater samråda med varandra i syfte att samordna sina insatser för en effektiv lagföring.
Artikel 12
Informationsutbyte
1. Medlemsstaterna skall antingen utse operativa kontaktpunkter eller också kan de använda befintliga operativa strukturer för informationsutbyte samt för annan kontakt mellan medlemsstaterna för att tillämpa detta rambeslut.
2. Varje medlemsstat skall meddela rådets generalsekretariat eller kommissionen vilket eller vilka organ som utgör kontaktpunkt enligt punkt 1. Generalsekretariatet skall meddela övriga medlemsstater vilka dessa kontaktpunkter är.
Artikel 13
Territoriell tillämpning
Detta rambeslut skall tillämpas i Gibraltar.
Artikel 14
Genomförande
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta rambeslut senast den 2 juni 2003.
2. Senast den 2 juni 2003 skall medlemsstaterna till rådets generalsekretariat och till Europeiska gemenskapernas kommission överlämna texten till de bestämmelser genom vilka de skyldigheter som åvilar dem enligt detta rambeslut överförs till nationell lag. Senast den 2 september 2003 skall rådet mot bakgrund av en rapport som upprättats på grundval av dessa upplysningar och en skriftlig rapport från kommissionen bedöma i vilken utsträckning medlemsstaterna har vidtagit nödvändiga åtgärder för att följa detta rambeslut.
Artikel 15
Ikraftträdande
Detta rambeslut träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets direktiv 2001/108/EG
av den 21 januari 2002
om ändring av rådets direktiv 85/611/EEG om samordning av lagar och andra författningar som avser företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag), vad gäller fondföretags investeringar
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 47.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Räckvidden av rådets direktiv 85/611/EEG(4) var ursprungligen begränsad till sådana företag för kollektiva investeringar av den öppna typen som utbjuder sina andelar till allmänheten inom gemenskapen och som har som enda syfte att investera i överlåtbara värdepapper (fondföretag). I ingressen till direktiv 85/611/EEG såg man framför sig att sådana företag för kollektiva investeringar som inte omfattades av direktivet skulle kunna bli föremål för samordning i ett senare skede.
(2) Med hänsyn till utvecklingen på marknaden bör fondföretagens investeringsmöjligheter utökas till att omfatta andra, tillräckligt likvida, finansiella instrument än överlåtbara värdepapper. Finansiella instrument som kan ingå som tillgångar i ett fondföretags värdepappersportfölj anges i detta direktiv. Att investera så att en portfölj återspeglar ett visst index är en förvaltningsteknik.
(3) Den i detta direktiv angivna definitionen av överlåtbara värdepapper gäller endast för detta direktiv och påverkar inte på något sätt de definitioner som används i nationell lagstiftning i andra sammanhang, exempelvis när det gäller beskattning. Denna definition omfattar följaktligen inte aktier och andra värdepapper som motsvarar aktier och som emitteras av sådana organ som hypoteksinstitut och industri- och utvecklingsfonder, där äganderätten i praktiken inte kan överföras på annat sätt än att det emitterande organet återköper dem.
(4) Penningmarknadsinstrument omfattar de kategorier av överlåtbara instrument som normalt inte handlas på reglerade marknader utan som omsätts på penningmarknaden, till exempel statsskuldväxlar, kommunala skuldväxlar, bankcertifikat, företagscertifikat, omsättningsbara medelfristiga skuldväxlar och bankaccepter.
(5) Det är lämpligt att säkerställa att begreppet "reglerad marknad" i detta direktiv stämmer överens med det i direktiv 93/22/EEG av den 10 maj 1993 om investeringstjänster inom värdepappersområdet(5).
(6) Fondföretag bör tillåtas att investera sina tillgångar i andelar i andra fondföretag och/eller andra företag för kollektiva investeringar av den öppna typen som också investerar i sådana likvida, finansiella tillgångar som omnämns i detta direktiv och som tillämpar principen om riskspridning. Det är nödvändigt att fondföretag och andra företag för kollektiva investeringar som fondföretag investerar i är föremål för effektiv tillsyn.
(7) Utvecklingen av möjligheterna för ett fondföretag att investera i fondföretag och i andra företag för kollektiva investeringar bör underlättas. Det är därför väsentligt att se till att en sådan investeringsverksamhet inte minskar skyddet för investerarna. På grund av fondföretagens ökade möjligheter att investera i andelar i andra fondföretag och/eller företag för kollektiva investeringar är det nödvändigt att fastställa vissa regler om kvantitativa begränsningar, tillhandahållande av information och förhindrande av uppkomsten av s.k. kaskadfonder.
(8) För att beakta marknadsutvecklingen och mot bakgrund av genomförandet av den ekonomiska och monetära unionen, bör fondföretag tillåtas att investera i inlåning. För att säkerställa en tillräcklig likviditet för sådana investeringar skall dessa tillgodohavanden kunna betalas ut på begäran eller kunna dras tillbaka. Om tillgodohavandena finns i ett kreditinstitut med säte i en icke-medlemsstat, bör detta institut omfattas av tillsynsregler likvärdiga med dem som gäller inom gemenskapslagstiftningen.
(9) Utöver det fall då ett fondföretag investerar i banktillgodohavanden i enlighet med sina fondbestämmelser eller sin bolagsordning kan det bli nödvändigt att tillåta alla fondföretag att inneha kompletterande likvida tillgångar, som exempelvis avistakonton. Innehav av sådana kompletterande likvida tillgångar kan exempelvis vara motiverat i följande fall, nämligen för att täcka löpande eller särskilda betalningar, vid försäljningar fram till dess att man kan återinvestera i överlåtbara värdepapper, penningmarknadsinstrument och/eller andra finansiella tillgångar som avses i detta direktiv samt för den tid under vilken det är absolut nödvändigt att uppskjuta investeringen i överlåtbara värdepapper, penningmarknadsinstrument eller andra finansiella tillgångar på grund av ogynnsamma marknadsvillkor.
(10) Av försiktighetsskäl är det nödvändigt att fondföretag, när det gäller investeringar som utsätter dem för en motpartsrisk, undviker orimlig koncentration till samma organ eller till organ som tillhör samma grupp.
(11) Fondföretag bör uttryckligen tillåtas att investera i finansiella derivatinstrument, såväl inom ramen för sin allmänna investeringspolicy som i syfte att säkra tillgångar, för att uppnå ett finansiellt mål eller den riskprofil som angetts i prospektet. För att säkerställa att investerarna skyddas är det nödvändigt att begränsa den maximala riskexponeringen i förhållande till finansiella derivatinstrument så att den inte överskrider det totala nettovärdet av fondföretagets portfölj. För att säkerställa ständig medvetenhet om riskerna och åtagandena vid derivattransaktioner och kontrollera att investeringsgränserna hålls, måste dessa risker och åtaganden fortlöpande mätas och övervakas. Slutligen, för att skapa ett skydd för investerarna genom tillhandahållande av information, bör fondföretagen beskriva sina strategier, metoder och sina investeringsgränser för derivattransaktioner.
(12) För OTC-derivat bör ytterligare krav ställas upp för lämplighetsbedömning av motparter och instrument, likviditet och fortlöpande värdering av positionen. Syftet med sådana ytterligare krav är att säkerställa ett tillräckligt skydd för investerarna, liknande det som de erhåller vid förvärv av derivat som handlas på reglerade marknader.
(13) Derivattransaktioner får aldrig användas för att kringgå principerna och reglerna i detta direktiv. För OTC-derivat måste det finnas ytterligare regler för riskspridningen som bör tillämpas vid exponering i förhållande till en enda motpart eller grupp av motparter.
(14) Vissa portföljförvaltningsmetoder för företag för kollektiva investeringar som främst investerar i aktier och/eller skuldebrev bygger på efterbildningen av aktieindex och/eller index för skuldebrev. Fondföretag bör tillåtas att efterbilda välkända och erkända aktieindex och/eller index för skuldförbindelser. Det kan därför vara nödvändigt att införa flexiblare riskspridningsregler för sådana fondföretag som investerar i aktier och/eller skuldförbindelser för detta ändamål.
(15) Företag för kollektiva investeringar som omfattas av detta direktiv bör inte användas för andra ändamål än kollektiva investeringar av medel från allmänheten, i enlighet med bestämmelserna i detta direktiv. I de fall som fastställs i detta direktiv får fondföretag ha dotterföretag endast när detta är nödvändigt för att utföra viss, i direktivet angiven verksamhet för fondföretagets räkning. Det är nödvändigt att säkerställa en effektiv tillsyn av fondföretag. Fondföretag skall därför tillåtas att etablera dotterföretag i tredje land endast i de fall och på de villkor som anges i detta direktiv. Den allmänna skyldigheten att uteslutande agera för att tillgodose andelsägarnas intressen och framför allt målet att förbättra kostnadseffektiviteten kan under inga omständigheter rättfärdiga åtgärder från fondföretagets sida som kan hindra de behöriga myndigheterna från att utöva en effektiv tillsyn.
(16) Det finns ett behov av att säkerställa fri saluföring över gränserna av andelar i ett större urval av företag för kollektiva investeringar, samtidigt som en enhetlig miniminivå för skydd av investerare tillhandahålls. De uppsatta målen kan därför endast nås genom att de överenskomna miniminormerna fastställs i ett bindande gemenskapsdirektiv. Detta direktiv gäller endast den erforderliga minimiharmoniseringen och går i enlighet med artikel 5 tredje stycket i fördraget inte utöver vad som är nödvändigt för att uppnå dessa mål.
(17) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(6).
(18) Kommissionen kan komma att överväga att föreslå kodifiering vid lämplig tidpunkt efter det att förslagen har antagits.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 85/611/EEG ändras härigenom på följande sätt:
1. Artikel 1.2 första strecksatsen skall ersättas med följande: "- som har till enda syfte att företa kollektiva investeringar i överlåtbara värdepapper och/eller i andra likvida finansiella tillgångar som avses i artikel 19.1 med kapital från allmänheten och som tillämpar principen om riskspridning, och"
2. I artikel 1 skall följande punkter införas: "8. I detta direktiv avses med 'överlåtbara värdepapper':
- aktier och andra värdepapper som motsvarar aktier (nedan kallade aktier),
- obligationer eller andra skuldförbindelser (nedan kallade skuldförbindelser),
- försäljningsbara värdepapper av annat slag som ger rätt att förvärva sådana överlåtbara värdepapper genom teckning eller utbyte,
med undantag för den teknik och de instrument som avses i artikel 21.
9. I detta direktiv avses med 'penningmarknadsinstrument' instrument som normalt omsätts på penningmarknaden och som är likvida och har ett värde som vid varje tidpunkt exakt kan fastställas."
3. Artikel 19.1 a skall ersättas med följande: "a) överlåtbara värdepapper och penningmarknadsinstrument som får omsättas eller omsätts på en sådan reglerad marknad som avses i artikel 1.13 i direktivet om investeringstjänster och/eller"
4. I artikel 19.1 b och c skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
5. Artikel 19.1 skall ändras på följande sätt:
- Orden "och/eller" skall läggas till i slutet av punkt d.
- Följande skall läggas till: "e) andelar i fondföretag som är auktoriserade i enlighet med detta direktiv och/eller andra företag för kollektiva investeringar enligt artikel 1.2 första och andra strecksatsen, oavsett om de är belägna i en medlemsstat eller ej, förutsatt att
- dessa andra företag för kollektiva investeringar är auktoriserade enligt lagstiftning som fastställer att de är föremål för tillsyn som av de behöriga myndigheterna med ansvar för fondföretaget anses motsvara den tillsyn som fastställs i gemenskapslagstiftningen och att det anses tillräckligt säkerställt att samarbete mellan myndigheterna sker, och
- skyddsnivån för andelsägare i det andra företaget för kollektiva investeringar motsvarar det skydd som ett fondföretags andelsägare har, särskilt genom att reglerna för separation av tillgångarna, in- och utlåning och försäljning av överlåtbara värdepapper och penningmarknadsinstrument som företaget inte innehar uppfyller villkoren i detta direktiv, och
- verksamheten i det andra företaget för kollektiva investeringar rapporteras halvårsvis och årsvis, så att det kan ske en värdering av tillgångar och skulder, intäkter och verksamhet under rapporteringsperioden, och
- de fondföretag eller andra företag för kollektiva investeringar i vars andelar förvärv planeras, enligt dessas fondbestämmelser eller bolagsordning, får investera högst 10 % av sina tillgångar i andelar i andra fondföretag eller andra företag för kollektiva investeringar, och/eller
f) inlåning i kreditinstitut, antingen som avistakonton eller som konton med högst 12 månaders uppsägningstid, under förutsättning att kreditinstitutet har sitt säte i en medlemsstat eller, om kreditinstitutet har sitt säte i tredje land, förutsatt att det omfattas av tillsynsregler som av behöriga myndigheter med ansvar för fondföretag anses motsvara dem som fastställs i gemenskapslagstiftningen, och/eller
g) finansiella derivat, inklusive motsvarande kontantavräknade instrument, som omsätts på en sådan reglerad marknad som avses i punkterna a, b och c, och/eller finansiella derivatinstrument som handlas direkt mellan parterna (nedan kallade OTC-derivat), förutsatt att
- de underliggande tillgångarna utgörs av sådana instrument som avses i denna punkt 1, finansiella index, räntesatser, växelkurser eller utländska valutor, i vilka fondföretaget kan investera utifrån de investeringsmål som det har angett i sina fondbestämmelser eller sin bolagsordning,
- motparterna vid affärer med OTC-derivat är institutioner som omfattas av tillsyn och tillhör de kategorier som godkänts av de behöriga myndigheterna med ansvar för fondföretaget, och
- OTC-derivaten är föremål för tillförlitlig och verifierbar värdering från dag till dag samt att de vid varje tidpunkt, på fondföretagets initiativ, kan säljas, lösas in eller avslutas genom en utjämnande transaktion till ett rimligt värde, och/eller
h) andra penningmarknadsinstrument än de som omsätts på en reglerad marknad och som faller under artikel 1.9, om själva emissionen eller emittenten av instrumenten reglerats i syfte att skydda investerare och sparmedel och under förutsättning att de har
- emitterats eller garanterats av en central, regional eller lokal myndighet, av en medlemsstats centralbank, av Europeiska centralbanken, av Europeiska unionen eller Europeiska investeringsbanken, av en icke-medlemsstat eller, i fråga om förbundsstater, av en av de stater som utgör förbundsstaten eller av en internationell offentlig organisation som en eller flera medlemsstater tillhör, eller
- emitterats av ett företag, vars värdepapper omsätts på de reglerade marknader som avses i punkterna a, b eller c, eller
- emitterats eller garanterats antingen av en inrättning som är föremål för tillsyn i enlighet med de kriterier som fastställs i gemenskapslagstiftningen eller av en inrättning som omfattas av och följer sådana tillsynsregler som av de behöriga myndigheterna anses minst lika stränga som de som fastställs i gemenskapslagstiftningen, eller
- emitterats av andra organ som tillhör de kategorier som godkänts av de behöriga myndigheterna med ansvar för fondföretaget förutsatt att investeringar i sådana instrument omfattas av ett investerarskydd som är likvärdigt med det som fastställs i första, andra eller tredje strecksatsen och att emittenten är ett bolag vars kapital och reserver uppgår till minst 10 miljoner euro och som lägger fram och offentliggör sin årsredovisning i enlighet med direktiv 78/660/EEG(7), är en enhet som inom en grupp företag som omfattar ett eller flera börsnoterade företag ägnar sig åt gruppens finansiering eller är en enhet som ägnar sig åt att finansiera värdepapperisering som omfattas av kreditförstärkning från en bank."
6. I artikel 19.2 a skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
7. Artikel 19.2 b och 19.3 skall utgå.
8. Artikel 20 skall utgå.
9. Artikel 21 skall ersättas med följande: "Artikel 21
1. Förvaltnings- eller investeringsbolaget måste använda ett förfarande för riskhantering som gör det möjligt för det att vid varje tidpunkt kontrollera och bedöma den risk som är knuten till positionerna och deras bidrag till portföljens allmänna riskprofil; bolaget måste använda ett förfarande som möjliggör en exakt och oberoende bedömning av värdet på OTC-derivat. Bolaget måste underrätta de behöriga myndigheterna regelbundet och i enlighet med de detaljerade regler de skall fastställa om de typer av derivatinstrument, underliggande risker, kvantitativa begränsningar liksom de metoder som valts för att beräkna de risker som åtföljer transaktioner med derivatinstrument för varje fondföretag som det förvaltar.
2. Medlemsstaterna får ge fondföretag tillstånd att använda sig av sådan teknik och sådana instrument som hänför sig till överlåtbara värdepapper och penningmarknadsinstrument på de villkor och inom de gränser medlemsstaterna föreskriver, förutsatt att sådan teknik och sådana instrument används i syfte att åstadkomma en effektiv förvaltning av värdepappersportföljen. Om denna verksamhet gäller användning av derivatinstrument skall dessa villkor och gränser överensstämma med bestämmelserna i detta direktiv.
Denna verksamhet får under inga omständigheter leda till att fondföretagen avviker från sina investeringsmål såsom de fastställts i fondföretagens fondbestämmelser, bolagsordning eller prospekt.
3. Ett fondföretag skall säkerställa att dess totala exponering som hänför sig till derivatinstrument inte överskrider dess portföljs totala nettovärde.
Exponeringen skall beräknas med hänsyn till det aktuella värdet av de underliggande tillgångarna, motpartsrisken, kommande marknadsrörelser och den tid som finns tillgänglig för att lösa in positionerna. Detta skall även gälla följande stycken.
Ett fondföretag får inom den gräns som anges i artikel 22.5 investera i finansiella derivatinstrument som ett led i sin investeringspolicy, förutsatt att exponeringen mot de underliggande tillgångarna inte sammanlagt överstiger de investeringsgränser som anges i artikel 22. När ett fondföretag investerar i indexbaserade finansiella derivatinstrument får medlemsstaterna medge att dessa investeringar sammanlagt inte behöver rymmas inom de gränser som anges i artikel 22.
När ett överlåtbart värdepapper eller ett penningmarknadsinstrument innefattar ett derivat måste detta beaktas när kraven i denna artikel skall uppfyllas.
4. Senast den 13 februari 2004 skall medlemsstaterna till kommissionen överlämna fullständig information om, och eventuella förändringar i, reglerna för de metoder som används för att beräkna riskexponering enligt punkt 3, inklusive riskexponeringen för en motpart vid transaktioner med OTC-derivat. Kommissionen skall vidarebefordra denna information till övriga medlemsstater. Sådan information kommer att vara föremål för överväganden inom kontaktkommittén i enlighet med förfarandet i artikel 53.4."
10. Artikel 22 skall ersättas med följande: "Artikel 22
1. Ett fondföretag får investera högst 5 % av sina tillgångar i överlåtbara värdepapper eller penningmarknadsinstrument som emitterats av samma organ. Ett fondföretag får investera högst 20 % av sina tillgångar i inlåning i samma organ.
Riskexponeringen mot ett fondföretags motpart vid en transaktion med OTC-derivat får inte överstiga:
- 10 % av fondföretagets tillgångar när motparten är ett kreditinstitut enligt artikel 19.1 f, eller
- 5 % av fondföretagets tillgångar i andra fall.
2. Medlemsstaterna får höja den 5-procentsgräns som anges i första meningen i punkt 1 till högst 10 %. I den mån fondföretaget investerar mer än 5 % av fondtillgångarna i överlåtbara värdepapper och penningmarknadsinstrument med samma utgivare, får det sammanlagda innehavet av sådana investeringar inte överstiga 40 % av fondtillgångarna. Begränsningen gäller inte inlåning hos och transaktioner med OTC-derivat med finansiella institut som står under tillsyn.
Trots de enskilda gränser som fastställs i punkt 1, får ett fondföretag inte kombinera
- investeringar i överlåtbara värdepapper eller penningmarknadsinstrument som emitterats av,
- inlåning hos, och/eller
4. Medlemsstaterna får höja den 5-procentsgräns som anges i punkt 1 första meningen till högst 25 % när det gäller vissa obligationer, om de är emitterade av ett kreditinstitut som har sitt säte i en medlemsstat och enligt lag omfattas av särskild offentlig tillsyn avsedd att skydda obligationsinnehavare. Särskilt skall iakttas att kapital som härrör från emissionen av sådana obligationer enligt lag måste investeras i tillgångar som, under obligationernas hela giltighetstid kan täcka de med obligationerna förenade fordringarna och som i händelse av emittentens oförmåga att fullgöra sina ekonomiska åtaganden skall med prioritet användas för återbetalning av kapital och upplupen ränta.
Om ett fondföretag investerar mer än 5 % av sina fondtillgångar i sådana obligationer som avses i första stycket och som har samma emittent, får det totala värdet av dessa investeringar inte överstiga 80 % av värdet av fondföretagets tillgångar.
Medlemsstaterna skall till kommissionen överlämna en förteckning över de ovan nämnda kategorier av obligationer och över de kategorier av emittenter, vilka enligt gällande lag och enligt sådana tillsynsregler som avses i första stycket, beviljas tillstånd att emittera sådana obligationer som uppfyller kriterierna ovan. Till förteckningen skall fogas uppgifter om vad slags garantier som erbjudits. Kommissionen skall till övriga medlemsstater genast vidarebefordra denna information jämte de kommentarer som bedömts erforderliga samt göra informationen tillgänglig för allmänheten. Sådana underrättelser kan göras till föremål för överväganden i kontaktkommittén i enlighet med förfarandet i artikel 53.4.
5. Vid beräkningen av den gräns på 40 % som anges i punkt 2 skall inte de överlåtbara värdepapper och penningmarknadsinstrument som anges i punkterna 3 och 4 beaktas.
De gränser som anges i punkterna 1, 2, 3 och 4 får inte kombineras, och investeringar i överlåtbara värdepapper och penningmarknadsinstrument emitterade av samma organ eller i inlåning eller derivatinstrument från detta organ enligt bestämmelserna i punkterna 1, 2, 3 och 4 får därför under inga förhållanden överstiga sammanlagt 35 % av ett fondföretags tillgångar.
Bolag som ingår i samma grupp för sammanställd redovisning enligt definitionen i direktiv 83/349/EEG(8) eller i enlighet med erkända internationella redovisningsregler räknas som ett organ vid beräkningen av gränserna i denna artikel.
Medlemsstaterna kan tillåta investeringar upp till en gräns på 20 % i överlåtbara värdepapper och penningmarknadsinstrument inom samma grupp."
11. Följande artikel skall läggas till: "Artikel 22a
1. Utan att det påverkar tillämpningen av de gränser som fastställs i artikel 25 får medlemsstaterna på följande villkor höja de gränser som anges i artikel 22 till högst 20 % för investeringar i aktier och/eller skuldförbindelser emitterade av samma organ, då fondföretagets investeringspolicy enligt fondbestämmelserna eller enligt bolagsordningen syftar till att efterbilda sammansättningen av ett visst aktieindex eller index för skuldförbindelser som är erkänt av de behöriga myndigheterna:
- Det skall ha en tillräckligt diversifierad sammansättning.
- Indexet skall utgöra en lämplig referens för den marknad det hänför sig till.
- Det skall offentliggöras på lämpligt vis.
2. Medlemsstaterna får höja den gräns som fastställs i punkt 1 till högst 35 % när det visar sig motiverat på grund av exceptionella marknadsvillkor särskilt på reglerade marknader där vissa överlåtbara värdepapper eller penningmarknadsinstrument i hög grad dominerar. Investeringar upp till denna gräns är bara tillåtna för en enda emittent."
12. I artikel 23.1 skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
13. Artikel 24 skall ersättas med följande: "Artikel 24
1. Ett fondföretag får förvärva andelar i fondföretag och/eller andra företag för kollektiva investeringar enligt artikel 19.1 e, under förutsättning att inte mer än 10 % av dess tillgångar investeras i andelar i ett enda fondföretag eller annat företag för kollektiva investeringar. Medlemsstaterna får höja denna gräns till högst 20 %.
2. Investeringar i andelar i företag för kollektiva investeringar som ej är fondföretag får sammanlagt inte överstiga 30 % av fondföretagets tillgångar.
Medlemsstaterna får, när ett fondföretag har förvärvat andelar i fondföretag och/eller andra företag för kollektiva investeringar, medge att värdet av dessa företags tillgångar inte behöver rymmas inom de gränser som anges i artikel 22.
3. När ett fondföretag investerar i andelar i andra fondföretag och/eller andra företag för kollektiva investeringar som direkt eller genom delegering förvaltas av samma förvaltningsbolag eller av ett annat bolag till vilket förvaltningsbolaget är anknutet via gemensam företagsledning eller ägarkontroll eller genom ett betydande direkt eller indirekt ägande får detta förvaltningsbolag eller det andra bolaget inte debitera några avgifter för teckning eller inlösen av fondföretagets investeringar i andelar i dessa andra fondföretag och/eller företag för kollektiva investeringar.
Ett fondföretag som investerar en betydande del av sina tillgångar i andra fondföretag och/eller företag för kollektiva investeringar, skall i sitt prospekt uppge maximinivån för de förvaltningskostnader som kan debiteras både fondföretaget självt och de andra fondföretag och/eller företag för kollektiva investeringar i vilka fondföretaget ämnar investera. Fondföretaget skall i sin årsrapport ange en maximal procentsats för de förvaltningskostnader som debiteras både fondföretaget självt och de fondföretag och/eller företag för kollektiva investeringar i vilka det investerar."
14. Följande artikel skall införas: "Artikel 24a
1. I prospektet skall anges vilka kategorier av tillgångar i vilka fondföretaget har tillstånd att investera. Det skall anges om transaktioner med finansiella derivatinstrument är tillåtna; i så fall måste det finnas en tydlig uppgift om huruvida dessa får utföras i syfte att säkra tillgångar eller i avsikt att nå investeringsmål och hur det möjliga resultatet av användningen av finansiella derivatinstrument kan påverka riskprofilen.
2. När ett fondföretag huvudsakligen investerar i någon annan kategori av de tillgångar som anges i artikel 19 än överlåtbara värdepapper och penningmarknadsinstrument eller efterbildar aktieindex eller index för skuldebrev enligt artikel 22a måste dess prospekt och i förekommande fall allt övrigt reklammaterial ange investeringspolicyn på framträdande plats.
3. Om nettovärdet av ett fondföretags tillgångar tenderar att ha hög volatilitet på grund av portföljens sammansättning och förvaltningsmetoderna måste detta anges på framträdande plats i prospektet och i förekommande fall i allt övrigt reklammaterial.
4. På begäran av en investerare måste förvaltningsbolaget också tillhandahålla kompletterande information om de kvantitativa gränser som gäller för fondföretagets riskhantering, de metoder som har valts för denna och den senaste utvecklingen av riskerna med och avkastningen från de viktigaste instrumentkategorierna."
15. Artikel 25.2 skall ändras enligt följande:
1. Tredje strecksatsen skall ersättas med följande: "- 25 % av andelarna i ett enskilt fondföretag och/eller annat företag för kollektiva investeringar enligt artikel 1.2 första och andra strecksatsen,"
2. Följande strecksats skall läggas till: "- 10 % av de penningmarknadsinstrument som emitterats av ett och samma organ."
16. Andra meningen i artikel 25.2 skall ersättas med följande: "De gränsvärden som anges i andra, tredje och fjärde strecksatserna behöver inte iakttas vid förvärvstillfället, om bruttomängden av skuldförbindelserna eller av penningmarknadsinstrumenten eller nettomängden av de värdepapper som är föremål för emission då inte kan beräknas."
17. I artikel 25.3 a, b och c skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
18. Artikel 25.3 e skall ersättas med följande: "e) Ett eller flera investeringsbolags aktieinnehav i dotterbolag vars verksamhet enbart består i förvaltning, rådgivning eller saluföring i det land där dotterbolaget är beläget, vid återköp av andelar på begäran av andelsägarna, uteslutande för investeringsbolagets eller investeringsbolagens räkning."
19. Artikel 26.1 skall ersättas med följande: "1. Fondföretag behöver inte iaktta de gränsvärden som anges i detta avsnitt när de nyttjar teckningsrätter för överlåtbara värdepapper eller penningmarknadsinstrument som ingår i fondtillgångarna.
Medlemsstaterna får, med beaktande av principen om riskspridning, tillåta nyligen auktoriserade fondföretag att under en tid av högst sex månader från auktorisationsdagen avvika från artiklarna 22, 22a, 23 och 24."
20. Artikel 41.2 skall ersättas med följande: "2. Bestämmelserna i punkt 1 skall inte hindra sådana företag från att förvärva överlåtbara värdepapper, penningmarknadsinstrument eller andra finansiella instrument som avses i artikel 19.1 e, g och h och som inte är till fullo betalda."
22. Efter artikel 53 skall följande artikel läggas till: "Artikel 53a
1. Utöver de funktioner som finns angivna i artikel 53.1 kan kontaktkommittén också sammanträda som en föreskrivande kommitté i enlighet med artikel 5 i beslut 1999/468/EG(9) för att bistå kommissionen med tekniska ändringar i detta direktiv på följande områden:
- Förtydligande av definitionerna för att säkerställa en enhetlig tillämpning av detta direktiv inom hela gemenskapen.
- Likriktning av definitionerna i fråga om terminologi och utformning i enlighet med senare rättsakter avseende fondföretag och närstående frågor.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning.".
Artikel 2
1. Senast den 13 februari 2005 skall kommissionen lägga fram en rapport för rådet och Europaparlamentet om tillämpningen av det ändrade direktiv 85/611/EEG tillsammans med eventuella förslag till ändringar. Rapporten skall särskilt innehålla
a) en analys av hur man kan fördjupa och vidga den inre marknaden för fondföretag, särskilt vad gäller gränsöverskridande marknadsföring av fondföretag (även tredjemansfonder), hur passet för förvaltningsföretag fungerar, hur det förenklade prospektet fungerar som informations- och marknadsföringsverktyg, en översyn av omfattningen av tillhörande verksamhet samt möjligheterna till förbättrat samarbete mellan kontrollmyndigheter vad gäller enhetlig tolkning och tillämpning av direktivet,
b) en översyn av direktivets tillämpningsområde vad gäller olika produkttyper (till exempel institutionella fonder, fastighetsfonder, matarfonder och hedgefonder); översynen bör särskilt inriktas på storleken på marknaden för sådana fonder, eventuell reglering av sådana fonder i medlemsstaterna och bedömning av behovet av ytterligare harmonisering av dessa fonder,
c) en utvärdering av hur fonderna organiseras, inklusive bestämmelser och metoder för delegering samt förhållandet mellan fondförvaltare och förvaringsinstitut,
d) en översyn av investeringsbestämmelserna för fondföretag, till exempel användningen av derivatinstrument och andra instrument samt tekniker för värdepapper, reglering av indexfonder, reglering av penningmarknadsinstrument, inlåning, reglering av fond-till-fond-investeringar liksom de olika investeringsgränserna,
e) en analys av konkurrenssituationen mellan fonder som förvaltas av förvaltningsföretag respektive investeringsföretag som sköter förvaltningen själva.
När kommissionen utarbetar denna rapport skall den i största möjliga utsträckning samråda med de olika branschintressena samt med konsumentorganisationer och tillsynsorgan.
2. Medlemsstaterna får bevilja fondföretag, som är verksamma vid tidpunkten för detta direktivs ikraftträdande, en frist om högst 60 månader från denna tidpunkt för att de skall kunna anpassa sig till den nya nationella lagstiftningen.
Artikel 3
Medlemsstaterna skall anta de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 13 augusti 2003. De skall genast underrätta kommissionen om detta.
De skall börja tillämpa dessa åtgärder senast den 13 februari 2004.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 4
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 70/2001
av den 12 januari 2001
om tillämpningen av artiklarna 87 och 88 i EG-fördraget på statligt stöd till små och medelstora företag
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 994/98 av den 7 maj 1998 om tillämpningen av artiklarna 92 och 93 i Fördraget om upprättandet av Europeiska gemenskapen på vissa slag av övergripande statligt stöd(1), särskilt artikel 1 a i och 1 b i denna,
efter att ha offentliggjort ett utkast till denna förordning(2),
efter samråd med Rådgivande kommittén för statligt stöd, och
av följande skäl:
(1) Genom förordning (EG) nr 994/98 bemyndigas kommissionen att i enlighet med artikel 87 i fördraget förklara att stöd till små och medelstora företag på vissa villkor skall vara förenliga med den gemensamma marknaden och undantagna från anmälningsskyldigheten enligt artikel 88.3 i fördraget.
(2) Genom förordning (EG) nr 994/98 bemyndigas också kommissionen att i enlighet med artikel 87 i fördraget förklara att stöd som är förenliga med den av kommissionen för varje medlemsstat godkända regionalstödskartan är förenliga med den gemensamma marknaden och undantagna från anmälningsskyldigheten enligt artikel 88.3 i fördraget.
(3) Kommissionen har i ett stort antal beslut tillämpat artiklarna 87 och 88 i fördraget på små och medelstora företag både inom och utanför stödområden och har också redogjort för sin politik på området, senast i gemenskapens riktlinjer för statligt stöd till små och medelstora företag(3), och i riktlinjerna för statligt stöd för regionala ändamål(4). För att säkerställa effektiv kontroll och förenklad administration utan att kommissionens kontroll försvagas bör kommissionen, mot bakgrund av dels sin stora erfarenhet av att tillämpa dessa artiklar på små och medelstora företag, dels de allmänna texter om små och medelstora företag och regionalstöd som den antagit på grundval av dessa artiklar, göra bruk av sina befogenheter enligt förordning (EG) nr 994/98.
(4) Denna förordning påverkar inte medlemsstaternas möjligheter att anmäla stöd till små och medelstora företag. Sådana anmälningar kommer att bedömas av kommissionen särskilt utifrån kriterierna i denna förordning. Riktlinjerna för statligt stöd till små och medelstora företag bör upphävas den dag då denna förordning träder i kraft, eftersom deras innehåll förs in i den här förordningen.
(5) Små och medelstora företag spelar en avgörande roll för att skapa arbetstillfällen och medverkar allmänt till social stabilitet och en dynamisk ekonomi. Brister i marknadens sätt att fungera kan emellertid hämma deras utveckling. De har ofta svårigheter att få tillgång till kapital och krediter till följd av obenägenheten att ta risker på vissa finansiella marknader och de begränsade garantier som dessa företag kan erbjuda. De små och medelstora företagens begränsade resurser kan också inskränka deras möjligheter att få tillgång till information, särskilt om ny teknik och nya marknader. Mot bakgrund av dessa överväganden bör det stöd som genom denna förordning undantas från anmälningsskyldigheten syfta till att underlätta utvecklingen av verksamheten i de små och medelstora företagen, under förutsättning att stödet inte påverkar handeln i negativ riktning i en omfattning som strider mot det gemensamma intresset.
(6) Genom denna förordning bör undantag medges för alla stöd som uppfyller förordningens samtliga tillämpliga krav, och för alla stödordningar, förutsatt att varje stöd som kan beviljas inom ramen för dessa ordningar uppfyller samtliga tillämpliga krav enligt förordningen. För att säkerställa effektiv kontroll och förenklad administration utan att kommissionens kontroll försvagas bör stödordningar och enskilda stöd som inte omfattas av någon stödordning innehålla en uttrycklig hänvisning till denna förordning.
(7) Denna förordning bör inte påverka tillämpningen av särskilda regler i förordningar och direktiv om statligt stöd inom vissa sektorer, såsom de gällande reglerna för varvssektorn, och den bör inte vara tillämplig inom jordbruks- samt fiske- och vattenbrukssektorn.
(8) För att vid tillämpningen av denna förordning eliminera olikheter som kan medföra snedvridningar av konkurrensen och för att underlätta samordningen mellan olika initiativ inom gemenskapen och på nationell nivå som rör små och medelstora företag samt av hänsyn till administrativ klarhet och rättssäkerhet, bör definitionen av små och medelstora företag i denna förordning vara densamma som fastställs i kommissionens rekommendation 96/280/EG av den 3 april 1996 om definitionen av små och medelstora företag(5). Den definitionen används också i gemenskapens riktlinjer för statligt stöd till små och medelstora företag(6).
(9) För att bättre säkerställa att stödet är proportionellt och begränsas till det belopp som är nödvändigt, bör tröskelvärdena i enlighet med kommissionens fastlagda praxis uttryckas som stödnivåer i förhållande till stödberättigande kostnader snarare än som maximala stödbelopp.
(10) För att fastställa huruvida stöd som omfattas av denna förordning är förenliga med den gemensamma marknaden, är det nödvändigt att ta hänsyn till stödnivån och således stödbeloppet uttryckt i bidragsekvivalenter. Vid beräkningen av bidragsekvivalenten av stöd som kan betalas ut i flera omgångar och stöd i form av mjuka lån måste de marknadsräntor som rådde när stödet beviljades användas. För att säkerställa en enhetlig, öppen och enkel tillämpning av reglerna för statligt stöd, bör med marknadsräntor i denna förordning avses referensräntorna, under förutsättning att det ställs normala säkerheter när det gäller mjuka lån och att dessa inte innebär ett onormalt risktagande. Referensräntorna bör vara de räntor som löpande fastställs av kommissionen på grundval av objektiva kriterier och som offentliggörs i Europeiska gemenskapernas officiella tidning samt på Internet.
(11) Med hänsyn till skillnaderna mellan små företag och medelstora företag bör olika stödtak fastställas för små företag respektive medelstora företag.
(12) Enligt kommissionens erfarenhet bör stödtaken fastställas till en nivå som ger en balans mellan målsättningen att skapa minsta möjliga snedvridning av konkurrensen inom den understödda sektorn och målsättningen att underlätta de små och medelstora företagens ekonomiska utveckling.
(13) Det är lämpligt att fastställa ytterligare villkor som bör uppfyllas av varje stödordning eller enskilt stöd som beviljas undantag med stöd av denna förordning. Med hänvisning till artikel 87.3 c i fördraget bör sådana stöd normalt inte ha som enda syfte att fortlöpande eller periodiskt minska de driftskostnader som stödmottagaren normalt skall stå för, och de bör stå i proportion till de hinder som måste övervinnas för att uppnå de sociala och ekonomiska fördelar som anses vara i gemenskapens intresse. Tillämpningsområdet för denna förordning bör därför begränsas till stöd som ges till vissa materiella och immateriella investeringar, vissa tjänster som tillhandahålls stödmottagarna och viss övrig verksamhet. Mot bakgrund av den överkapacitet inom transportsektorn som råder i gemenskapen, med undantag för rullande järnvägsmateriel, bör transportmedel och transportutrustning inte ingå i de stödberättigande investeringskostnaderna för företag som har sin huvudsakliga ekonomiska verksamhet inom transportsektorn.
(14) Genom denna förordning bör stöd till små och medelstora företag undantas från anmälningsskyldigheten oberoende av var företagen är belägna. Investeringar och skapande av arbetstillfällen kan bidra till den ekonomiska utvecklingen i gemenskapens mindre gynnade regioner. Små och medelstora företag i dessa regioner har strukturella nackdelar på grund av sin lokalisering och svårigheter på grund av sin begränsade storlek. De bör därför beviljas högre stödtak.
(15) För att inte gynna kapitalfaktorn på bekostnad av arbetsfaktorn i samband med en investering, bör i denna förordning föreskrivas en möjlighet att mäta investeringsstöd på grundval av antingen investeringskostnader eller kostnader för nyanställningar i samband med att ett investeringsprojekt genomförs.
(16) Mot bakgrund av Världshandelsorganisationens (WTO) avtal om subventioner och kompensatoriska åtgärder(7) bör exportstöd och stöd som gynnar inhemska produkter på bekostnad av importerade produkter inte undantas enligt denna förordning. Bidrag till kostnaderna för deltagande i handelsmässor eller för undersökningar eller konsulttjänster som behövs för att lansera en ny produkt eller en befintlig produkt på en ny marknad utgör normalt inte exportstöd.
(17) Med hänsyn till behovet att uppnå balans mellan minsta möjliga snedvridning av konkurrensen inom den understödda sektorn och denna förordnings mål bör enskilda stöd som överskrider ett fastställt maximibelopp inte medges undantag enligt denna förordning, oavsett om de omfattas av en stödordning som har beviljats undantag enligt denna förordning eller inte.
(18) För att säkerställa att stödet är nödvändigt och fungerar som ett incitament för att utveckla en viss verksamhet bör undantag enligt denna förordning inte beviljas för verksamhet som stödmottagaren även skulle bedriva på rena marknadsvillkor.
(19) Undantag bör enligt denna förordning inte medges stöd som kumuleras med annat statligt stöd, inbegripet stöd från nationella, regionala eller lokala myndigheter, eller med gemenskapsbidrag, om, i förhållande till samma stödberättigande kostnader, ett sådant kumulerat stöd, överstiger de tröskelvärden som anges i denna förordning.
(20) I syfte att säkerställa insyn och effektiv kontroll i enlighet med artikel 3 i förordning (EG) nr 994/98 är det lämpligt att utarbeta ett standardformulär som medlemsstaterna bör använda för att förse kommissionen med sammanfattande information för offentliggörande i Europeiska gemenskapernas officiella tidning, varje gång en stödordning genomförs eller ett enskilt stöd som inte täcks av någon sådan stödordning beviljas enligt denna förordning. Av samma skäl är det lämpligt att fastställa regler för de register som medlemsstaterna bör föra över stöd som har beviljats undantag enligt denna förordning. Beträffande den årliga rapport som medlemsstaterna är skyldiga att överlämna till kommissionen, är det lämpligt att kommissionen fastställer de närmare kraven på rapportens utformning, inbegripet information i elektronisk form, då den teknik som krävs för detta är allmänt tillgänglig.
(21) Med hänsyn till kommissionens erfarenhet på detta område, särskilt av hur ofta det i allmänhet är nödvändigt att se över politiken på området för statligt stöd, bör tillämpningsperioden för denna förordning begränsas. Om denna förordnings giltighetstid skulle löpa ut utan att förlängas, bör stödordningar som redan undantagits enligt denna förordning fortsätta att vara undantagna i sex månader.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Tillämpningsområde
1. Denna förordning gäller för statligt stöd som beviljas små och medelstora företag inom alla sektorer, utan att det påverkar tillämpningen av särskilda gemenskapsförordningar eller gemenskapsdirektiv enligt EG-fördraget vilka styr beviljandet av statligt stöd till särskilda sektorer, oavsett om de är mer eller mindre restriktiva än denna förordning.
2. Denna förordning får inte tillämpas på
a) verksamheter i samband med produktion, bearbetning eller marknadsföring av de produkter som förtecknas i bilaga I till fördraget,
b) exportrelaterade stöd, d.v.s. stöd som är direkt knutna till exporterade volymer, till upprättandet eller driften av ett distributionsnät eller till andra löpande uppgifter som har samband med exportverksamhet,
c) stöd som förutsätter att inhemska produkter används på bekostnad av importerade produkter.
Artikel 2
Definitioner
I denna förordning används följande beteckningar med de betydelser som här anges:
a) stöd: varje åtgärd som uppfyller samtliga kriterier som anges i artikel 87.1 i fördraget.
b) små och medelstora företag: företag som definieras i bilaga I.
c) investering i materiella tillgångar: investering i materiella anläggningstillgångar som hänför sig till skapandet av en ny anläggning, utvidgning av en existerande anläggning, eller igångsättande av en verksamhet som innebär en grundläggande förändring av en existerande anläggningsprodukt eller produktionsprocess (genom rationalisering, omställning eller modernisering). En investering i anläggningstillgångar som genomförs i form av övertagande av en anläggning som har lagts ned eller som skulle ha lagts ned om den inte hade förvärvats skall också betraktas som en materiell investering.
d) investering i immateriella tillgångar: investering i överföring av teknik genom förvärv av patenträttigheter, licenser, know-how eller icke patentskyddad teknisk kunskap.
e) stödnivå brutto: stödbeloppet uttryckt i procent av projektets stödberättigande kostnader. Alla siffror som används skall avse belopp före eventuella avdrag för direkt skatt. Om stöd beviljas i någon annan form än som bidrag, skall stödbeloppet vara lika med stödets bidragsekvivalent. Stöd som betalas ut i flera omgångar skall aktualiseras till sitt värde vid tidpunkten för beviljandet. Den ränta som skall användas för nuvärdesberäkningar och för att räkna ut stödbeloppet i ett mjukt lån skall vara den gällande referensräntan vid den tidpunkt då lånet beviljades.
f) stödnivå netto: stödbeloppet efter avdrag för skatt i procent av projektets stödberättigande kostnader.
g) antal anställda: antalet arbetskraftsenheter per år, dvs. antalet heltidsanställda under ett år, medan deltidsarbete eller säsongsarbete utgör delar av arbetskraftsenheter.
Artikel 3
Förutsättningar för undantag
1. Enskilda stöd som inte omfattas av någon stödordning och som uppfyller samtliga villkor enligt denna förordning skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget, under förutsättning att stöden innehåller en uttrycklig hänvisning till denna förordning, med angivande av förordningens titel och en hänvisning till dess offentliggörande i Europeiska gemenskapernas officiella tidning.
2. Stödordningar som uppfyller samtliga villkor enligt denna förordning skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget, under förutsättning att
a) varje stöd som skulle kunna beviljas inom ramen för stödordningen uppfyller samtliga villkor i denna förordning,
b) stödordningen innehåller en uttrycklig hänvisning till denna förordning, med angivande av förordningens titel och en hänvisning till dess offentliggörande i Europeiska gemenskapernas officiella tidning.
3. Stöd som beviljas enligt en sådan stödordning som avses i punkt 2 skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget, under förutsättning att det beviljade stödet direkt uppfyller samtliga villkor i denna förordning.
Artikel 4
Investeringar
1. Stöd till investeringar i materiella och immateriella tillgångar inom och utom gemenskapen skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskraven i artikel 88.3 i fördraget om det uppfyller villkoren i punkterna 2-6.
2. Stödnivån brutto får inte överskrida
a) 15 % för små företag, eller
b) 7,5 % för medelstora företag.
3. Om investeringen äger rum i områden som är berättigade till regionalstöd får stödnivån inte överstiga det tak för regionalt investeringsstöd som fastställts i den karta som kommissionen har godkänt för varje medlemsstat med mer än
a) 10 procentenheter brutto i de områden som omfattas av artikel 87.3 c, under förutsättning att den totala stödnivån netto inte överstiger 30 %, eller
b) 15 procentenheter brutto i de områden som omfattas av artikel 87.3 a, under förutsättning att den totala stödnivån netto inte överstiger 75 %.
De högre regionala stödtaken skall endast gälla om stödet beviljas på villkor att investeringen bibehålls i den stödmottagande regionen under minst fem år och att stödmottagarens bidrag till finansieringen av investeringen uppgår till minst 25 %.
4. De tak som fastställs i punkterna 2 och 3 skall gälla stödnivån beräknad antingen som en procentandel av investeringens stödberättigande kostnader eller som en procentandel av lönekostnaden för den sysselsättning som skapas till följd av investeringen (stöd till skapande av arbetstillfällen) eller en kombination av båda, under förutsättning att stödet inte överstiger det högsta belopp som endera av beräkningssätten resulterar i.
5. Om stödet beräknas på grundval av investeringskostnaderna, skall de stödberättigande kostnaderna för materiella investeringar utgöra kostnader som avser investeringar i mark, byggnader, maskiner och utrustning. Inom transportsektorn får, med undantag för rullande järnvägsmateriel, transportmedel och transportutrustning inte ingå i de stödberättigande kostnaderna. Stödberättigande kostnader för immateriella investeringar skall vara kostnader för förvärv av teknologi.
6. Om stödet beräknas på grundval av skapade arbetstillfällen skall stödbeloppet uttryckas i procent av lönekostnaderna för den sysselsättning som skapats under en tvåårsperiod enligt följande villkor:
a) Den skapade sysselsättningen måste ha samband med genomförandet av ett investeringsprojekt i materiella eller immateriella tillgångar. Arbetstillfällena måste skapas inom tre år från det att investeringen har slutförts.
b) Investeringsprojektet måste leda till en nettoökning av antalet sysselsatta i den berörda anläggningen i förhållande till det genomsnittliga antalet anställda under de senaste tolv månaderna.
c) Den skapade sysselsättningen måste bibehållas under en period av minst fem år.
Artikel 5
Rådgivningsverksamhet och andra tjänster och verksamheter
Stöd till små och medelstora företag som uppfyller följande villkor skall vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget:
a) För tjänster som tillhandahålls av utomstående konsulter får stödet brutto inte överstiga 50 % av kostnaderna för dessa tjänster. De berörda tjänsterna får varken vara av fortlöpande eller periodiskt slag eller röra företagets ordinarie driftsutgifter, som t.ex. rutinmässig skatterådgivning, regelbunden juridisk rådgivning eller annonskostnader.
b) För deltagande i mässor och utställningar får stödet brutto inte överstiga 50 % av merkostnaderna för hyra, uppförande och drift av utställningsmontern. Detta undantag skall endast gälla för ett företags första deltagande i en viss mässa eller utställning.
Artikel 6
Beviljande av stora enskilda stöd
Ett enskilt stöd som uppfyller ett av följande tröskelvärden får inte beviljas undantag enligt denna förordning:
a) de totala stödberättigande kostnaderna för hela projektet är minst 25 miljoner euro, och
i) stödnivån brutto i områden som inte är berättigade till regionalstöd är minst 50 % av de stödnivåer som anges i artikel 4.2,
ii) stödnivån netto i områden som är berättigade till regionalstöd är minst 50 % av stödtaket netto enligt regionalstödskartan för området i fråga, eller
b) det totala stödbeloppet brutto är minst 15 miljoner euro.
Artikel 7
Villkor för stödet
Stöd får beviljas undantag enligt denna förordning endast om medlemsstaten innan arbetet på det berörda projektet inleds
- har fått en ansökan om stöd från stödmottagaren, eller
- har antagit bestämmelser som fastställer en laglig rätt till stöd enligt objektiva kriterier och utan vidare diskretionär prövningsrätt för medlemsstaten
Artikel 8
Kumulering
1. De stödtak som fastställs i artiklarna 4, 5 och 6 skall tillämpas oavsett om stödet helt finansieras med statliga medel eller samfinansieras av gemenskapen.
2. Stöd som undantas genom denna förordning får inte kumuleras med något annat statligt stöd i den mening som avses i artikel 87.1 i fördraget eller med annan gemenskapsfinansiering, i förhållande till samma stödberättigande kostnader, om en sådan kumulering skulle leda till en högre stödnivå än den som fastställs i denna förordning.
Artikel 9
Insyn och kontroll
1. Vid genomförandet av en stödordning eller vid beviljandet av ett enskilt stöd som inte omfattas av någon stödordning, skall medlemsstaterna, om stödordningen eller stödet är undantaget enligt denna förordning, till kommissionen inom tjugo arbetsdagar överlämna en sammanfattning av uppgifterna om stödordningen eller det enskilda stödet enligt det formulär som anges i bilaga II för offentliggörande i Europeiska gemenskapernas officiella tidning.
2. Medlemsstaterna skall föra detaljerade register över de stödordningar som undantas genom denna förordning, de enskilda stöd som beviljas enligt dessa stödordningar, och de enskilda stöd som undantas enligt denna förordning och som beviljas vid sidan om en befintlig stödordning. Dessa register skall innehålla alla uppgifter som behövs för att det skall vara möjligt att fastställa att de villkor för beviljande av undantag som anges i denna förordning har uppfyllts inbegripet uppgifter om företagets status som litet eller medelstort företag. Medlemsstaterna skall bevara ett register över ett enskilt stöd under tio år från den dag då stödet beviljades, och, när det gäller en stödordning, under tio år från den dag då det sista enskilda stödet beviljades enligt stödordningen. En berörd medlemsstat skall på skriftlig begäran inom tjugo arbetsdagar, eller inom en längre tidsfrist som anges i begäran, förse kommissionen med alla uppgifter den anser sig behöva för att kunna bedöma om villkoren i denna förordning har följts.
3. Medlemsstaterna skall sammanställa en rapport om tillämpningen av denna förordning för varje helt kalenderår eller del av kalenderår under vilket denna förordning gäller, enligt den förlaga som anges i bilaga III och även i elektronisk form. Medlemsstaterna skall överlämna en sådan rapport till kommissionen senast tre månader efter utgången av den period som rapporten avser.
Artikel 10
Ikraftträdande och giltighetstid
1. Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 283/2001
av den 9 februari 2001
om ändring av förordning (EG) nr 562/2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 1254/1999 vad avser systemen för offentliga interventionsuppköp inom nötköttssektorn och förordning (EG) nr 2734/2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1254/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för nötkött(1), särskilt artikel 47.8 i denna, och
av följande skäl:
(1) Genom kommissionens förordning (EG) nr 2734/2000 av den 14 december 2000 om ändring av förordning (EEG) nr 1627/89 om uppköp av nötkött genom anbudsinfordran och om undantag från eller ändring av förordning (EG) nr 562/2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 1254/1999 vad avser systemen för offentliga interventionsuppköp inom nötköttssektorn(2), ändrad genom förordning (EG) nr 3/2001(3), fastställdes ett antal ändringar av eller undantag från kommissionens förordning (EG) nr 562/2000(4) med anledning av den exceptionella situationen på marknaden till följd av den senaste händelseutvecklingen i samband med bovin spongiform encefalopati (BSE).
(2) Med hänsyn till den exceptionella situationen på marknaden och för att de interventionsåtgärder som föreskrivs i förordning (EG) nr 2734/2000 skall ha större effekt bör det medges undantag från artikel 4.2 g i förordning (EG) nr 562/2000 vad gäller den maximala vikten för slaktkroppar genom att inte fastställa någon viktbegränsning för de två anbudsförfarandena under februari månad och genom att öka vikten till 430 kg för de resterande anbudsförfarandena under det första kvartalet 2001 och samtidigt tillåta uppköp av tyngre djur, men då begränsa priset för dessa till det pris som betalas för den högsta tillåtna vikten.
(3) Följaktligen bör förordning (EG) nr 2734/2000 ändras.
(4) Med hänsyn till att produkter som köps upp för intervention även får säljas efter den 1 januari 2002, när det obligatoriska märkningssystemet enligt Europaparlamentets och rådets förordning av den 17 juli 2000 om upprättande av ett system för identifiering och registrering av nötkreatur samt märkning av nötkött och nötköttsprodukter och om upphävande av rådets förordning (EG) nr 820/97(5) skall börja tillämpas, bör det för avtal som sluts från och med den 12 februari, dvs. från och med februari månads första anbudsförfarande, vara obligatoriskt att i märkningen ange det eller de länder där de berörda djuren är födda eller har fötts upp enligt artikel 13.5 i förordning (EG) nr 1760/2000, och i förekommande fall de uppgifter som föreskrivs i artikel 2.2 i kommissionens förordning 1825/2000 om tillämpningsföreskrifter för Europaparlamentets och rådets förordning (EG) nr 1760/2000(6).
(5) I bilaga III till förordning (EG) nr 562/2000 fastställs de bestämmelser som hela och halva slaktkroppar samt kvartsparter måste följa om de skall få köpas upp för offentlig intervention. För att anpassa bestämmelserna till gällande handelssed bör beskrivningen av halva slaktkroppar i den bilagan ändras så att den tillåter viss variation.
(6) Följaktligen bör förordning (EG) nr 562/2000 ändras.
(7) Med hänsyn till händelseutvecklingen bör denna förordning träda i kraft omedelbart.
(8) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för nötkött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 6.1 i förordning (EG) nr 2734/2000 skall ersättas med följande:
"1. Trots vad som sägs i artikel 4.2 g i förordning (EG) nr 562/2000 skall den maximala vikten för de slaktkroppar som avses i ovannämnda bestämmelse vara 430 kg. Dock
- skall ingen begränsning av den maximala vikten för slaktkroppar tillämpas för de två anbudsförfarandena i februari månad.
- får slaktkroppar med en vikt över 430 kg köpas för intervention vid de resterande anbudsförfarandena under det första kvartalet 2001, men i sådana fall skall uppköpspriset högst vara det som betalas för den maximala vikten."
Artikel 2
Förordning (EG) nr 562/2000 ändras på följande sätt:
1. Artikel 4.3 d skall ersättas med följande:
"d) De har försetts med etiketter i enlighet med det system som införs genom Europaparlamentets och rådets förordning (EG) nr 1760/2000(7), samt för avtal som sluts från och med den 12 februari 2001 även de uppgifter som anges i artikel 13.5 i den förordningen."
2. I bilaga III skall punkt 2 b ersättas med följande:
"b) halv slaktkropp: de produkter som erhålls genom symmetrisk delning av den slaktkropp som avses i a ovan genom mitten av hals-, rygg-, länd- och korskotorna och genom mitten av bröstbenet och bäckenbensfogen. Under uppslaktning och hantering av slaktkroppen får inte rygg- och ländkotorna tydligt förskjutas. Tillhörande muskler och senor får inte skadas allvarligt av såg eller kniv."
Artikel 3
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 749/2001
av den 18 april 2001
om ändring av bilaga II till rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), senast ändrad genom kommissionens förordning (EG) nr 2908/2000(2), särskilt artiklarna 7 och 8 i denna, och
av följande skäl:
(1) I enlighet med förordning (EEG) nr 2377/90 måste gränsvärden för högsta tillåtna restmängder successivt fastställas för samtliga farmakologiskt verksamma substanser som används inom gemenskapen veterinärmedicinska läkemedel som är avsedda att ges till livsmedelsproducerande djur.
(2) Gränsvärden bör fastställas först efter det att Kommittén för veterinärmedicinska läkemedel har granskat all relevant information beträffande säkerheten med restmängder av ämnet i fråga för den som konsumerar livsmedel med animaliskt ursprung samt restmängdernas påverkan på den industriella bearbetningen av livsmedel.
(3) Vid fastställandet av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung är det nödvändigt att ange de djurarter i vilka restmängder kan förekomma, vilka mängder som kan förekomma i var och en av de relevanta vävnaderna från det behandlade djuret (målvävnad) samt vilket slag av restmängd som är relevant vid övervakningen av restmängder (restmarkör).
(4) För kontroll av resthalter bör enligt tillämplig gemenskapslagstiftning gränsvärden vanligtvis fastställas för målvävnaderna lever eller njure. I den internationella handeln avlägsnas dock ofta lever och njure från slaktkroppen, och gränsvärden bör därför alltid fastställas även för muskel- eller fettvävnader.
(5) För veterinärmedicinska läkemedel som är avsedda för äggläggande fåglar, mjölkdjur eller honungsbin, måste gränsvärden även fastställas för ägg, mjölk eller honung.
(6) Tiamylal och Tiopentalnatrium skall införas i bilaga II till förordning (EEG) nr 2377/90.
(7) En tillräckligt lång tidsfrist bör fastställas innan denna förordning träder i kraft så att medlemsstaterna kan göra de nödvändiga anpassningarna till bestämmelserna i denna förordning av tillstånden att släppa ut de berörda veterinärmedicinska läkemedlen på marknaden, vilka beviljats enligt rådets direktiv 81/851/EEG(3), senast ändrat genom kommissionens direktiv 2000/37/EG(4).
(8) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga II till förordning (EEG) nr 2377/90 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 939/2001
av den 14 maj 2001
om tillämpningsföreskrifter till rådets förordning (EG) nr 104/2000 beträffande beviljande av schablonmässigt stöd för vissa fiskeriprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 104/2000 av den 17 december 1999 om den gemensamma organisationen av marknaden för fiskeri- och vattenbruksprodukter(1), särskilt artikel 24.8 i denna, och
av följande skäl:
(1) I artikel 24 i förordning (EG) nr 104/2000, som upphävde rådets förordning (EEG) nr 3759/92(2) med verkan från och med den 1 januari 2001, föreskrivs att ett schablonmässigt stöd på vissa villkor skall beviljas producentorganisationer som återtar produkter som förtecknas i bilaga IV till den förordningen.
(2) I syfte att harmonisera och förenkla bör de förfaranden som krävs inom ramen för det schablonmässiga stödet vara analoga med dem som gäller för den ekonomiska ersättningen och förädlingsstödet, såsom följer av kommissionens förordning (EG) nr 2509/2000 av den 15 november 2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 104/2000 beträffande beviljande av ekonomisk ersättning för återtag från marknaden av vissa fiskeriprodukter(3), och kommissionens förordning (EG) nr 2814/2000 av den 21 december 2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 104/2000 beträffande beviljande av förädlingsstöd för vissa fiskeriprodukter(4). Villkoren för att bevilja schablonmässigt stöd bör följaktligen fastställas på denna grund och kommissionens förordning (EG) nr 4176/88 av den 28 december 1988 om tillämpningsföreskrifter för beviljande av fast stöd för vissa fiskeri- och vattenbruksprodukter(5), senast ändrad genom förordning (EG) nr 3516/93(6), bör upphöra att gälla.
(3) I artikel 6.1 i rådets förordning (EG) nr 2406/96 av den 26 november 1996 om fastställande av gemensamma marknadsnormer för saluföring av vissa fiskeriprodukter(7), senast ändrad genom förordning (EG) nr 2578/2000(8), föreskrivs att produkter i kategori B inte skall berättiga till ekonomiskt stöd i samband med intervention inom ramen för den gemensamma organisationen av marknaden. I den mån som endast produkter av kvalitet Extra, "E" och "A" berättigar till schablonmässigt stöd enligt artikel 24 i förordning (EG) nr 104/2000, bör beräkningen av stödberättigande kvantiteter uteslutande göras på grundval av dessa produktkategorier.
(4) Det bör fastställas bestämmelser som producentorganisationerna skall följa när det gäller schablonmässigt stöd.
(5) Det schablonmässiga stödet får betalas ut först efter fiskeårets slut. Det bör emellertid införas en möjlighet att bevilja förskott, förutsatt att säkerhet ställs.
(6) För beräkningen av det schablonmässiga stödet bör medlemsstaterna tillåtas att fastställa ett schablonvärde, fördelat på de återtagna produkternas avsättning enligt kommissionens förordning (EEG) nr 1501/83 av den 9 juni 1983 om omhändertagande av vissa fiskeriprodukter som varit föremål för marknadsstabiliserande åtgärder(9), ändrad genom förordning (EEG) nr 1106/90(10).
(7) För att säkerställa produkternas kvalitet och underlätta deras avsättning på marknaden bör det fastställas vilka minimikrav för beredningen som skall vara tillgodosedda och vilka villkor som skall gälla för lagring och återförande till marknaden av de bearbetade produkterna.
(8) Stödmottagarna bör föra lagerbokföring (i kg) över de varor som varje månad bjuds ut till försäljning, återtas och förädlas för att effektiviteten i kontrollerna skall kunna ökas och de bör meddela dessa uppgifter till medlemsstaten. För ett väl fungerande system är det tillräckligt att kräva lagerbokföring under den kortast tillåtna lagringsperioden.
(9) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fiskeriprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
Allmänna villkor
Artikel 1
Artikel 2
Det schablonmässiga stödet skall betalas ut till den berörda producentorganisationen först sedan medlemsstatens behöriga myndighet har konstaterat att de kvantiteter för vilka stödet har sökts inte överstiger den högsta nivå som anges i artikel 24.5 i förordning (EG) nr 104/2000.
KAPITEL II
Villkor för att bevilja schablonmässigt stöd enligt artikel 24.2 i förordning (EG) nr 104/2000 (nedan kallat schablonersättning)
Artikel 3
Villkoren i artiklarna 1-4 och artikel 7 i förordning (EG) nr 2509/2000 skall i tillämpliga delar gälla för beviljande av schablonersättning.
Artikel 4
Medlemsstaterna skall fastställa ett schablonvärde för att beräkna schablonersättning och tillhörande förskott, fördelat på de återtagna produkternas avsättning enligt artikel 1 b, c och d i förordning (EEG) nr 1501/83.
För alla producentorganisationer som medlemsstaten har erkänt skall det fastställas ett schablonvärde vid fiskeårets början på grundval av de genomsnittliga inkomster som i samband med dessa avsättningar uppnåtts och konstaterats i de berörda medlemsstaterna under sex månader innan detta schablonvärde fastställs. Värdet skall emellertid ändras om väsentliga och bestående inkomstvariationer konstateras på medlemsstatens marknad.
KAPITEL III
Villkor för att bevilja schablonmässigt stöd enligt artikel 24.4 i förordning (EG) nr 104/2000 (nedan kallat schablonbidrag)
Artikel 5
1. Schablonbidraget skall fastställas innan fiskeåret börjar enligt artikel 38.2 i förordning (EG) nr 104/2000. Beloppet skall fastställas per viktenhet och gälla för nettovikten av de produkter som anges i bilaga IV till förordning (EG) nr 104/2000.
2. Schablonbidraget skall beräknas på grundval av de faktiska tekniska och ekonomiska kostnader för nödvändiga åtgärder vid stabiliseringsbehandling och lagring av produkterna i fråga som noterats i gemenskapen under det föregående fiskeåret.
3. Följande skall betraktas som tekniska kostnader:
a) Kostnader för energi.
b) Arbetskostnader i samband med lagring och uttag från lager.
c) Kostnader för material vid direktförpackning.
d) Beredningskostnader (ingredienser).
e) Transportkostnader från landningsställe till plats där beredningen sker.
4. De ekonomiska kostnaderna skall utgöras av ett schablonbelopp på 10 euro per ton för 2001. Därefter skall schablonbeloppet justeras årligen enligt den räntesats som årligen fastställs i enlighet med artikel 5 i rådets förordning (EEG) nr 1883/78(11).
5. Det schablonbidrag som fastställs för ett fiskeår skall gälla för produkter som började lagras under det året, oavsett när lagringen upphör.
Artikel 6
Bestämmelserna i artikel 3.1 och 3.2 samt artikel 4 i förordning (EG) nr 2814/2000 skall i tillämpliga delar gälla för beviljande av schablonbidrag.
Artikel 7
Schablonbidraget skall betalas ut till den berörda producentorganisationen först sedan medlemsstatens behöriga myndighet har konstaterat att de kvantiteter för vilka bidraget har sökts antingen beretts och lagrats eller konserverats och sedan återförts till marknaden i enlighet med bestämmelserna i artikel 4 i förordning (EG) nr 2814/2000.
KAPITEL IV
Slutbestämmelser
Artikel 8
1. Ansökningar om utbetalning av schablonmässigt stöd skall av producentorganisationerna överlämnas till de behöriga myndigheterna i medlemsstaten inom fyra månader från det aktuella fiskeårets slut. Ansökningarna skall minst innehålla de uppgifter som anges i bilagan.
2. Efter ansökan av en berörd producentorganisation skall förskott beviljas varje månad för återtagna eller förädlade kvantiteter, under förutsättning att producentorganisationen ställer en säkerhet som minst motsvarar 105 % av förskottsbeloppet.
3. Förskotten skall fastställas på grundval av det under perioden rådande preliminära förhållandet mellan återtagna och saluförda kvantiteter. Beräkningen av beloppet skall justeras två månader efter den aktuella månaden på grundval av de transaktioner som faktiskt genomförts och skall redovisas enligt den förlaga som finns i bilagan.
4. De nationella myndigheterna skall betala ut det schablonmässiga stödet senast åtta månader efter fiskeårets slut. Varje medlemsstat skall underrätta övriga medlemsstater och kommissionen om namn på och adress till det organ som utsetts att betala ut det schablonmässiga stödet.
Artikel 9
1. Medlemsstaterna skall införa en ordning för att kontrollera att den information som lämnas i ansökningarna om utbetalning överensstämmer med de kvantiteter som producentorganisationen i fråga faktiskt har salufört och återtagit från marknaden.
2. Producentorganisationerna skall se till att stödmottagarna för lagerbokföring i enlighet med den förlaga som finns i bilagan.
3. Producentorganisationen skall i fråga om de produkter som återtagits eller förädlats varje månad underrätta medlemsstaten om datum, art och kvantitet.
Artikel 10
Medlemsstaterna skall underrätta kommissionen om de åtgärder som vidtagits för tillämpningen av den här förordningen så snart de antagits, och i vart fall senast den 1 juli 2001. De skall senast den 1 juli 2001 underrätta kommissionen om redan gällande åtgärder på det område som omfattas av artikel 9.1.
Artikel 11
Förordning (EEG) nr 4176/88 skall upphöra att gälla.
Artikel 12
Europaparlamentets och rådets förordning (EG) nr 999/2001
av den 22 maj 2001
om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 152.4 b i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Flera olika typer av transmissibel spongiform encefalopati (TSE) har sedan flera år tillbaka konstaterats oberoende av varandra hos människor och djur. Bovin spongiform encefalopati (BSE) upptäcktes först hos nötkreatur 1986 och under följande år också hos andra djurarter. En ny variant av Creutzfeldt-Jakobs sjukdom (CJS) beskrevs 1996. Det samlas ständigt nya bevis för likheten mellan BSE-smittämnet och det smittämne som förorsakar den nya varianten av Creutzfeldt-Jakobs sjukdom.
(2) Sedan 1990 har gemenskapen beslutat om en rad åtgärder för att skydda människor och djur mot BSE-risken. Dessa åtgärder grundar sig på skyddsbestämmelserna i direktiven om kontrollåtgärder på veterinärområdet. Med hänsyn till omfattningen av den hälsorisk som människor och djur utsätts för genom vissa typer av TSE är det lämpligt att anta särskilda bestämmelser om förebyggande, kontroll och utrotning av dessa.
(3) Denna förordning har direkt avseende på folkhälsan och har betydelse för hur den inre marknaden fungerar. Den omfattar produkter som ingår i bilaga I till fördraget men även produkter som inte ingår i denna bilaga. Det är därför lämpligt att välja artikel 152.4 b i fördraget som rättslig grund.
(4) Kommissionen har erhållit vetenskapliga yttranden om flera aspekter av TSE, bland annat från Vetenskapliga styrkommittén och Vetenskapliga kommittén för veterinära åtgärder till skydd för människors hälsa. Vissa av dessa yttranden avser åtgärder för att minska den potentiella risken för att människor och djur skall utsättas för produkter från infekterade djur.
(5) Dessa bestämmelser bör gälla produktion och avyttring av levande djur och animaliska produkter. De behöver däremot inte gälla kosmetiska eller medicinska produkter, medicintekniska produkter, deras utgångsmaterial eller mellanprodukter, för vilka andra särskilda bestämmelser gäller, särskilt avseende förbud mot användning av vissa typer av riskmaterial. De bör inte heller gälla animaliska produkter som inte innebär någon hälsorisk för människor och djur eftersom de är avsedda att användas till annat än livsmedel, foder eller gödningsmedel. Det är däremot nödvändigt att säkerställa att animaliska produkter som inte omfattas av denna förordning hålls åtskilda från dem som omfattas av förordningen, om de inte uppfyller minst samma hälsovillkor som de sistnämnda.
(6) Det bör införas bestämmelser om att kommissionen får vidta skyddsåtgärder om den behöriga myndigheten i en medlemsstat eller i ett tredje land inte har hanterat TSE-risken på lämpligt sätt.
(7) Ett förfarande bör fastställas för att bestämma den epidemiologiska statusen för en medlemsstat, ett tredje land och en av dess regioner (nedan kallade länder eller regioner) med hänsyn till BSE på grundval av en bedömning av risken för förekomst (på engelska: incident risk), spridning och risk för att människor utsätts för smitta, utifrån tillgänglig information. Medlemsstater och tredje land som väljer att inte ansöka om att få sin status fastställd bör av kommissionen placeras i en kategori, på grundval av all information som kommissionen har tillgång till.
(8) Medlemsstaterna bör införa utbildningsprogram för dem som har till uppgift att förebygga och bekämpa TSE, liksom för veterinärer, jordbrukare och personer som har hand om transport, avyttring och slakt av livsmedelsproducerande djur.
(9) Medlemsstaterna måste årligen genomföra ett övervakningsprogram för BSE och scrapie och meddela kommissionen och de övriga medlemsstaterna resultaten härav samt om någon annan form av TSE har uppträtt.
(10) Vissa vävnader från idisslare bör betecknas som specificerat riskmaterial på grundval av de olika TSE-typernas patogener och den epidemiologiska statusen för det land eller den region där det berörda djuret har sitt ursprung eller sin hemvist. De specificerade riskmaterialen måste avlägsnas och destrueras på ett sådant sätt att människor och djur inte utsätts för några hälsorisker. Framför allt bör de inte avyttras för att användas vid tillverkning av livsmedel, foder eller gödningsmedel. Bestämmelser bör emellertid införas om möjlighet att uppnå en likvärdig hälsoskyddsnivå, med hjälp av ett TSE-test som utförs på enskilda djur, sedan full validitet fastställts. Slakttekniker som innebär en risk för att material från hjärnan infekterar andra vävnader bör inte tillåtas i andra länder eller regioner än de där BSE-risken är lägst.
(11) Åtgärder bör vidtas för att förhindra att TSE överförs till människor och djur genom förbud mot att utfodra vissa kategorier djur med vissa kategorier djurprotein, samt genom förbud mot att använda vissa material från idisslare i livsmedel. Dessa förbud bör stå i proportion till de risker det handlar om.
(12) Det bör föreskrivas att varje misstanke om någon form av TSE hos något djur skall anmälas till den behöriga myndigheten, som omedelbart skall vidta alla lämpliga åtgärder, och i synnerhet fastställa restriktioner för förflyttning av det misstänkta djuret i väntan på resultatet av undersökningen eller låta slakta det under officiell övervakning. Om den behöriga myndigheten inte kan utesluta möjligheten att djuret är smittat med TSE, bör den se till att lämpliga undersökningar görs och hålla slaktkroppen under officiell övervakning till dess att en diagnos har ställts.
(13) Om förekomst av TSE bekräftas officiellt, bör den behöriga myndigheten vidta alla nödvändiga åtgärder, i synnerhet låta destruera slaktkroppen, och genomföra en undersökning för att identifiera alla riskdjur och fastställa restriktioner för förflyttning av djur och animaliska produkter för vilka smittorisk konstaterats. Ägarna bör utan dröjsmål ersättas för förlust av djur och animaliska produkter som destruerats enligt denna förordning.
(14) Medlemsstaterna bör upprätta beredskapsplaner i vilka de nationella åtgärder som skall vidtas vid ett utbrott av BSE anges. Beredskapsplanerna bör godkännas av kommissionen. Bestämmelser bör införas för att kunna utsträcka denna bestämmelse till att gälla andra typer av TSE än BSE.
(15) Det bör fastställas bestämmelser om avyttring av vissa levande djur och animaliska produkter. I nuvarande gemenskapslagstiftning om identifiering och registrering av nötkreatur finns bestämmelser om ett system som gör det möjligt att, enligt internationella normer, spåra djuren tillbaka till moderdjuret och ursprungsbesättningen. Det bör införas bestämmelser om likvärdiga garantier i fråga om nötkreatur som importeras från tredje land. Djur och animaliska produkter som omfattas av nämnda lagstiftning och som förflyttas vid handel inom gemenskapen eller importeras från tredje land bör åtföljas av de intyg som krävs enligt gemenskapslagstiftningen, vid behov kompletterade i enlighet med denna förordning.
(16) Avyttring av vissa animaliska produkter som härrör från nötkreatur i högriskregioner bör förbjudas. Detta förbud bör dock inte gälla vissa animaliska produkter som framställs under kontrollerade förhållanden och som kommer från djur för vilka det kan fastställas att de inte utgör någon hög risk för infektion med TSE.
(17) För att säkerställa att reglerna om förebyggande, kontroll och utrotning av TSE respekteras är det lämpligt att ta prover för laboratorietester på grundval av ett på förhand fastställt protokoll som kan ge en fullständig epidemiologisk bild av läget när det gäller TSE. För att garantera att testförfarandena och testresultaten är enhetliga bör referenslaboratorier inrättas, nationellt och på gemenskapsnivå; därtill måste det införas tillförlitliga vetenskapliga metoder, bland annat specifika snabbtest för TSE. Man bör i möjligaste mån använda snabbtest.
(18) Det är nödvändigt att genomföra gemenskapsinspektioner i medlemsstaterna för att garantera en enhetlig tillämpning av kraven när det gäller förebyggande, kontroll och utrotning av TSE samt även föreskriva tillämpning av kontrollförfaranden. För att säkerställa att de garantier som lämnas av tredje land vid import av levande djur och animaliska produkter till gemenskapen är likvärdiga med dem som är i kraft inom gemenskapen bör gemenskapsinspektioner och -kontroller genomföras på plats för att kontrollera att importvillkoren uppfylls av exporterande tredje land.
(19) Handelsåtgärderna när det gäller TSE bör bygga på internationella standarder, riktlinjer eller rekommendationer, om sådana finns. Åtgärder som är vetenskapligt underbyggda och som säkerställer ett bättre sanitärt skydd får dock vidtas om de åtgärder som är grundade på relevanta internationella standarder, riktlinjer eller rekommendationer inte skulle säkerställa ett lämpligt hälsoskydd.
(20) Det bör föreskrivas att denna förordning skall ses över när nya vetenskapliga uppgifter blir tillgängliga.
(21) De övergångsåtgärder som är nödvändiga för att i synnerhet reglera användningen av de typer av riskmaterial som anges i denna förordning bör fastställas.
(22) De åtgärder som krävs för att genomföra denna förordning bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(4).
(23) I syfte att genomföra denna förordning bör förfaranden fastställas för ett nära och effektivt samarbete mellan kommissionen och medlemsstaterna inom Ständiga veterinärkommittén, Ständiga foderkommittén och Ständiga livsmedelskommittén.
(24) Eftersom tillämpningsföreskrifterna för denna förordning är åtgärder med allmän räckvidd enligt artikel 2 i rådets beslut 1999/468/EG, bör de antas enligt det föreskrivande förfarandet i artikel 5 i det beslutet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
ALLMÄNNA BESTÄMMELSER
Artikel 1
Tillämpningsområde
1. I denna förordning fastställs bestämmelser för förebyggande, kontroll och utrotning av transmissibel spongiform encefalopati (TSE) hos djur. Den skall tillämpas på framställning och avyttring, samt i vissa särskilda fall export, av levande djur och animaliska produkter.
2. Denna förordning skall inte tillämpas på
a) kosmetiska, medicinska eller medicintekniska produkter, eller utgångsmaterial och mellanprodukter till dessa,
b) produkter, eller utgångsmaterial och mellanprodukter till dessa, som inte är avsedda att användas i livsmedel, foder eller gödningsmedel,
c) animaliska produkter som är avsedda för utställning, undervisning, forskning, specialstudier eller analyser, förutsatt att de inte slutligen kan konsumeras eller användas av människor eller andra djur än de som används för de aktuella forskningsprojekten,
d) levande djur som används vid eller är avsedda för forskning.
Artikel 2
Separering av levande djur och animaliska produkter
För att undvika korskontaminering eller substitution av levande djur eller animaliska produkter som avses i artikel 1.1, med de animaliska produkter som avses i artikel 1.2 a-1.2 c eller de levande djur som avses i artikel 1.2 d, skall de hållas permanent åtskilda, såvida inte dessa levande djur eller dessa animaliska produkter har framställts under åtminstone likvärdiga hälsoskyddsvillkor när det gäller TSE.
Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
Artikel 3
Definitioner
1. I denna förordning används följande beteckningar med de betydelser som här anges:
a) TSE: samtliga former av transmissibel spongiform encefalopati utom de som människor kan drabbas av.
b) avyttring: all verksamhet som har till syfte att sälja levande djur eller animaliska produkter som omfattas av denna förordning, till tredje man inom gemenskapen, eller varje annan form av överlåtelse mot eller utan betalning till en sådan tredje man, eller lagring i syfte att senare tillhandahålla en sådan tredje man produkterna.
c) animaliska produkter: alla produkter som härrör från eller innehåller en produkt som härrör från något av de djur som omfattas av bestämmelserna i direktiv 89/662/EEG(5) eller direktiv 90/425/EEG(6).
d) utgångsmaterial: råvaror eller andra animaliska produkter från vilka eller med vars hjälp de produkter som avses i artikel 1.2 a och 1.2 b framställs.
e) behörig myndighet: den centrala myndighet i en medlemsstat som har till uppgift att se till att kraven i denna förordning efterlevs, eller varje annan myndighet till vilken den centrala myndigheten har delegerat nämnda uppgift, särskilt för foderkontroll. Denna definition skall också, i förekommande fall, omfatta motsvarande myndighet i tredje land.
f) kategori: någon av de klassificeringskategorier som avses i kapitel C i bilaga II.
g) specificerat riskmaterial: de vävnader som specificeras i bilaga V. Om inte annat anges, skall produkter som innehåller eller härrör från dessa vävnader inte inbegripas i denna definition.
h) djur som misstänks vara smittade med TSE: levande, slaktade eller döda djur som uppvisar eller har uppvisat neurologiska eller beteendemässiga störningar eller ett gradvis försämrat allmäntillstånd som har samband med en störning i centrala nervsystemet och för vilka ingen alternativ diagnos kan fastställas på grundval av information som inhämtats på grundval av en klinisk undersökning, svar på behandling, obduktion eller laboratorieanalys före eller efter djurets död. Alla nötkreatur som har gett positivt resultat i ett snabbtest för bovin spongiform encefalopati (BSE) skall också misstänkas vara smittade med BSE.
i) anläggning: varje anläggning eller plats där djur som omfattas av denna förordning hålls, föds upp och hanteras eller visas upp för allmänheten.
j) provtagning: provtagning, med statistiskt korrekt underlag, från djur eller deras omgivning eller från animaliska produkter för att ställa en sjukdomsdiagnos eller fastställa släktskap, övervaka hälsan samt kontrollera frånvaron av mikrobiologiska agenser eller vissa material i animaliska produkter.
k) gödningsmedel: varje ämne som innehåller animaliska produkter som används på mark för att främja tillväxten. Det får innehålla rötningsrester från biogasproduktion eller kompostering.
l) snabbtest: de analysmetoder som avses i kapitel C.4 i bilaga X och som ger ett resultat inom 24 timmar.
m) alternativt test: de test som avses i artikel 8.2 och som används i stället för avlägsnande av specificerat riskmaterial.
2. De särskilda definitionerna i bilaga I skall också gälla.
3. Om en term i denna förordning inte har definierats i punkt 1 eller i bilaga I, skall de relevanta definitionerna i förordning (EG) nr 1760/2000(7) och de definitioner som finns i eller som har fastställts med stöd av direktiven 64/432/EEG(8), 89/662/EEG, 90/425/EEG och 91/68/EEG(9) tillämpas i den utsträckning som det hänvisas till dem i denna text.
Artikel 4
Skyddsåtgärder
1. När det gäller genomförandet av skyddsåtgärder skall principerna och bestämmelserna i artikel 9 i direktiv 89/662/EEG, artikel 10 i direktiv 90/425/EEG, artikel 18 i direktiv 91/496/EEG(10) och artikel 22 i direktiv 97/78/EG(11) tillämpas.
2. Skyddsåtgärderna skall antas i enlighet med det förfarande som avses i artikel 24.2 och Europaparlamentet skall samtidigt underrättas om dessa åtgärder och om motiveringen till dem.
KAPITEL II
FASTSTÄLLANDE AV BSE-STATUS
Artikel 5
Klassificering
1. BSE-status för en medlemsstat, ett tredje land eller en region i en medlemsstat eller ett tredje land (nedan kallade länder eller regioner), kan endast fastställas på grundval av kriterierna i kapitel A i bilaga II och resultaten av en riskanalys som identifierar samtliga potentiella faktorer för uppkomsten av BSE, angivna i kapitel B i bilaga II, samt deras utveckling över tiden.
Medlemsstaterna och de tredje länder som vill stå kvar på förteckningarna över tredje länder som är godkända för att till gemenskapen exportera de levande djur eller de produkter som avses i denna förordning, skall till kommissionen lämna en ansökan om fastställande av deras BSE-status, tillsammans med relevanta uppgifter avseende kriterierna i kapitel A i bilaga II och de potentiella riskfaktorerna i kapitel B i bilaga II samt deras utveckling över tiden.
2. Ett beslut om att fatta ett avgörande om varje ansökan för att klassificera den medlemsstat eller det tredje land eller den region i medlemsstaten eller det tredje landet som har lämnat in ansökan såsom hörande till någon av kategorierna i kapitel C i bilaga II, skall fattas med beaktande av de kriterier och potentiella riskfaktorer som anges i punkt 1, i enlighet med det förfarande som avses i artikel 24.2.
Detta beslut skall antas inom sex månader efter det att ansökan samt de relevanta upplysningar som avses i punkt 1, andra stycket, har lämnats in. Om kommissionen finner att underlaget inte innehåller den information som fastställs i kapitlen A och B i bilaga II, skall den begära ytterligare information inom en tidsfrist som skall fastställas. Det slutliga beslutet skall sedan fattas inom sex månader efter det att den fullständiga informationen lämnats.
Efter det att Internationella byrån för epizootiska sjukdomar har fastställt ett förfarande för klassificering av länder i kategorier och om den har placerat det ansökande landet i någon av dessa kategorier, får det beslutas om en förnyad bedömning av den gemenskapskategorisering som genomförts för det berörda landet i enlighet med första stycket i denna punkt, i förekommande fall i enlighet med det förfarande som avses i artikel 24.2.
3. Om kommissionen finner att den information som en medlemsstat eller ett tredje land har lämnat i enlighet med kapitlen A och B i bilaga II är otillräcklig eller oklar, kan den i enlighet med det förfarande som avses i artikel 24.2 fastställa BSE-status för den berörda medlemsstaten eller det berörda tredje landet på grundval av en fullständig riskanalys.
Denna analys skall innehålla en avgörande statistisk undersökning av den epidemiologiska situationen avseende TSE i den ansökande medlemsstaten eller det ansökande tredje landet, vilken skall genomföras med snabbtest med hjälp av ett screeningförfarande. Kommissionen skall beakta de klassificeringskriterier som Internationella byrån för epizootiska sjukdomar har fastställt.
Snabbtest skall godkännas för detta ändamål enligt det förfarande som avses i artikel 24.2 och införas i en förteckning i kapitel C.4 i bilaga X.
Detta screeningförfarande kan även utnyttjas av de medlemsstater eller tredje länder som vill att kommissionen - enligt det förfarande som avses i artikel 24.2 - skall godkänna den klassificering som de gjort på denna grund.
Den berörda medlemsstaten eller det berörda tredje landet skall stå för kostnaderna för detta förfarande.
4. De medlemsstater eller tredje länder som inte lämnat in någon ansökan enligt punkt 1 inom sex månader från och med den 1 juli 2001 skall, när det gäller export från deras territorier av levande djur eller animaliska produkter, betraktas som länder i kategori 5 enligt kapitel C i bilaga II så länge de inte har lämnat in någon ansökan.
5. Medlemsstaterna skall utan dröjsmål till kommissionen anmäla alla epidemiologiska bevis eller annan information som skulle kunna leda till förändringar i deras BSE-status, särskilt resultaten av de övervakningsprogram som föreskrivs i artikel 6.
6. Bibehållandet av ett tredje land i någon av förteckningarna enligt gemenskapens bestämmelser om tillstånd att till Europeiska gemenskapen exportera levande djur och animaliska produkter, för vilka det finns särskilda bestämmelser i denna förordning, beslutas enligt det förfarande som anges i artikel 24.2 och under förutsättning att, med hänsyn till tillgänglig information eller om TSE förmodas förekomma - den information som föreskrivs i punkt 1 lämnas. Om sådan information inte lämnas inom tre månader från det att kommissionen begärt den, skall bestämmelserna i punkt 4 i denna artikel tillämpas så länge informationen inte har lämnats och inte har kunnat utvärderas i enlighet med punkt 2 eller punkt 3.
För att tredje land skall få exportera levande djur eller animaliska produkter för vilka det finns särskilda bestämmelser i denna förordning till gemenskapen enligt de villkor som grundar sig på den kategori som kommissionen fastställt, skall de förbinda sig att utan dröjsmål till kommissionen skriftligen anmäla alla epidemiologiska eller andra bevis som skulle kunna leda till ändringar i deras BSE-status.
7. Ett beslut får antas i enlighet med det förfarande som avses i artikel 24.2 om att ändra BSE(klassificeringen för en medlemsstat eller ett tredje land eller någon av deras regioner i enlighet med resultaten av de kontroller som föreskrivs i artikel 21.
8. De beslut som avses i punkterna 2, 3, 4, 6 och 7 skall grundas på en riskbedömning med hänsyn till de rekommenderade kriterier som fastställs i kapitlen A och B i bilaga II.
KAPITEL III
FÖREBYGGANDE AV TSE
Artikel 6
Övervakningssystem
1. Varje medlemsstat skall genomföra ett årligt övervakningsprogram för BSE och scrapie i enlighet med kapitel A i bilaga III. Ett screeningförfarande med hjälp av snabbtest skall ingå i detta program.
Snabbtest skall godkännas för detta ändamål enligt det förfarande som avses i artikel 24.2 och införas i en förteckning i kapitel C.4 i bilaga X.
2. Medlemsstaterna skall underrätta kommissionen och de övriga medlemsstaterna i Ständiga veterinärkommittén om uppkomst av annan TSE än BSE.
3. Alla officiella undersökningar och laboratorieprov skall registreras enligt kapitel B.1 bilaga III.
4. Medlemsstaterna skall förelägga kommissionen en årlig rapport som skall innehålla åtminstone den information som avses i kapitel B.I i bilaga III. Rapporten för varje kalenderår skall överlämnas senast den 31 mars nästkommande år. Inom tre månader efter det att de nationella rapporterna har mottagits, skall kommissionen för Ständiga veterinärkommittén lägga fram en sammanfattning av dessa rapporter, som skall innehålla åtminstone den information som avses i kapitel B.II i bilaga III.
Artikel 7
Förbud avseende foder
1. Det är förbjudet att utfodra idisslare med protein som härrör från däggdjur.
2. Dessutom skall det förbud som avses i punkt 1 även gälla djur och animaliska produkter i enlighet med punkt 1 i bilaga IV.
3. Punkterna 1 och 2 skall tillämpas utan att det påverkar tillämpningen av punkt 2 i bilaga IV.
4. De medlemsstater eller regioner i medlemsstaterna som har placerats i kategori 5 skall inte tillåtas att exportera eller lagra sådant foder för livsmedelsproducerande djur som innehåller protein som härrör från däggdjur, eller foder som är avsett för däggdjur, med undantag av hundar och katter, och som innehåller bearbetat protein som härrör från däggdjur.
Tredje land eller regioner i tredje land som har placerats i kategori 5 skall inte tillåtas att till gemenskapen exportera sådant foder för livsmedelsproducerande djur som innehåller protein som härrör från däggdjur eller foder som är avsett för däggdjur, med undantag av hundar och katter, och som innehåller bearbetat protein som härrör från däggdjur.
5. Tillämpningsföreskrifterna för denna artikel, inbegripet reglerna om förebyggande av korskontaminering och om de metoder för provtagning och provanalys som krävs för att kontrollera att denna artikel efterlevs, skall antas enligt det förfarande som avses i artikel 24.2.
Artikel 8
Specificerat riskmaterial
1. Det specificerade riskmaterialet skall avlägsnas och destrueras i enlighet med punkterna 2, 3, 4 och 8 i bilaga V.
Dessa specificerade riskmaterial eller bearbetade material av dessa får endast avyttras eller, i förekommande fall, exporteras för slutlig destruktion i enlighet med punkterna 3 och 4 eller i förekommande fall punkt 7 c eller punkt 8 i bilaga V. De får inte importeras till gemenskapen. Transitering genom gemenskapens territorium skall ske i överensstämmelse med kraven i artikel 3 i direktiv 91/496/EEG.
2. Punkt 1 skall inte tillämpas på vävnader från djur som har genomgått ett alternativt test som godkänts för detta särskilda syfte i enlighet med det förfarande som avses i artikel 24.2 och som införts i förteckningen i kapitel C.5 i bilaga X och tillämpas enligt de villkor som anges i punkt 5 i bilaga V, och där testresultaten är negativa.
De medlemsstater som godkänner detta alternativa test skall underrätta de övriga medlemsstaterna och kommissionen om detta.
3. I de medlemsstater eller regioner inom dessa som har placerats i kategorierna 2, 3, 4 och 5 enligt kapitel C i bilaga II får laceration, efter bedövning, av vävnad från centrala nervsystemet med ett avlångt, stavformigt instrument som förs in i hjärnskålen inte användas för nötkreatur, får eller getter vars kött är avsett som livsmedel eller foder.
4. De uppgifter om ålder som anges i bilaga V skall anpassas regelbundet. Denna anpassning skall genomföras på grundval av de senaste säkra vetenskapliga rönen om den statistiska sannolikheten för att TSE förekommer inom de berörda åldersgrupperna av gemenskapens bestånd av nötkreatur, får och getter.
5. Trots vad som sägs i punkterna 1-4 kan ett beslut antas i enlighet med det förfarande som avses i artikel 24.2 om den dag då bestämmelserna i artikel 7.1 skall börja gälla eller i förekommande fall i tredje land om den dag förbudet skall träda i kraft mot användning av proteiner som härrör från däggdjur i foder för idisslare i samtliga länder eller regioner som placerats i kategori 3 eller 4, i syfte att begränsa tillämpningen av denna artikel till djur som har fötts före denna dag i dessa länder eller regioner.
Trots vad som sägs i artiklarna 1-4, kan efter samråd med den behöriga vetenskapliga kommittén och på grundval av en bedömning av risken för förekomst eller spridning av sjukdomen eller för att människor utsätts för smitta, ett beslut likaså fattas i enlighet med det förfarande som avses i artikel 24.2 om att tillåta att kotpelare och dorsala rotganglier från nötkreatur i eller från de länder eller regioner som placerats i kategori 5, används i livsmedel, foder och gödningsämnen.
6. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
Artikel 9
Animaliska produkter som härrör från eller innehåller material från idisslare
1. De animaliska produkter som räknas upp i bilaga VI får inte framställas av material som härrör från idisslare från länder eller regioner som är placerade i kategori 5, såvida de inte framställs i enlighet med de produktionsprocesser som har godkänts i enlighet med det förfarande som avses i artikel 24.2.
2. Skallben och kotpelare från nötkreatur, får och getter från länder eller regioner som är placerade i kategori 2, 3, 4 eller 5 får inte användas för framställning av mekaniskt urbenat kött.
3. Bestämmelserna i punkterna 1 och 2 skall, när det gäller kriterierna i punkt 5 i bilaga V, inte tillämpas på idisslare som har genomgått ett alternativt test som godkänts enligt det förfarande som avses i artikel 24.2 och där testresultaten är negativa.
4. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
Artikel 10
Utbildningsprogram
1. Medlemsstaterna skall se till att personalen vid den behöriga myndigheten, diagnostiska laboratorier samt utbildningsanstalter för lantbruk och veterinärmedicin, officiella veterinärer, praktiserande veterinärer, slakteripersonal samt personer som föder upp, håller och hanterar djur får utbildning när det gäller kliniska tecken, epidemiologi samt, när det gäller personal som har ansvar för inspektionerna, utbildning i att tolka laboratorieresultat som rör TSE.
2. För att de utbildningsprogram som avses i punkt 1 skall kunna genomföras effektivt får gemenskapen bevilja ekonomiskt stöd. Beloppet för ett sådant stöd skall bestämmas enligt det förfarande som avses i artikel 24.2.
KAPITEL IV
KONTROLL OCH UTROTNING AV TSE
Artikel 11
Anmälan
Utan att det påverkar tillämpningen av direktiv 82/894/EEG(12) skall medlemsstaterna se till att alla djur som misstänks vara smittade med TSE omedelbart anmälas till de behöriga myndigheterna.
Medlemsstaterna skall regelbundet underrätta övriga medlemsstater och kommissionen om anmälda fall av TSE.
Den behöriga myndigheten skall utan dröjsmål vidta de åtgärder som fastställs i artikel 12 i denna förordning, liksom alla andra nödvändiga åtgärder.
Artikel 12
Åtgärder vid misstänkta fall
1. Alla djur som misstänks vara smittade med TSE skall vara föremål för officiella restriktioner vad avser förflyttning i avvaktan på att resultaten av den behöriga myndighetens kliniska och epidemiologiska undersökning blir tillgängliga, eller avlivas för laboratorieundersökning under officiell kontroll.
Om man misstänker BSE hos ett nötkreatur på en anläggning i en medlemsstat, skall alla övriga nötkreatur på denna anläggning vara föremål för officiella restriktioner vad avser förflyttning i avvaktan på att resultaten av undersökningen blir tillgängliga.
Om man misstänker BSE hos ett får eller en get på en anläggning i en medlemsstat på grundval av objektiva faktorer såsom resultaten av ett test som på ett praktiskt sätt kan göra åtskillnad mellan olika typer av TSE, skall alla övriga får och getter på anläggningen vara föremål för officiella restriktioner vad avser förflyttning i avvaktan på att resultaten av undersökningen blir tillgängliga.
Om det kan styrkas att den anläggning där djuret befann sig när man misstänkte BSE förmodligen inte är den anläggning där djuret kan ha exponerats för BSE, får den behöriga myndigheten besluta att bara det djur som misstänks vara smittat skall vara föremål för en officiell restriktion vad avser förflyttning. Om den behöriga myndigheten anser det nödvändigt, får den också besluta att övriga anläggningar eller endast den anläggning där exponeringen förekom skall ställas under officiell övervakning, beroende på den tillgängliga epidemiologiska informationen.
En medlemsstat får, enligt det förfarande som avses i artikel 24.2 och med avvikelse från kraven i andra, tredje och fjärde styckena i denna punkt, undantas från tillämpning av officiella restriktioner vad avser förflyttning av djur, om medlemsstaten tillämpar åtgärder som erbjuder likvärdiga garantier.
2. Om den behöriga myndigheten beslutar att det inte kan uteslutas att ett djur har smittats av TSE, skall djuret - om det fortfarande är vid liv - avlivas; dess hjärna, liksom alla övriga vävnader som den behöriga myndigheten bestämmer, skall avlägsnas och skickas till ett officiellt godkänt laboratorium, det nationella referenslaboratoriet enligt artikel 19.1 eller gemenskapens referenslaboratorium enligt artikel 19.2, för att undersökas där enligt de testmetoder som anges i artikel 20.
3. Alla delar av det misstänkta djurets kropp, inklusive huden, skall hållas under officiell övervakning till dess en negativ diagnos har ställts, eller destrueras i enlighet med punkt 3 eller 4 i bilaga V.
4. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
Artikel 13
Åtgärder vid bekräftad förekomst av TSE
1. Om förekomst av TSE har bekräftats officiellt, skall följande åtgärder vidtas utan dröjsmål:
a) Samtliga delar av det smittade djurets kropp skall destrueras fullständigt i enlighet med bilaga V, med undantag för det material som skall bevaras för registren i enlighet med kapitel B.III.2 i bilaga III.
b) En undersökning skall genomföras för att identifiera alla riskdjur i enlighet med punkt 1 i bilaga VII.
c) Alla djur och animaliska produkter som avses i punkt 2 i bilaga VII och som vid den undersökning som avses i punkt b har konstaterats vara riskdjur, skall avlivas och destrueras fullständigt i enlighet med punkterna 3 och 4 i bilaga V.
En medlemsstat får, trots bestämmelserna i detta stycke, tillämpa andra åtgärder som erbjuder motsvarande skyddsnivå, om dessa åtgärder har godkänts enligt det förfarande som avses i artikel 24.2.
2. I avvaktan på att de åtgärder som avses i punkterna 1 b och 1 c genomförs, skall den anläggning där djuret befann sig när förekomsten av TSE bekräftades ställas under officiell övervakning och all förflyttning från eller till anläggningen av djur som riskerar att ha smittats med TSE samt av animaliska produkter från dessa djur godkännas av den behöriga myndigheten, så att djuren och de berörda animaliska produkterna omedelbart skall kunna spåras och identifieras.
Om det kan styrkas att anläggningen där det smittade djuret befann sig när TSE bekräftades förmodligen inte är den anläggning där djuret exponerats för TSE, får den behöriga myndigheten besluta att båda anläggningarna eller bara den anläggning där djuret exponerats skall placeras under officiell övervakning.
3. De medlemsstater som har genomfört ett alternativt system som erbjuder likvärdiga garantier enligt artikel 12.1 femte stycket får, enligt det förfarande som avses i artikel 24.2 och med avvikelse från kraven i punkterna 1 b och 1 c, undantas från skyldigheten att tillämpa det officiella förbudet mot förflyttning av djuren och från kravet på att avliva och destruera djuren.
4. Ägarna skall utan dröjsmål ersättas för förlusten av de djur som har avlivats och de animaliska produkter som har destruerats i enlighet med artikel 12.2 och punkterna 1 a och 1 c i denna artikel.
5. Utan att det påverkar tillämpningen av direktiv 82/894/EEG skall varje bekräftat fall av en annan typ av TSE än BSE anmälas till kommissionen på årlig basis.
6. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
Artikel 14
Beredskapsplan
1. Medlemsstaterna skall - i enlighet med de allmänna kriterierna i gemenskapens bestämmelser för kontroll av djursjukdomar - utarbeta riktlinjer som specificerar vilka nationella åtgärder som skall genomföras och ange behörighet och ansvar om TSE-fall bekräftas.
2. Om det är nödvändigt för att möjliggöra en enhetlig tillämpning av gemenskapslagstiftningen får riktlinjerna harmoniseras enligt det förfarande som avses i artikel 24.2.
KAPITEL V
AVYTTRING OCH EXPORT
Artikel 15
Levande djur, deras sperma, embryon och ägg
1. Avyttring eller i förekommande fall export av nötkreatur, får eller getter och deras sperma, embryon och ägg skall omfattas av de villkor som anges i bilaga VIII eller, vid import, de villkor som anges i bilaga IX. De levande djuren och deras embryon och ägg skall åtföljas av de relevanta hälsointyg som föreskrivs i gemenskapslagstiftningen i enlighet med artikel 17 eller, vid import, i enlighet med artikel 18.
2. Avyttring av den första generationen avkomma, sperma, embryon och ägg från djur som misstänks eller bekräftats vara smittade med TSE skall omfattas av de villkor som anges i kapitel B i bilaga VIII.
3. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
Artikel 16
Avyttring av animaliska produkter
1. Följande animaliska produkter från friska idisslare skall inte vara föremål för restriktioner när de avyttras eller i förekommande fall exporteras enligt denna artikel och enligt bestämmelserna i kapitlen C och D i bilaga VIII och i kapitlen A, C, F och G i bilaga IX:
a) Animaliska produkter som omfattas av bestämmelserna i artikel 15, särskilt sperma, embryon och ägg.
b) i) Rå mjölk enligt definitionen i direktiv 92/46/EEG(13).
ii) Mjölk avsedd för framställning av mjölkbaserade produkter enligt definitionen i direktiv 92/46/EEG.
iii) Värmebehandlad konsumtionsmjölk enligt definitionen i direktiv 92/46/EEG.
iv) Dikalciumfosfat (utan spår av protein eller fett).
v) Hudar och skinn i den mening som avses i direktiv 92/118/EEG(14).
vi) Gelatin i den mening som avses i direktiv 92/118/EEG som härrör från hudar och skinn enligt punkt v.
vii) Kollagen som härrör från hudar och skinn enligt punkt v.
2. Animaliska produkter från tredje land som har placerats i kategorierna 2, 3, 4 och 5 skall härröra från nötkreatur, får och getter som inte har utsatts för sådan laceration av vävnad från centrala nervsystemet som anges i artikel 8.3, eller avlivats med gas som har injicerats i hjärnskålen.
3. Animaliska produkter som innehåller material från nötkreatur med ursprung i en medlemsstat, en region i en medlemsstat eller ett tredje land som placerats i kategori 5 får inte avyttras utom i de fall då de härrör från
a) djur som är födda efter den dag då förbudet mot utfodring av idisslare med bearbetat protein som härrör från däggdjur började gälla,
b) djur som är födda, har fötts upp och hållits i besättningar som bevisligen varit BSE-fria sedan minst 7 år tillbaka i tiden.
Animaliska produkter får inte skickas från en medlemsstat eller en region i en medlemsstat som placerats i kategori 5, från en annan medlemsstat eller importeras från ett tredje land som placerats i kategori 5. Detta förbud gäller inte sådana animaliska produkter som avses i kapitel C i bilaga VIII och som uppfyller kraven i kapitel C i bilaga VIII. De skall åtföljas av ett hälsointyg som utfärdats av en officiell veterinär som intygar att de framställts i enlighet med denna förordning.
4. Om ett djur förflyttas från ett land eller en region till ett annat land eller en annan region placerade i en annan kategori, skall det klassificeras i den högsta kategorin för de länder eller regioner där det har vistats mer än ett dygn, såvida inte tillräckliga garantier om att djuret inte har utfodrats med foder från detta land eller denna region som klassificerats i den högsta kategorin kan lämnas.
5. De animaliska produkter för vilka det anges särskilda regler i denna artikel skall åtföljas av sådana lämpliga hälsointyg eller handelsdokument som föreskrivs i gemenskapslagstiftningen i enlighet med artiklarna 17 och 18 eller, om det inte finns något sådant krav i gemenskapslagstiftningen, av ett hälsointyg eller ett handelsdokument, för vilka modeller skall fastställas i enlighet med det förfarande som avses i artikel 24.2.
6. För import till gemenskapen skall animaliska produkter uppfylla kraven i kapitlen A, C, F och G i bilaga IX.
7. Enligt det förfarande som avses i artikel 24.2 får bestämmelserna i punkterna 1-6 utvidgas till att omfatta andra animaliska produkter. Tillämpningsföreskrifter för denna artikel skall fastställas enligt samma förfarande.
Artikel 17
Enligt det förfarande som avses i artikel 24.2 skall de hälsointyg som avses i bilaga F till direktiv 64/432/EEG och i modellerna II och III i bilaga E till rådets direktiv 91/68/EEG, samt de lämpliga hälsointyg som föreskrivs i gemenskapslagstiftningen om handel med sperma, ägg och embryon från nötkreatur, får eller getter vid behov kompletteras med en uppgift om kategori med angivande av den klassificering av medlemsstaten eller ursprungsregionen som gjorts enligt artikel 5.
Lämpliga handelsdokument för handel med animaliska produkter skall i förekommande fall kompletteras med en uppgift om den kategori som kommissionen i enlighet med artikel 5 placerat medlemsstaten eller ursprungsregionen i.
Artikel 18
Lämpliga hälsointyg för import som föreskrivs i gemenskapslagstiftningen skall, enligt det förfarande som avses i artikel 24.2, kompletteras med de särskilda kraven i bilaga IX när det gäller tredje länder som klassificerats i en kategori i enlighet med artikel 5, så snart detta beslut om klassificering har antagits.
KAPITEL VI
REFERENSLABORATORIER, PROVTAGNING, UNDERSÖKNINGAR OCH KONTROLLER
Artikel 19
Referenslaboratorier
1. De nationella referenslaboratorierna i varje medlemsstat samt deras behörighet och uppgifter fastställs i kapitel A i bilaga X.
2. Gemenskapens referenslaboratorium, dess behörighet och uppgifter fastställs i kapitel B i bilaga X.
Artikel 20
Provtagning och metoder för laboratorieanalyser
1. Provtagning och laboratorieundersökningar för att fastställa förekomst av TSE skall genomföras enligt de metoder och protokoll som anges i kapitel C i bilaga X.
2. När så krävs för att möjliggöra en enhetlig tillämpning av denna artikel, skall tillämpningsföreskrifter - inbegripet metoden för att bekräfta förekomst av BSE hos får och getter - fastställas enligt det förfarande som avses i artikel 24.2.
Artikel 21
Gemenskapskontroller
1. Experter från kommissionen får, när så krävs för en enhetlig tillämpning av denna förordning, i samarbete med de behöriga myndigheterna i medlemsstaterna genomföra kontroller på plats. Den medlemsstat på vars territorium en kontroll utförs skall ge all nödvändig hjälp till experterna så att de kan fullgöra sina uppgifter. Kommissionen skall underrätta den behöriga myndigheten om resultaten av de utförda kontrollerna.
Tillämpningsföreskrifter för denna artikel, särskilt sådana som syftar till att reglera formerna för samarbete med de nationella myndigheterna, skall fastställas enligt det förfarande som avses i artikel 24.2.
2. Gemenskapskontrollerna vad avser tredje land skall ske i enlighet med artiklarna 20 och 21 i direktiv 97/78/EG.
KAPITEL VII
ÖVERGÅNGSBESTÄMMELSER OCH SLUTBESTÄMMELSER
Artikel 22
Övergångsbestämmelser för specificerat riskmaterial
1. Bestämmelserna i del A i bilaga XI skall tillämpas under en period på minst sex månader räknat från den 1 juli 2001; denna period upphör samma dag som ett beslut har antagits i enlighet med bestämmelserna i artikel 5.2 eller 5.4; från och med den dagen skall artikel 8 tillämpas.
2. Resultaten av en avgörande statistisk undersökning, som under övergångsperioden utförs i enlighet med bestämmelserna i artikel 5.3, skall utnyttjas för att bekräfta eller vederlägga slutsatserna från den riskanalys som avses i artikel 5.1, varvid de klassificeringskriterier som fastställts av Internationella byrån för epizootiska sjukdomar skall beaktas.
3. Detaljerade bestämmelser om denna statistiska undersökning skall, efter samråd med den relevanta vetenskapliga kommittén, antas enligt det förfarande som avses i artikel 24.2.
4. De minimikriterier som denna statistiska undersökning skall uppfylla fastställs i del B i bilaga XI.
Artikel 23
Ändring av bilagorna och övergångsbestämmelser
Efter samråd med den relevanta vetenskapliga kommittén om sådana frågor som kan ha konsekvenser för folkhälsan skall bilagorna ändras eller kompletteras och lämpliga övergångsbestämmelser antas, i enlighet med det förfarande som avses i artikel 24.2.
Enligt det förfarandet skall övergångsbestämmelser antas för en period på högst två år för att möjliggöra en övergång från nuvarande ordning till den ordning som fastställs i denna förordning.
Artikel 24
Kommittéer
1. Kommissionen skall biträdas av Ständiga veterinärkommittén. I frågor som uteslutande rör foder skall kommissionen dock biträdas av Ständiga foderkommittén, och i frågor som uteslutande rör livsmedel skall kommissionen biträdas av Ständiga livsmedelskommittén.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader, och när det gäller skyddsåtgärder enligt artikel 4.2 i denna förordning skall tiden vara 15 dagar.
3. Varje kommitté skall själva anta sin arbetsordning.
Artikel 25
Samråd med vetenskapliga kommittéer
De relevanta vetenskapliga kommittéerna skall höras i alla frågor som omfattas av tillämpningsområdet för denna förordning och som kan ha konsekvenser för folkhälsan.
Artikel 26
Ikraftträdande
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1282/2001
av den 28 juni 2001
om tillämpningsföreskrifter för rådets förordning (EG) nr 1493/1999 om framtagning av uppgifter för produktinformation och marknadsuppföljning inom vinsektorn och om ändring av förordning (EG) nr 1623/2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1493/1999 av 17 maj 1999 om den gemensamma organisationen av marknaden för vin(1), senast ändrad genom förordning (EG) nr 2826/2000(2), särskilt artiklarna 23, 33 och 73 i denna, och
av följande skäl:
(1) I artikel 18 i förordning (EG) nr 1493/1999 föreskrivs att producenter av druvor avsedda för vinframställning och producenter av druvmust och vin varje år skall deklarera vilka mängder som producerats av den senaste skörden, samt att både producenter av druvmust och vin och andra näringsidkare än detaljhandlare varje år skall deklarera sina lager av druvmust och vin.
(2) I samma artikel föreskrivs att medlemsstaterna även får kräva att försäljare av druvor varje år skall deklarera vilka mängder som saluförts från den senaste skörden.
(3) För att underlätta förvaltningen av marknaden för vin måste ett datum anges då deklarationerna skall göras. Eftersom skörden äger rum vid olika tidpunkter i de olika medlemsstaterna bör tidsfristerna för inlämning av producenternas deklarationer spridas över en lämplig period. Även de aktörer som levererar vinprodukter före de angivna deklarationsdatumen bör åläggas att lämna deklarationer.
(4) Det är inte nödvändigt att kräva två deklarationer från producenter som kan lämna alla nödvändiga uppgifter i produktionsdeklarationen. Småproducenter kan undantas från deklarationsskyldighet eftersom deras sammanlagda produktion utgör en relativt blygsam andel av produktionen inom gemenskapen.
(5) Medlemsstaterna får själva närmare besluta om på vilket sätt företagen skall lämna de uppgifter som skall ingå i deklarationen, men för att underlätta tillämpningen av denna förordning bör det föreskrivas att uppgifterna skall lämnas i tabellform. Det är också nödvändigt att fastställa tidsfrister inom vilka medlemsstaterna skall sammanställa och överlämna de insamlade uppgifterna till kommissionen, samt att ange på vilket sätt de skall överlämnas.
(6) Kategorin "annat vin" bör definieras i förhållande till den klassificering av druvsorter som får odlas inom gemenskapen som fastställs i artikel 19 i förordning (EG) nr 1493/1999.
(7) Uppgifterna om vinarealerna kan vara oriktiga på grund av att deklaranten inte har haft de kontrollmöjligheter som krävs. I sådana fall bör påföljden stå i proportion till hur grava felen är i den inlämnade deklarationen.
(8) Påföljdssystemet bör tillåta en tillräcklig grad av proportionalitet för de av vinproducenternas deklarationer som vid kontroll har visats vara ofullständiga eller oriktiga. Påföljden bör anpassas efter de rättelser som görs i en deklaration.
(9) Tillräcklig information om produktion och lager inom vinsektorn återfinns för närvarande bara i de skörde- och lagerdeklarationer som lämnas av de berörda parterna. Lämpliga åtgärder bör därför vidtas för att säkerställa att dessa deklarationer lämnas av vederbörande och att de är fullständiga och korrekta. Det bör ges möjlighet till påföljder för den händelse att deklarationer inte lämnas eller är felaktiga eller ofullständiga. För att förenkla behandlingen av deklarationsuppgifterna bör varje deklaration som lämnas in i den behöriga administrativa enheten anses vara oberoende av andra deklarationer som samma producent kan ha lämnat in till andra av medlemsstatens administrativa enheter.
(10) Enligt rådets förordning (EEG) nr 2392/86(3), senast ändrad genom förordning (EG) nr 1631/98(4), skall ett gemenskapsregister över vinodlingar upprättas. De medlemsstater som förfogar över ett fullständigt register bör tillåtas att använda vissa uppgifter ur registret om de inte finns i deklarationen.
(11) Vissa uppgifter om vinmarknaden är nödvändiga för marknadsuppföljningen. Utöver uppgifter från sammanställningar av de olika deklarationerna måste även tillgängliga mängden, deras användning samt vinpriser uppges. Därför bör det föreskrivas att medlemsstaterna skall samla in uppgifterna och överlämna dem till kommissionen senast vissa angivna datum.
(12) I detta sammanhang är det lämpligt att erinra om att det är nödvändigt att respektera de tidsfrister som fastställs för överföring av uppgifterna för att säkerställa marknadsuppföljningen och se till att effektiva åtgärder inom ramen för budgeten kan vidtas i rätt tid.
(13) För att uppnå nödvändig överensstämmelse mellan de påföljder som föreskrivs i denna förordning och påföljderna enligt kommissionens förordning (EG) nr 1623/2000(5), senast ändrad genom förordning (EG) nr 545/2001(6), är det lämpligt att ändra sistnämnda förordning och införa en lämplig formulering om påföljderna.
(14) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för vin.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Denna förordning gäller tillämpningsföreskrifter för förordning (EG) nr 1493/1999, främst när det gäller framtagning av uppgifter som ökar produktkunskapen och som kan användas för marknadsuppföljning inom vinsektorn.
Artikel 2
1. Fysiska eller juridiska personer eller sammanslutningar av sådana personer som odlar druvor, nedan kallade skördare, skall varje år till de behöriga myndigheter som har utsetts av medlemsstaterna överlämna en skördedeklaration till den administrativa enhet som fastställs. Skördedeklarationen skall minst innehålla de uppgifter som framgår av tabell A och, i förekommande fall, tabell B i bilagan.
I förekommande fall får medlemsstaterna tillåta att en deklaration lämnas per jordbruksföretag.
2. Följande personer behöver emellertid inte lämna in någon skördedeklaration:
a) Skördare vars hela produktion av druvor är avsedd för konsumtion i färskt tillstånd, för torkning eller för omedelbar bearbetning till druvsaft.
b) Skördare vars jordbruksföretag omfattar mindre än 10 ar vinodlingsareal och som varken har sålt eller kommer att sälja någon del av sin produktion i någon form.
c) Skördare vars jordbruksföretag omfattar mindre än 10 ar vinodlingsareal och som levererar hela skörden till ett vinkooperativ eller en sammanslutning som de tillhör eller är associerade med. I sådana fall skall skördarna till jordbrukskooperativen eller sammanslutningarna lämna deklarationer med uppgift om
i) vinodlarens förnamn, efternamn och adress,
ii) den mängd druvor som levereras,
iii) den berörda vinodlingens areal och läge.
I det sista fallet skall vinkooperativet eller sammanslutningen kontrollera att uppgifterna i deklarationen stämmer med de uppgifter som kooperativet har.
3. Med undantag från punkt 1 första stycket, och utan att detta påverkar de skyldigheter som följer av artikel 4, får medlemsstaterna undanta följande personer från skyldigheten att lämna skördedeklarationer:
a) Skördare som själva bearbetar hela sin druvskörd till vin eller som låter bearbeta den för egen räkning.
b) Skördare som är anslutna till eller tillhör ett vinkooperativ eller en sammanslutning och som levererar hela sin skörd, i form av vin eller druvmust, till detta vinkooperativ eller denna sammanslutning, inklusive sådana skördare som avses i artikel 4.4.
Artikel 3
Artikel 4
1. Fysiska eller juridiska personer eller sammanslutningar av sådana personer, inbegripet vinkooperativ, som av innevarande vinårs skörd har framställt vin och/eller vid de tidpunkter som anges i artikel 11.1 innehar andra produkter än vin, skall varje år till de behöriga myndigheter som har utsetts av medlemsstaterna överlämna en produktionsdeklaration som innehåller minst de uppgifter som skall anges enligt tabell C i bilagan.
2. Medlemsstaterna får föreskriva att fysiska eller juridiska personer eller sammanslutningar av sådana personer, inbegripet vinkooperativ, som före de tidpunkter som anges i artikel 11.1 har behandlat eller salufört produkter i tidigare produktionsled än vin under innevarande vinår, till de behöriga myndigheterna skall lämna in behandlings- eller saluföringsdeklarationer som minst skall innehålla uppgifterna enligt tabell C.
3. De skördare som avses i artikel 2.2 samt de producenter som i egna anläggningar av inköpta produkter framställer mindre än tio hektoliter vin, som varken har saluförts eller kommer att saluföras i någon form, är inte skyldiga att lämna någon produktions-, eller i förekommande fall behandlings- eller saluföringsdeklaration.
4. Undantagna från skyldigheten att lämna produktionsdeklaration är även skördare som tillhör ett vinkooperativ som skall lämna produktionsdeklaration och som levererar hela sin druvskörd till kooperativet, men som förbehåller sig rätten att för sin familjs bruk framställa mindre än 10 hektoliter vin.
5. Beträffande fysiska eller juridiska personer eller sammanslutningar av sådana personer, som överlåter vinprodukter i produktionsleden före vin, skall medlemsstaterna vidta nödvändiga åtgärder för att se till att producenter som skall lämna deklarationer har tillgång till de uppgifter som skall ingå.
Artikel 5
Oaktat bestämmelserna i artikel 4 får medlemsstater, som i enlighet med förordning (EEG) nr 2392/86 har upprättat ett fullständigt register över vinodlingar som uppdateras varje år eller ett annat liknande administrativt kontrollinstrument, undanta de fysiska eller juridiska personer, sammanslutningar av sådana personer eller skördare som avses i denna artikel från skyldigheten att deklarera areal.
I dessa fall skall de behöriga myndigheter som har utsetts av medlemsstaten själva fylla i de deklarationer som avses i denna artikel med uppgifter om arealen som bygger på uppgifterna i vinodlingsregistret.
Artikel 6
1. Fysiska eller juridiska personer eller sammanslutningar av sådana personer, med undantag av privata konsumenter och detaljister, skall varje år till de behöriga myndigheter som har utsetts av medlemsstaterna deklarera de lager av druvmust, koncentrerad druvmust, rektifierad koncentrerad druvmust och vin som de innehar den 31 juli. Vinprodukter från gemenskapen skall inte tas med i denna deklaration om de framställts av druvor som skördats under innevarande kalenderår.
Medlemsstater med en årlig vinproduktion av högst 25000 hektoliter får emellertid utöver detaljister undanta även andra handelsidkare som innehar små lager från skyldigheten att lämna de deklarationer som avses i första stycket, förutsatt att de behöriga myndigheterna kan ge kommissionen en statistisk uppskattning av dessa lagers storlek i medlemsstaten.
2. I punkt 1 avses med detaljister fysiska eller juridiska personer eller sammanslutningar av sådana personer vars affärsverksamhet omfattar försäljning av vin i små mängder direkt till konsumenten, med undantag för de detaljister som har vinkällare avsedda för lagring och tappning av stora mängder vin.
De mängder som avses i första stycket skall fastställas enskilt av varje medlemsstat med hänsyn till handelns och distributionens särskilda egenskaper.
3. Den deklaration som avses i punkt 1 skall innehålla minst de uppgifter som framgår av tabell D i bilagan.
Artikel 7
1. Medlemsstaterna skall utarbeta formulär för de olika deklarationerna och säkerställa att dessa innehåller minst de uppgifter som anges i tabellerna A, B, C och D i bilagan.
Formulären behöver inte innehålla någon uttrycklig hänvisning till areal om medlemsstaten med säkerhet kan bestämma denna med hjälp av andra uppgifter som lämnas i deklarationen eller i vinodlingsregistret, särskilt produktionsarealen och jordbruksföretagets totala skörd.
Den information som innefattas i de deklarationer som avses i första stycket skall behandlas centralt på nationell nivå.
Medlemsstaterna skall besluta om nödvändiga kontrollåtgärder för att säkerställa att deklarationerna överensstämmer med verkligheten.
De skall underrätta kommissionen om dessa åtgärder och översända de formulär som utarbetas enligt första stycket.
2. Medlemsstater vars vinodlingsareal inte överstiger 100 ha och som har
- fått vissa av de uppgifter som skall anges i deklarationerna enligt kapitlen I och II från andra administrativa handlingar behöver inte kräva att dessa uppgifter skall finnas med i deklarationerna,
- fått alla de uppgifter som skall anges i deklarationerna enligt kapitlen I och II från andra administrativa handlingar får undanta aktörerna i fråga från skyldigheten att lämna in en eller flera av deklarationerna.
De medlemsstater i vilka kapitlen I och II i avdelning II i förordning (EG) nr 1493/1999 inte tillämpas i enlighet med artikel 21 i den förordningen och som har
- fått vissa av de uppgifter som skall anges i deklarationerna enligt kapitel III från andra administrativa handlingar behöver inte kräva att dessa uppgifter skall finnas med i deklarationerna,
- fått alla de uppgifter som skall anges i deklarationerna enligt kapitel III från andra administrativa handlingar får undanta aktörerna i fråga från skyldigheten att lämna in deklarationerna.
Artikel 8
Vid utformningen av deklarationer enligt artiklarna 2 och 4 skall följande viner betraktas som "annat vin" vara vin som härrör från druvsorter som i medlemsstaternas klassificering i enlighet med artikel 19 i förordning (EG) nr 1493/1999, samtidigt för samma administrativa enhet anges som druvsorter för vinframställning och i förekommande fall som bordsdruvor, som druvsorter som är avsedda att torkas eller som sorter avsedda för framställning av vinsprit.
När det gäller den deklaration som avses i artikel 4 skall emellertid endast sådant vin betraktas som "annat vin" enligt första stycket som enbart skall användas för framställning av vinsprit med skyddad ursprungsbeteckning eller sådan obligatorisk destillation som avses i artikel 28 i förordning (EG) nr 1493/1999.
Artikel 9
De produktmängder som skall tas upp i de deklarationer som avses i artiklarna 2, 4 och 6 skall uttryckas i hektoliter vin. De mängder koncentrerad druvmust och rektifierad koncentrerad druvmust som skall tas upp i de deklarationer som avses i artikel 4 skall uttryckas i hektoliter.
Medlemsstaterna får dock föreskriva att mängderna skall uttryckas i deciton i stället för i hektoliter i de deklarationer som avses i artikel 2.
Medlemsstaterna får fastställa koefficienter för konvertering av mängder så att andra produkter kan uttryckas som hektoliter vin. Koefficienterna får anpassas efter olika objektiva kriterier som påverkar konverteringen. Medlemsstaterna skall meddela kommissionen koefficienterna samtidigt som det sammandrag lämnas in som avses i artikel 14.
Den mängd vin som skall anges i de produktionsdeklarationer som föreskrivs i artikel 4 skall vara den totala mängd som erhålls efter huvudjäsningen, inklusive vindruv.
Artikel 10
Denna förordning skall inte påverka medlemsstaternas bestämmelser om skörde-, produktions-, behandlingsoch/eller saluförings- eller lagerdeklarationer som är avsedda att ge mer fullständig information, i synnerhet genom att de omfattar en bredare krets av personer än de som avses i artiklarna 2, 4 och 6.
Artikel 11
1. De deklarationer som avses i artiklarna 2 och 4 skall lämnas senast den 10 december. Medlemsstaterna får emellertid fastställa ett eller flera tidigare datum. De får dessutom fastställa ett visst datum vid vilket de kvantiteter som innehas skall tas med i deklarationen.
2. De deklarationer som avses i artikel 6 skall lämnas senast den 10 september för de kvantiteter som innehas den 31 juli. Medlemsstaterna får emellertid fastställa ett eller flera tidigare datum.
Artikel 12
Personer som skall lämna in skörde-, produktions-, saluförings- och/eller behandlings- eller lagerdeklarationer och som inte har lämnat in dessa vid de tidpunkter som anges i artikel 11 skall, utom i fall av force majeure, inte omfattas av de åtgärder som föreskrivs i artiklarna 24, 29, 30, 34 och 35 i förordning (EG) nr 1493/1999 för innevarande och närmast därpå följande vinår.
Dock gäller att om de frister som avses i första stycket överskrids med högst fem arbetsdagar skall de belopp som skall utbetalas för innevarande vinår minskas med 15 %. Om fristerna överskrids med högst tio arbetsdagar skall beloppen minskas med 30 %.
Artikel 13
1. Personer som skall lämna in skörde-, produktions-, saluförings-, behandlings- eller lagerdeklarationer och som lämnar in deklarationer som de behöriga myndigheterna i medlemsstaterna finner ofullständiga eller oriktiga får endast omfattas av de åtgärder som avses i artiklarna 24, 29, 30, 34 och 35 i förordning (EG) nr 1493/1999 om de uppgifter som saknas eller som är oriktiga inte är avgörande för ett korrekt genomförande av åtgärderna i fråga.
2. Om medlemsstaternas behöriga myndigheter finner att de deklarationer som avses i denna förordning är ofullständiga eller oriktiga, och om de felaktiga eller ej införda uppgifterna är nödvändiga för en korrekt tillämpning av de åtgärder som avses i punkt 1 skall medlemsstaten, utom i fall av force majeure, tillämpa följande påföljder, utan att det påverkar nationella påföljder.
a) När det gäller de åtgärder som avses i artiklarna 24, 34 och 35 i förordning (EG) nr 1493/1999, skall stödet minskas med
- samma procentsats som det konstaterade felet om felet medför att den deklarerade volymen justeras med 5 % eller mindre,
- två gånger det konstaterade felets procentsats om felet medför att den deklarerade volymen justeras med mer än 5 % men högst 20 %.
Stöd skall inte betalas ut om felet medför att den deklarerade volymen justeras med mer än 20 %, vare sig för vinåret i fråga eller för det därpå följande vinåret.
Om den oriktighet som fastställts i deklarationen kan hänföras till uppgifter från andra aktörer eller anslutna vilkas namn finns med i de föreskrivna handlingarna och inte kan kontrolleras i förväg av deklaranten skall stödet endast minskas med procentsatsen för justeringen.
b) När det gäller de åtgärder som avses i artiklarna 29 och 30 i förordning (EEG) nr 1493/1999 skall det pris som destillatören skall betala till den deklarerande producenten, om det vin som levereras till destillation ännu inte har betalats, minskas i följande omfattning:
- Med samma procentsats som det konstaterade felet om felet medför att den deklarerade volymen justeras med 5 % eller mindre.
Dessa priser skall inte betalas om felet medför att den deklarerade volymen justeras med mer än 20 %, vare sig för vinåret i fråga eller för det därpå följande vinåret.
Om den oriktighet som fastställts i deklarationen kan hänföras till information från andra aktörer eller anslutna vilkas namn finns med i de föreskrivna handlingarna och inte kan kontrolleras i förväg av deklaranten skall priserna endast minskas med procentsatsen för justeringen.
De behöriga myndigheterna skall anpassa de stöd som skall utbetalas till destillatören i förhållande till det pris som betalats till producenten.
Artikel 14
Medlemsstaterna skall vid datum som möjliggör för de meddelanden enligt artikel 16 upprätta följande:
a) En sammanställning på nationell nivå av de produktionsdeklarationer som avses i artikel 4 i denna förordning och om sådana finns, också av de koefficienter som används för att konvertera volymer av andra produkter än vin uttryckta i deciton till hektoliter vin för de olika produktionsområdena.
b) En sammanställning på nationell nivå av de lagerdeklarationer som avses i artikel 6 i denna förordning.
c) En bedömning för pågående vinår av den volym vinprodukter som kan förväntas framställas i medlemsstaten.
d) En bedömning för pågående vinår av uppgifter som gör det möjligt att uppskatta de tillgängliga mängderna vinprodukter och deras användning i medlemsstaten.
e) En provisorisk försörjningsbalans för senast föregående vinår och en slutlig försörjningsbalans för det näst senaste vinåret.
Artikel 15
1. För prisnoteringarna skall medlemsstaterna, förutom de i vilka kapitlen I och II i avdelning II i förordning (EG) nr 1493/1999 inte tillämpas i enlighet med artikel 21 i den förordningen, definiera sammanhängande produktionsområden som omfattar flera mindre produktionsområden vars produktion är tillräckligt homogen.
2. För varje produktionsområde skall medlemsstaterna välja plats för prisnoteringen.
3. På de valda platserna skall var fjortonde dag priset på vita och röda bordsviner utan geografisk beteckning och den saluförda volymen av dessa viner noteras på lämpligt sätt.
4. Ovannämnda priser skall gälla en nettovara fritt producenten.
Artikel 16
1. Medlemsstaterna skall meddela kommissionen
a) senast den 15 september och den 30 november under innevarande vinår, en bedömning av den volym vinprodukter som kan förväntas framställas i medlemsstaten enligt artikel 14 c,
b) senast den 30 november, en sammanställning av lagerdeklarationerna enligt artikel 14 b,
c) senast den 30 november, de uppgifter som gör det möjligt att uppskatta de tillgängliga mängderna vinprodukter och deras användning i medlemsstaten enligt artikel 14 d,
d) den provisoriska försörjningsbalansen för senast föregående vinår senast den 15 november och den slutliga försörjningsbalansen för det näst senaste vinåret senast den 15 mars, enligt artikel 14 e; försörjningsbalanserna skall skickas till Eurostat, gemenskapens statistikkontor.
e) senast den 15 februari, en sammanställning av produktionsdeklarationerna enligt artikel 14 a, eller en preliminär sammanställning. I det senare fallet skall det slutliga resultatet meddelas senast den 15 april.
2. Medlemsstaterna skall meddela kommissionen
a) före den 1 augusti 2001:
- Definitionen av de fastställda produktionsområdena.
- En beräkning av produktionen under de fem senaste vinåren för de områden som samlats inom produktionsområdet.
- De platser som valts i varje produktionsområde för prisnotering.
- Bestämmelserna för prisnotering.
b) Från och med den 1 augusti 2001 skall medlemsstaterna varannan tisdag meddela kommissionen priser och volymer för saluförda produkter tillsammans med alla övriga uppgifter som bedöms vara till hjälp för att bedöma marknadsutvecklingen i produktionsområdet.
Artikel 17
Medlemsstaterna skall underrätta kommissionen om alla nya omständigheter av betydelse som i nämnvärd grad kan påverka den bedömning av tillgängliga mängder och deras användning som görs på grundval av den slutgiltiga informationen från tidigare år.
Artikel 18
Utöver att de används för statistiska ändamål används uppgifterna i deklarationerna även vid tillämpningen av förordning (EG) nr 1493/1999. Särskilt uppgifter om uppdelningen av produktionen i bordsvin, kvalitetsvin fso och annat vin avgör rättigheter och skyldigheter för producenterna vid tillämpning av den förordningen.
Artikel 19
Kommissionen ansvarar för att de uppgifter som mottas i enlighet med denna förordning sprids.
Artikel 20
Artikel 74.4 i förordning (EG) nr 1623/2000 skall ersättas med följande: "4. Interventionsorganet skall från producenten återvinna ett belopp som motsvarar en del eller hela det stöd som betalats ut till destillatören i de fall producenten inte uppfyller kraven i gemenskapens bestämmelser för destillationen i fråga, och orsaken är något av följande:
a) Producenten har inte lämnat in skörde-, produktions- eller lagerdeklarationen inom fastställda tidsfrister.
Det belopp som skall återvinnas fastställs enligt reglerna i artikel 12 i kommissionens förordning (EG) nr 1282/2001(7).
b) Producenten har lämnat in en deklaration enligt punkt a ovan som medlemsstatens behöriga myndigheter anser vara ofullständig eller felaktig, och de uppgifter som saknas eller är felaktiga anses vara av väsentlig betydelse för tillämpningen av den berörda åtgärden.
Det belopp söm skall återvinnas fastställs enligt reglerna i artikel 13 i förordning (EG) nr 1282/2001.
c) Producenten har inte fullgjort skyldigheterna i artikel 37 i förordning (EG) nr 1493/1999 och överträdelsen har konstaterats eller meddelats destillatören efter det att det lägsta priset har betalats på grundval av tidigare deklarationer.
Hela det stöd som har betalats ut till destillatören skall återvinnas."
Artikel 21
Upphävanden
Kommissionens förordning (EEG) nr 2396/84(8) och (EG) nr 1294/96(9) upphör att gälla.
Artikel 22
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1322/2001
av den 29 juni 2001
om ändring av bilagorna I och III i rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), senast ändrad genom kommissionens förordning (EG) nr 807/2001(2), särskilt artikel 6, 7 och 8 i denna, och
av följande skäl:
(1) I enlighet med förordning (EEG) nr 2377/90 måste gränsvärden för högsta tillåtna restmängder successivt fastställas för samtliga farmakologiskt verksamma substanser som används inom gemenskapen i veterinärmedicinska läkemedel som är avsedda att ges till livsmedelsproducerande djur.
(2) Gränsvärden bör fastställas först efter det att Kommittén för veterinärmedicinska läkemedel har granskat all relevant information beträffande säkerheten med restmängder av ämnet i fråga för den som konsumerar livsmedel med animaliskt ursprung samt restmängdernas påverkan på den industriella bearbetningen av livsmedel.
(3) Vid fastställandet av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemdel i livsmedel med animaliskt ursprung är det nödvändigt att ange de djurarter i vilka restmängder kan förekomma, vilka mängder som kan förekomma i var och en av de relevanta vävnaderna från det behandlade djuret (målvävnad) samt vilket slag av restmängd som är relevant vid övervakningen av restmängder (restmarkör).
(4) För kontroll av resthalter bör enligt tillämplig gemenskapslagstiftning gränsvärden vanligtvis fastställas för målvävnaderna lever eller njure. I den internationella handeln avlägsnas dock ofta lever och njure från slaktkroppen, och gränsvärden bör därför alltid fastställas även för muskel- eller fettvävnader.
(5) För veterinärmedicinska läkemedel som är avsedda för äggläggande fåglar, mjölkdjur eller honungsbin, måste gränsvärden även fastställas för ägg, mjölk eller honung.
(6) Florfenikol bör införas i bilaga I till förordning (EEG) nr 2377/90.
(7) För att möjliggöra komplettering av vetenskapliga studier, bör giltighetstiden för temporär MRL, tidigare definierad i bilaga III till förordning (EEG) nr 2377/90, förlängas för cefalonium, morantel och metamizol.
(8) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I och III till förordning (EEG) nr 2377/90 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1637/2001
av den 23 juli 2001
om ändring av rådets förordning (EEG) nr 3880/91 om avlämnande av statistikuppgifter om nominell fångst för medlemsstater som bedriver fiske i Nordatlantens östra del
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3880/91 av den 17 december 1991 om avlämnande av statistikuppgifter över nominell fångst för medlemsstater som bedriver fiske i Nordatlantens östra del(1), särskilt artikel 2.3 och artikel 4 i denna, och
av följande skäl:
(1) Vid det nionde sammanträdet med parterna i Konventionen om internationell handel med utrotningshotade arter av vilda djur och växter (CITES) 1994 krävdes att åtgärder för bevakning av uppgifter om fångster av och handel med arter av Elasmobranchii-fiskar (hajar och rockor) skulle vidtas av FN:s livsmedels- och jordbruksorganisation (FAO) och av regionala fiskeorganisationer.
(2) Vid sitt 87:e stadgeenliga sammanträde 1999 beslöt Internationella rådet för utnyttjande av havet (ICES) att uppta de artgrupper av Elasmobranchii-fiskar, som beskrivs i rapporten från arbetsgruppen om Elasmobranchii-arter, och uppmana FAO att införa dessa arter i sitt Statlant 27A-frågeformulär om fångststatistik för nordöstra Atlanten.
(3) ICES har utvidgat sin förteckning över de arter vilkas fångst i nordöstra Atlanten skall inläggas i ICES:s databas och där medlemsstaterna när det gäller dessa ytterligare arter således skall uppmuntras att lämna tillgänglig fångststatistik.
(4) I artikel 4.2 i förordning (EEG) nr 3880/91 föreskrivs att medlemsstaterna efter att i förväg ha inhämtat medgivande från Eurostat, får lämna uppgifter i annan form eller med annat medium än enligt vad som föreskrivs i bilaga IV till förordningen.
(5) Flera medlemsstater har begärt att få inlämna uppgifter i annan form eller med annat medium än enligt vad som som föreskrivs i bilaga IV till förordning (EG) nr 3880/91 (som motsvarar ovannämnda Statlant-frågeformulär).
(6) De åtgärder, som föreskrivs i denna förordning står i överensstämmelse med yttrandet från Ständiga kommittén för jordbruksstatistik inrättad genom rådets förordning 72/279/EEG(2).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till förordning (EEG) nr 3880/91 skall ersättas med bilaga I till denna förordning.
Artikel 2
Medlemsstaterna får inlämna uppgifter i enlighet med det format som specificeras i bilaga II till denna förordning.
Artikel 3
Denna förordning träder i kraft den tjugonde dagen efter det att den offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1660/2001
av den 16 augusti 2001
om ändring av förordning (EG) nr 1623/2000 om tillämpningsföreskrifter för rådets förordning (EG) nr 1493/1999 om den gemensamma organisationen av marknaden för vin, vad beträffar marknadsmekanismerna
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1493/1999 av 17 maj 1999 om den gemensamma organisationen av marknaden för vin(1), senast ändrad genom förordning (EG) nr 2826/2000(2), särskilt artiklarna 33 och 36 i denna, och
av följande skäl:
(1) I artikel 58 i kommissionens förordning (EG) nr 1623/2000 av den 25 juli 2000 om tillämpningsföreskrifter för rådets förordning (EG) nr 1493/1999 om den gemensamma organisationen av marknaden för vin, vad beträffar marknadsmekanismerna(3), senast ändrad genom förordning (EG) nr 1282/2001(4), föreskrivs vinproducenters skyldigheter vid levererans av resterande kvantiteter till destillerier. Erfarenheten visar att tidsfristen bör senareläggas.
(2) I artikel 63 föreskrivs inrättandet av en stödordning för destillation av vin till spritdrycker. Denna ordning tilllämpades första gången under vinåret 2000/2001. Mot bakgrund av de erfarenheter som gjorts under det första tillämpningsåret bör ändringar införas. Bland annat bör destillationen inledas senare på året och andelen av vinproducentens produktion som får gå till denna destillation bör sänkas. Dessutom bör ett slutdatum införas för destillation.
(3) I artiklarna 86-102 föreskrivs avsättningsregler för alkohol som innehas av interventionsorganen. Vissa sakfel bör rättas, bland annat bör priset för prover ändras. Vidare bör det för rektifieringsprodukter beviljas samma avvikelse för bioetanol som för nya industriella användningsområden.
(4) Förvaltningskommittén för vin har inte avgivit något yttrande inom den tid som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.!
Artikel 1
Förordning (EG) nr 1623/2000 ändras på följande sätt:
1. Artikel 58 första stycket skall ersättas med följande: "De producenter som omfattas av någon av skyldigheterna enligt artiklarna 45 och 52 i den här förordningen och som före den 15 juli innevarande vinår har levererat minst 90 % av sin ålagda kvantitet kan uppfylla denna skyldighet genom att leverera resterande kvantitet före ett datum som den behöriga nationella myndigheten skall fastställa, dock inte senare än den 31 juli påföljande vinår."
2. Artikel 63 skall ändras på följande sätt:
a) Punkterna 1 och 2 skall ersättas med följande: "1. För bordsvin och vin som lämpar sig för framställning av bordsvin skall destillationen enligt artikel 29 i förordning (EG) nr 1493/1999 börja från och med den 16 oktober varje vinår.
2. Kvantiteten bordsvin, och vin som lämpar sig för framställning av bordsvin, som varje producent får lämna till destillation, skall begränsas till 30 % av dennes maximiproduktion av dessa viner som deklarerats under de tre senaste vinåren, inklusive det innevarande om deklarationen redan lämnats. Om den ovan angivna procentsatsen tillämpas, skall den producerade mängden bordsvin vara den som anges som vin i kolumnen 'bordsvin' i produktionsdeklarationen enligt artikel 18.1 i förordning (EG) nr 1493/1999."
b) Följande punkt skall läggas till som punkt 10: "10. Det vin som levereras till destilleri skall destilleras senast den 30 september påföljande vinår."
3. Artikel 86 första stycket skall ersättas med följande: "Kommissionen skall enligt förfarandet i artikel 75 i förordning (EG) nr 1493/1999 kvartalsvis inleda flera anbudsinfordringar som var och en skall omfatta minst 50000 hektoliter vinalkohol, och kvartalsvis tillsammans högst 600000 hektoliter hundraprocentig alkohol, för export till vissa tredje länder för slutlig användning endast inom bränslesektorn."
4. Artikel 91.12 skall ersättas med följande: "12. Säkerheten för att garantera att alkoholen exporteras skall, av det interventionsorgan som innehar den, frisläppas för varje kvantitet som bevisligen har exporterats inom föreskriven tidsfrist. Om tidsfristen för export överskrids skall, genom undantag från artikel 23 i förordning (EEG) nr 2220/85, och utom i fall av force majeure, denna exportsäkerhet på 3 euro per hektoliter hundraprocentig alkoholvara förverkas
a) under alla förhållanden till 15 %,
b) per dag efter den överskridna exporttidsfristen till 0,33 % av återstående belopp, efter avdrag av de tidigare 15 %."
5. Artikel 95.2 andra och tredje styckerna skall ersättas med följande: "Alkohol i behållare som inte anges i meddelandena om anbudsinfordran och offentlig auktion, eller i det beslut av kommissionen som avses i artiklarna 83-93 i den här förordningen, skall inte omfattas av detta förbud.
Interventionsorgan som innehar alkohol kan, i synnerhet av logistikskäl, ersätta alkohol i de behållare som anges i medlemsstaternas meddelande enligt punkt 1 i den här artikeln med en annan alkohol, som är av samma typ eller som blandats med annan alkohol som levererats till interventionsorganet fram till dess att en uttagsorder utfärdas. Medlemsstaternas interventionsorgan skall meddela kommissionen om att alkoholen ersatts."
6. Artikel 98 skall ändras på följande sätt:
a) Punkt 1 skall ersättas med följande: "1. Från och med offentliggörandet av ett meddelande om anbudsförfarande och fram till sista dagen för inlämnande av anbud kan alla intresserade parter, mot betalning av 10 euro per liter, erhålla prover av den alkohol som bjuds ut. Kvantiteten per intresserad part får inte överstiga 5 liter per behållare. För avsättningen enligt delavsnitt III kan varuprovet erhållas, mot samma betalning, inom 30 dagar efter meddelandet om offentlig auktion."
b) Punkt 2 skall ersättas med följande: "2. Efter tidsfristen för inlämnande av anbud eller efter trettio dagar efter meddelandet om offentlig auktion
a) får anbudsgivare eller godkända företag enligt artikel 92 erhålla prover av den tilldelade alkoholen,
b) får de anbudsgivare som erbjudits en ersättningsmängd enligt artikel 83.3 i den här förordningen erhålla prover av den alkohol som erbjuds som ersättning.
Dessa prover kan fås från interventionsorganet mot betalning av 10 euro per liter, varvid kvantiteten skall begränsas till 5 liter per behållare."
7. Artikel 100.2 c skall ersättas med följande: "c) Beträffande alkohol som vid offentlig auktion tilldelas för nya industriella användningsområden i syfte att användas som bioetanol inom gemenskapens bränslesektor och som måste rektifieras före den slutliga användningen, skall en användning för de föreskrivna ändamålen anses vara fullständig när minst 90 % av de totala alkoholkvantiteter som avhämtats i samband med anbudsinfordran eller offentlig auktion har använts för ändamålen i fråga. Anbudstagaren, eller det godkända företaget, som accepterat att köpa upp alkohol skall informera kommissionen och interventionsorganet om kvantiteten, ändamålet och användningen av de produkter som erhålls genom rektifieringen. Förlusterna får emellertid inte överskrida gränserna enligt b ovan."
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1681/2001
av den 22 augusti 2001
om ändring av förordning (EG) nr 174/1999 om fastställande av särskilda tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 i fråga om exportlicenser och exportbidrag inom sektorn för mjölk och mjölkprodukter och av förordning (EG) nr 1498/1999 om tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 beträffande meddelanden mellan medlemsstaterna och kommissionen med avseende på mjölk och mjölkprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), senast ändrad genom förordning (EG) nr 1670/2000(2), särskilt artikel 26.3, artikel 30, artikel 31.14 och artikel 40 i denna, och
av följande skäl:
(1) I artikel 1 i kommissionens förordning (EG) nr 174/1999 av den 26 januari 1999 om fastställande av särskilda tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 i fråga om exportlicenser och exportbidrag inom sektorn för mjölk och mjölkprodukter(3), senast ändrad genom förordning (EG) nr 1370/2001(4), fastställs som generell regel att en exportlicens skall uppvisas vid all export av mjölkprodukter för vilken exportbidrag begärs. För att få en effektiv förvaltning av den inre marknaden för skummjölkspulver, en produkt för vilken interventionsåtgärder kan bli aktuella, är det nödvändigt att exportlicensen blir obligatorisk och att medlemsstaterna skall ha skyldighet att meddela kommissionen uppgifter om dessa licenser. Därför bör kommissionens förordning (EG) nr 1498/1999 av den 8 juli 1999 om tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 beträffande meddelanden mellan medlemsstaterna och kommissionen med avseende på mjölk och mjölkprodukter(5), senast ändrad genom förordning (EG) nr 732/2001(6), ändras.
(2) En rättelse bör göras av ett fel som insmugit sig i artikel 9 i förordning (EG) nr 174/1999.
(3) För mjölkprodukter beaktas inte innehållet av sackaros när grundbeloppet för bidraget för mjölkhalten är fastställt till noll. Denna bestämmelse bör utvidgas till att gälla även om det inte fastställts något bidrag för mjölkhalten.
(4) För slutliga licenser för export utan bidrag till Förenta staterna inom den tilläggskvot som är en följd av jordbruksavtalet inom ramen för GATT:s Uruguayrunda(7) (nedan kallat jordbruksavtalet) behöver ingen säkerhet ställas. För att se till att denna kvot i möjligaste mån utnyttjas fullt ut och att de licenser som utfärdats används, bör en säkerhet ställas.
(5) För att förenkla säkerheterna för de tillfälliga licenser som avses i artikel 20 är det lämpligt att justera säkerheterna för sådana licenser och att precisera hur säkerheterna för slutliga licenser skall fungera.
(6) Förvaltningskommittén för mjölk och mjölkprodukter har inte yttrat sig inom den tid som dess ordföranden har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 174/1999 ändras på följande sätt:
1. I artikel 1.1 skall följande stycke läggas till: "Genom undantag från första stycket skall emellertid en exportlicens uppvisas vid all export av sådana produkter som avses i bilaga I kategori II."
2. I artikel 9 skall led a ersättas med följande: "a) 5 % för produkter med KN-nummer 0405."
3. Artikel 16.3 andra stycket skall ersättas med följande: "Innehållet av sackaros skall emellertid inte beaktas om grundbeloppet för den mjölkhalt som avses i punkt 2 andra stycket är fastställt till noll, eller om det inte har fastställts något grundbelopp."
4. I artikel 20.2 andra stycket skall "9 euro" ersättas med "6 euro".
5. Artikel 20.10 skall ersättas med följande: "10. Före utgången av det år för vilket de tillfälliga licenserna utfärdats skall den berörda parten, även om det rör sig om delkvantiteter, ansöka om en slutlig exportlicens som skall utfärdas omedelbart, varvid den säkerhet som avses i punkt 2 skall höjas till det totalbelopp som föreskrivs i artikel 9 för de kvantiteter för vilka licenser tilldelas. I ansökan om slutlig licens och i licensen skall följande anges i fält 20: 'För export till Amerikas förenta stater: artikel 20 i förordning (EG) nr 174/1999.'
De slutliga licenserna gäller endast för sådan export som avses i punkt 1.
Säkerheten för den slutliga licensen får endast frisläppas mot uppvisande av det bevis som avses i artikel 35.5 i förordning (EG) nr 1291/2000(8)."
Artikel 2
Artikel 9.1 i förordning (EG) nr 1498/1999 skall ersättas med följande: "1. varje arbetsdag före kl. 18.00, utom för kvantiteter för vilka exportlicens begärts, antingen enligt artikel 18 eller artikel 19.5 i förordning (EG) nr 174/1999, eller för leveranser av livsmedelshjälp enligt artikel 10.4 i Uruguayrundans jordbruksavtal, översända uppgifter om följande:
a) De kvantiteter, fördelade efter nummer i exportbidragsnomenklaturen för mjölkprodukter och efter kod för bestämmelseort, för vilka licens har begärts samma dag,
i) som avses i artikel 1 i förordning (EG) nr 174/1999, med undantag för sådana produkter som avses i artikel 17 i den förordningen (kod för IDES-meddelanden: 1),
b) De kvantiteter, fördelade efter begäran, efter nummer i exportbidragsnomenklaturen för mjölkprodukter och efter kod för bestämmelseort, för vilka det samma dag begärts sådan tillfällig licens som avses i artikel 8 i förordning (EG) nr 174/1999, med angivande av sista dag för att lämna in anbud samt kvantiteten i anbudsinfordran, eller, om det rör sig om en anbudsinfordran som öppnats av de väpnade styrkorna i enlighet med artikel 36.1 c i kommissionens förordning (EG) nr 800/19991(1) i vilken någon kvantitet inte specificeras, med angivande av den beräknade kvantiteten, fördelad enligt vad som sägs ovan (kod för IDES-meddelande: 2).
c) De kvantiteter, fördelade efter nummer i exportbidragsnomenklaturen för mjölkprodukter och efter kod för bestämmelseort, för vilka sådana tillfälliga licenser som avses i artikel 8 i förordning (EG) nr 174/1999 slutligt utfärdats eller dragits in samma dag, med angivande av från vilket organ anbudsinfordran kommer, samt dessutom datum och kvantitet för den tillfälliga licensen.
d) I förekommande fall den justerade kvantiteten i en anbudsinfordran enligt b ovan."
Artikel 3
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Rådets förordning (EG) nr 2136/2001
av den 23 oktober 2001
om ändring av rådets förordning (EG) nr 723/97 om genomförande av medlemsstaternas åtgärdsprogram på området för kontroll av utgifterna för EUGFJ:s garantisektion
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2), och
av följande skäl:
(1) Enligt artikel 1 i förordning (EG) nr 723/97(3) skall gemenskapen delta i de kostnader som medlemsstaterna ådragit sig för att genomföra de nya åtgärdsprogram som följer av nya skyldigheter gentemot gemenskapen, vilka har godkänts av kommissionen och vars syfte är att förbättra strukturen hos och effektiviteten av kontrollen när det gäller utgifterna för EUGFJ:s garantisektion. Enligt artikel 4 i förordningen skall det finansiella bidraget från gemenskapen beviljas per kalenderår under en tid av fem år i följd räknat från år 1997. Det skall beviljas inom ramen för de årliga anslag som beviljas av budgetmyndigheten inom ramen för budgetplanen.
(2) Kommissionen har lämnat en rapport till rådet om tilllämpningen av förordning (EG) nr 723/97 under perioden 1997-2000. Av de utvärderingsrapporter som sammanställts av medlemsstaterna och de genomförda programmens effektivitet drar kommissionen slutsatsen att medlemsstaterna bör få fortsatt finansiellt bidrag för att genomföra programmen enligt artikel 1 i förordning (EG) nr 723/97.
(3) Särskilt eftersom nya dyra tekniska metoder har införts genom rådets förordning (EG) nr 1593/2000 av den 17 juli 2000 om ändring av förordning (EEG) nr 3508/92 om ett integrerat system för administration och kontroll av vissa stödsystem inom gemenskapen(4), i form av förbättringar av systemet för identifiering av jordbruksskiften med hjälp av GIS-system och digitala ortofotosystem, är ett bidrag från gemenskapen motiverat för att täcka en del av medlemsstaternas kostnader för de nya åtgärdsprogrammen inom detta område. För den juridiska tydlighetens skull bör därför sista strecksatsen i artikel 5 i förordning (EG) nr 723/97 strykas.
(4) Den period under vilken det finansiella bidraget från gemenskapen kan betalas bör därför förlängas med två år.
(5) Förordning (EG) nr 723/97 bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 723/97 ändras på följande sätt:
2. I första meningen i artikel 4.1 skall orden "fem år i följd" ersättas med orden "sju år i följd".
Kommissionens förordning (EG) nr 2601/2001
av den 28 december 2001
om komplettering av bilagan till förordning (EG) nr 2400/96 om upptagandet av vissa namn i Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar som föreskrivs i rådets förordning (EEG) nr 2081/92 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel(1), senast ändrad genom kommissionens förordning (EG) nr 2796/2000(2), särskilt artikel 6.3 och 6.4 i denna, och
av följande skäl:
(1) Spanien har i enlighet med artikel 5 i förordning (EEG) nr 2081/92 till kommissionen översänt en ansökan om registrering av "Manzana Reineta del Bierzo" som ursprungsbeteckning och en ansökan om registrering av "Salchichón de Vic" "Llonganissa de Vic" som geografisk beteckning.
(2) Det har i enlighet med artikel 6.1 i nämnda förordning konstaterats att de två ansökningarna är förenliga med den förordningen, särskilt eftersom de omfattar alla komponenter som avses i artikel 4.
(3) Inga invändningar enligt artikel 7 i förordning (EEG) nr 2081/92 har framställts till kommissionen till följd av offentliggörandet i Europeiska gemenskapernas officiella tidning(3) av de produktnamn som anges i bilagan till den här förordningen.
(4) Dessa produktnamn kan därför tas upp i Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar och därmed vara skyddade inom gemenskapen såsom skyddad ursprungsbeteckning eller skyddad geografisk beteckning.
(5) Bilagan till denna förordning kompletterar bilagan till kommissionens förordning (EG) nr 2400/96(4), senast ändrad genom förordning (EG) nr 2372/2001(5).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (EG) nr 2400/96 skall kompletteras med de produktnamn som anges i bilagan till denna förordning och dessa namn skall tas upp i Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar såsom skyddad ursprungsbeteckning (SUB) eller skyddad geografisk beteckning (SGU) i enlighet med artikel 6.3 i förordning (EEG) nr 2081/92.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens beslut
av den 4 februari 2002
(Text av betydelse för EES)
(2002/79/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 93/43/EEG av den 14 juni 1993 om livsmedelshygien(1), särskilt artikel 10.1 i detta, och
av följande skäl:
(1) Jordnötter som har sitt ursprung i eller försänds från Kina har vid ett flertal tillfällen visat sig innehålla alltför höga halter av aflatoxin B1 eller alltför hög total aflatoxinhalt.
(2) Vetenskapliga livsmedelskommittén har konstaterat att aflatoxin B1 även i extremt låga doser orsakar levercancer och dessutom är genotoxisk.
(3) I kommissionens förordning (EG) nr 194/97 av den 31 januari 1997 om fastställande av högsta tillåtna halt för vissa främmande ämnen i livsmedel(2), senast ändrad genom förordning (EG) nr 1566/1999(3), fastställs högsta tillåtna halter för vissa främmande ämnen i livsmedel, särskilt för aflatoxiner. Dessa gränsvärden har vida överskridits i prov tagna från jordnötter som har sitt ursprung i eller försänds från Kina.
(4) Detta utgör en allvarlig fara för folkhälsan inom gemenskapen. Det är därför nödvändigt att anta skyddsåtgärder på gemenskapsnivå.
(5) Den 8-21 maj 2001 besökte kommissionens kontor för livsmedels- och veterinärfrågor Kina för att bedöma de befintliga kontrollsystemen för att hindra aflatoxinkontaminering av jordnötter avsedda för export till Europeiska gemenskapen. Vid detta besök konstaterades bland annat att kontrollen av aflatoxinhalten i jordnötter var minimal såväl i produktionen som i den allmänna bearbetningen. Brister i laboratoriehanteringen konstaterades också. För att garantera ett fullgott skydd för folkhälsan bör därför särskilda villkor införas för jordnötter och produkter framställda av jordnötter som har sitt ursprung i eller försänds från Kina.
(6) Jordnötter och produkter framställda av jordnötter måste produceras, sorteras, hanteras, bearbetas, förpackas och transporteras under goda hygieniska förhållanden. Halterna av aflatoxin B1 och den totala aflatoxinhalten måste fastställas i prover som tas ur sändningar just innan de lämnar Kina.
(7) De kinesiska myndigheterna bör se till att alla sändningar av jordnötter som har sitt ursprung i eller försänds från Kina åtföljs av skriftlig dokumentation som anger under vilka förhållanden varorna producerats, sorterats, hanterats, bearbetats, förpackats och transporterats samt resultaten från en laboratorieanalys av halterna av aflatoxin B1 och den totala aflatoxinhalten i sändningen.
(8) Av resultaten från det ovannämnda besöket framgår att de kinesiska myndigheterna för närvarande inte kan garantera att provresultaten är tillförlitliga eller att certifieringen avser hela sändningen. Det är därför mycket tveksamt hur tillförlitliga intyg är som avser jordnötter med ursprung i Kina.
(9) För att skydda folkhälsan måste därför de behöriga myndigheterna i den importerande medlemsstaten ta prover på alla sändningar av jordnötter som har sitt ursprung i eller försänds från Kina och som importeras till Europeiska gemenskapen och analysera dessa prover med avseende på aflatoxinhalten, innan jordnötterna släpps ut på marknaden. Eftersom denna åtgärd tar en betydande del av medlemsstaternas kontrollresurser i anspråk, kommer resultaten av åtgärden att utvärderas efter en kort period och åtgärderna ändras vid behov.
(10) Ständiga livsmedelskommittén rådfrågades den 2 april 2001 och den 19 juli 2001.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Medlemsstaterna får inte importera produkter som tillhör nedanstående kategorier och som har sitt ursprung i eller försänds från Kina och är avsedda som livsmedel eller att användas som ingrediens i livsmedel, om inte sändningen åtföljs av resultaten av en officiell provtagning och analys samt av ett sådant hälsointyg som återges i bilaga I, ifyllt och undertecknat av en företrädare för den kinesiska myndigheten State Administration for Entry/Exit Inspection and Quarantine:
- Jordnötter som omfattas av KN-nummer 1202 10 90 eller 1202 20 00.
- Jordnötter som omfattas av KN-nummer 2008 11 94 (i förpackningar med en nettovikt på mer än 1 kg) eller 2008 11 98 (i förpackningar med en nettovikt på mindre än 1 kg).
- Rostade jordnötter som omfattas av KN-nummer 2008 11 92 (i förpackningar med en nettovikt på mer än 1 kg) och KN-nummer 2008 11 96 (i förpackningar med en nettovikt på mindre än 1 kg).
2. Sändningar får importeras till gemenskapen endast genom de införselplatser som anges i bilaga II.
3. Varje sändning skall märkas med samma beteckning som den som anges i hälsointyget och i den bifogade rapporten med resultaten från den officiella provtagningen och analysen som avses i punkt 1.
4. De behöriga myndigheterna i varje medlemsstat skall se till att handlingarna för importerade jordnötter som har sitt ursprung i eller försänds från Kina kontrolleras, för att garantera att de krav på hälsointyg och provresultat som avses i punkt 1 är uppfyllda.
5. Medlemsstaterna skall ta prover ur alla sändningar och analysera halterna av aflatoxin B1 och den totala aflatoxinhalten i sändningen innan denna släpps ut på marknaden från införselplatsen, och skall underrätta kommissionen om resultaten.
Artikel 2
Europaparlamentets beslut
av den 14 mars 2002
om ändring av Europaparlamentets beslut 94/262/EGKS, EG, Euratom om föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning
(2002/262/EG, EKSG, Euratom)
EUROPAPARLAMENTET HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 195.4,
med beaktande av Fördraget om upprättandet av Europeiska kol- och stålgemenskapen, särskilt artikel 20 d.4,
med beaktande av Fördraget om upprättandet av Europeiska kol- och stålgemenskapen, särskilt artikel 107 d.4,
med beaktande av Europaparlamentets resolution av den 17 november 2000 om ändring av Europaparlamentets beslut av den 9 mars 1994 om föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning(1),
med beaktande av kommissionens yttrande,
med rådets godkännande, och
av följande skäl:
(1) Enligt artikel 22.5 i budgetförordningen av den 21 december 1977 för Europeiska gemenskapernas allmänna budget(2) skall ombudsmannen vid tillämpningen av denna förordning behandlas som en institution.
(2) Genom rådets förordning (EG, EKSG, Euratom) nr 2673/1999 om ändring av budgetförordningen inrättades ett särskilt avsnitt för ombudsmannen i Europeiska unionens allmänna budget och i konsekvens med detta ändrades berörda bestämmelser i budgetförordningen.
(3) Det är därför nödvändigt att ändra beslut 94/262/EKSG, EG, Euratom och Europaparlamentet av den 9 mars 1994 om föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning(3) eftersom det i detta beslut föreskrivs att ombudsmannens budget skall utgöra bilaga till avsnitt I (Europaparlamentet) i Europeiska gemenskaperna allmänna budget.
(4) Följaktligen bör artiklarna 12 och 16 i detta beslut utgå.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artiklarna 12 och 16 i beslut 94/262/EKSG, EG och Euratom skall utgå.
Artikel 2
Kommissionens beslut
av den 29 juli 2002
om att bilda Europeiska gruppen av regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation
(Text av betydelse för EES)
(2002/627/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, och
av följande skäl:
(1) Ett nytt regelverk för nät och tjänster inom området elektronisk kommunikation har inrättats i enlighet med följande direktiv från Europaparlamentet och rådet: 2002/21/EG av den 7 mars 2002 om ett gemensamt regelverk för elektroniska kommunikationsnät och kommunikationstjänster ("ramdirektivet")(1), 2002/19/EG av den 7 mars 2002 om tillträde till och samtrafik mellan elektroniska kommunikationsnät och tillhörande utrustning ("samtrafikdirektivet")(2), 2002/20/EG av den 7 mars 2002 om auktorisation för elektroniska kommunikationsnät och kommunikationstjänster ("tillståndsdirektivet")(3) samt 2002/22/EG av den 7 mars 2002 om samhällsomfattande tjänster och användares rättigheter avseende elektroniska kommunikationsnät och kommunikationstjänster ("direktivet om samhällsomfattande tjänster")(4).
(2) För genomförandet av de regleringsuppgifter som anges i dessa direktiv har nationella regleringsmyndigheter inrättats i samtliga medlemsstater, och dessa myndigheter skall anmälas till kommissionen i enlighet med artikel 3.6 i ramdirektivet. Enligt ramdirektivet skall medlemsstaterna också garantera den oberoende ställningen hos sina nationella regleringsmyndigheter genom att sörja för att de hålls rättsligt åtskilda från och verksamhetsmässigt oberoende av alla organisationer som tillhandahåller nät, utrustning eller tjänster för elektronisk kommunikation. Medlemsstater som behåller äganderätten till eller kontrollen över företag som tillhandahåller elektroniska kommunikationsnät eller kommunikationstjänster skall också sörja för att en praktiskt fungerande organisatorisk åtskillnad görs mellan regleringsverksamhet och sådan verksamhet som har samband med ägande eller kontroll.
(3) De sätt på vilka de nationella regleringsmyndigheternas ansvar och uppgifter är fastlagda i detalj skiljer sig åt mellan medlemsstaterna, men gemensamt är att alla har minst en nationell regleringsmyndighet som har som uppdrag att tillämpa bestämmelserna - särskilt dem som rör den löpande tillsynen över marknaden - när de väl har omsatts i nationell lagstiftning.
(4) Att bestämmelserna tillämpas på ett enhetligt sätt i alla medlemsstater är av avgörande betydelse för att man skall lyckas med att utveckla en gemensam marknad för nät och tjänster inom området elektronisk kommunikation. I det nya regelverket fastställs mål och ramar för de nationella regleringsmyndigheternas åtgärder, samtidigt som de får handlingsutrymme för att inom bestämda områden väga in nationella särdrag vid tillämpningen av bestämmelserna.
(5) En europeisk grupp av regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation (nedan kallad gruppen) bör bildas. Avsikten är att den skall fungera som förmedlande länk för samråd med och experthjälp åt kommissionen inom området elektronisk kommunikation.
(6) Gruppen bör fungera som en förmedlande länk mellan nationella regleringsmyndigheter och kommissionen på sådant sätt att den bidrar till den inre marknadens utveckling. I gruppen bör medlemsstaterna också kunna bedriva öppet redovisat samarbete med nationella regleringsmyndigheter och kommissionen för att på så sätt sörja för att regelverket för nät och tjänster inom området elektronisk kommunikation tillämpas på ett enhetligt sätt i alla medlemsstater.
(7) Gruppen bör fungera som ett organ som bistår kommissionen med utredningar, diskussioner och rådgivning inom området elektronisk kommunikation, däribland även i frågor som rör genomförande och revidering av rekommendationer avseende relevanta produkt- och tjänstemarknader samt när det gäller att utforma beslutet om transnationella marknader.
(8) Gruppen bör bedriva nära samarbete med den kommunikationskommitté som inrättats i enlighet med ramdirektivet. Gruppen bör verka på ett sådant sätt så att den inte inkräktar på kommitténs arbete.
(9) Verksamheten bör samordnas med arbetet i den radiospektrumkommitté som inrättats i enlighet med Europaparlamentets och rådets beslut nr 676/2002/EG av den 7 mars 2002 om ett regelverk för radiospektrumpolitiken i Europeiska gemenskapen (det s.k. radiospektrumbeslutet)(5), i den grupp för radiospektrumpolitik som inrättats i enlighet med kommissionens beslut 2002/622/EG av den 26 juli 2002 om inrättande av en grupp för radiospektrumpolitik(6) samt i den kontaktkommitté för television utan gränser som inrättats i enlighet med Europaparlamentets och rådets direktiv 97/36/EG av den 30 juni 1997 om samordning av vissa bestämmelser som fastställts i medlemsstaternas lagar och andra författningar om utförandet av sändningsverksamhet för television(7).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Innehåll
Härmed inrättas en rådgivande grupp som skall bestå av oberoende nationella regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation och vars namn skall vara Europeiska gruppen av regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation (nedan kallad gruppen).
Artikel 2
Definition
I detta direktiv avses med regleringsmyndighet: myndighet som inrättats i respektive medlemsstat för övervakning av den löpande tolkningen och tillämpningen av bestämmelserna i de direktiv som rör elektroniska kommunikationsnät och elektroniska kommunikationstjänster såsom de är definierade i ramdirektivet.
Artikel 3
Arbetsuppgifter
Gruppen skall vara rådgivare till kommissionen och bistå den när det gäller att befästa den inre marknaden för nät och tjänster inom området elektronisk kommunikation.
Gruppen skall fungera som en förmedlande länk mellan nationella regleringsmyndigheter och kommissionen på sådant sätt att den bidrar till den inre marknadens utveckling och till att regelverket för nät och tjänster inom området elektronisk kommunikation tillämpas på ett enhetligt sätt i alla medlemsstater.
Artikel 4
Ledamöter
Gruppen skall vara sammansatt av cheferna för respektive medlemsstaters nationella regleringsmyndigheter eller av deras ombud.
Kommissionen skall vara företrädd på en nivå som är avpassad till gruppens uppgifter, och kommissionen skall även tillhandahålla ett sekretariat för gruppens behov.
Artikel 5
Arbetsordning
Gruppen skall - på eget initiativ eller på kommissionens begäran - ge råd till och bistå kommissionen i alla frågor som rör nät och tjänster inom området elektronisk kommunikation.
Gruppen skall inom sig utse en ordförande. Verksamheten får i tillämpliga fall organiseras så att den fördelas på undergrupper och sakkunniggrupper.
Ordföranden skall kalla gruppen till sammanträde efter överenskommelse med kommissionen.
Gruppen skall enhälligt anta sin arbetsordning eller, om enhällighet inte kan uppnås, genom omröstning med två tredjedels majoritet, varvid varje medlemsstat har en röst, och arbetsordningen skall godkännas av kommissionen.
Kommissionen skall vara företrädd vid gruppens samtliga möten och ha möjlighet att närvara vid samtliga de möten som undergrupperna och sakkunniggrupperna håller.
Sakkunniga från EES-länder samt från kandidatländerna för anslutning till Europeiska unionen får delta som observatörer i gruppen. Gruppen får kalla andra sakkunniga och observatörer att närvara vid sina möten.
Artikel 6
Samråd
Gruppen skall i ett tidigt skede genomföra omfattande samråd med marknadsaktörer, konsumenter och slutförbrukare på ett sätt som garanterar öppenhet och insyn.
Artikel 7
Sekretess
Utan att det påverkar tillämpningen av bestämmelserna i artikel 287 i fördraget, skall gruppens ledamöter, liksom dess observatörer och alla andra personer - i de fall kommissionen upplyser dem om att de rådgivande yttranden som begärts in eller de frågor väckts är av konfidentiell art - vara förpliktade att inte röja uppgifter som har kommit till deras kännedom genom arbetet i gruppen, dess undergrupper eller sakkunniggrupper. Kommissionen får i sådana fall besluta att enbart gruppens ledamöter får närvara vid mötena i fråga.
Artikel 8
Årsberättelse
Gruppen skall lämna en årsberättelse över sin verksamhet till kommissionen. Kommissionen skall överlämna årsberättelsen till Europaparlamentet och rådet, i tillämpliga fall med sina kommentarer bifogade.
Artikel 9
Ikraftträdande
Detta beslut träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Kommissionens beslut
av den 21 november 2002
om ändring av beslut 94/652/EG om uppdatering av inventeringen och uppgifterna inom ramen för medlemsstaternas samarbete vid den vetenskapliga granskningen av livsmedelsfrågor
(2002/916/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 93/5/EEG av den 25 februari 1993 om hjälp till kommissionen och samarbete från medlemsstaternas sida vid den vetenskapliga granskningen av livsmedelsfrågor(1), särskilt artikel 3.2 fjärde strecksatsen i detta, och
av följande skäl:
(1) I kommissionens beslut 94/458/EG(2) fastställs bestämmelser om den administrativa organisationen av samarbetet vid den vetenskapliga granskningen av livsmedelsfrågor.
(2) I kommissionens beslut 94/652/EG(3), senast ändrat genom beslut 2001/773/EG(4), fastställs inventeringen och fördelningen av uppgifterna inom ramen för medlemsstaternas samarbete vid den vetenskapliga granskningen av livsmedelsfrågor.
(3) Uppdateringen av inventeringen av uppgifterna bör ta hänsyn till behovet av människors hälsa inom gemenskapen och till gemenskapslagstiftningens krav inom livsmedelssektorn.
(4) Uppgifterna bör fördelas med hänsyn till den vetenskapliga kompetens och de resurser som finns i medlemsstaterna och särskilt de institut som kommer att delta i det vetenskapliga samarbetet.
(5) Beslut 94/652/EG bör ändras i enlighet med detta.
(6) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga livsmedelskommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till beslut 94/652/EG ersätts med texten i bilagan till det här beslutet.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Europaparlamentets och rådets direktiv 2002/14/EG
av den 11 mars 2002
om inrättande av en allmän ram för information till och samråd med arbetstagare i Europeiska gemenskapen
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 137.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
med beaktande av Regionkommitténs yttrande(3),
i enlighet med förfarandet i artikel 251(4), på grundval av det gemensamma utkast som förlikningskommittén godkände den 23 januari 2002 och
av följande skäl:
(1) Enligt artikel 136 i fördraget skall gemenskapen och medlemsstaterna särskilt ha som mål att främja en dialog mellan arbetsmarknadens parter.
(2) I punkt 17 i gemenskapsstadgan om arbetstagares grundläggande sociala rättigheter föreskrivs bland annat att "information till, samråd med och deltagande av arbetstagare måste utvecklas på ett lämpligt sätt med hänsyn till gällande förfaranden i de olika medlemsstaterna".
(3) Kommissionen har samrått med arbetsmarknadens parter på gemenskapsnivå om den möjliga inriktningen av en gemenskapsåtgärd för information till och samråd med arbetstagare i företag inom gemenskapen.
(4) Kommissionen ansåg efter detta samråd att en gemenskapsåtgärd var önskvärd och samrådde på nytt med arbetsmarknadens parter om det planerade förslagets innehåll; arbetsmarknadens parter har inkommit med yttranden till kommissionen.
(5) Efter denna andra samrådsetapp har arbetsmarknadens parter inte underrättat kommissionen om att de önskar inleda det förfarande som kan leda till att ett avtal ingås.
(6) De rättsliga ramar som finns på nationell nivå och på gemenskapsnivå för att säkerställa arbetstagarnas deltagande i företagets angelägenheter och i de beslut som berör dem har inte alltid kunnat förhindra att ingripande beslut som påverkar arbetstagarna har fattats och offentliggjorts utan att lämpliga förfaranden för information och samråd ägt rum i förväg.
(7) Det finns behov av att förstärka den sociala dialogen och öka det ömsesidiga förtroendet inom företagen för att göra det lättare att föregripa risker, göra arbetsorganisationen mer flexibel och underlätta arbetstagarnas tillgång till utbildning inom företaget under trygga förhållanden, öka arbetstagarnas medvetenhet om behoven av anpassning, stimulera arbetstagarna att medverka i åtgärder och insatser för att öka deras anställbarhet, främja arbetstagarnas medverkan i företagets verksamhet och framtid samt stärka företagets konkurrenskraft.
(8) Det finns i synnerhet ett behov av att främja och stärka informationen och samrådet om den rådande situationen och den förväntade utvecklingen av sysselsättningen inom företaget och, när arbetsgivaren bedömer att sysselsättningen i företaget kan komma att hotas, om vilka eventuella föregripande åtgärder som planeras, i synnerhet i form av utbildning och kompetensutveckling för arbetstagarna, för att motverka den negativa utvecklingen eller mildra dess följder samt för att öka anställbarheten och anpassningsförmågan hos de arbetstagare som kan komma att påverkas.
(9) Det är en förutsättning att information ges och samråd äger rum i god tid i förväg om företagens omstrukturering och anpassning till de nya villkor som globaliseringen av ekonomin skapar skall kunna bli framgångsrik, bland annat genom att nya former för arbetets organisation utvecklas.
(10) Gemenskapen har utarbetat och genomfört en sysselsättningsstrategi som vilar på begreppen "föregripande", "förebyggande" och "anställbarhet", som skall bli hörnstenar i all offentlig politik som kan inverka positivt på sysselsättningen, även den som utformas inom företagen, genom en intensifiering av dialogen mellan arbetsmarknadens parter för att främja sådana förändringar som är förenliga med bibehållandet av det prioriterade sysselsättningsmålet.
(11) Den inre marknaden måste utvecklas på ett balanserat sätt med bibehållande av de viktiga värderingar som ligger till grund för våra samhällen, och genom att alla medborgare får del av den ekonomiska utvecklingen.
(12) Inträdet i den tredje etappen av den ekonomiska och monetära unionen har medfört en fördjupad och ökad konkurrens på europeisk nivå. Detta kräver att stödåtgärder vidtas på nationell nivå.
(13) Gemenskapens och medlemsstaternas nuvarande rättsliga ramar för information till och samråd med arbetstagare är ofta i alltför hög grad inriktade på hur man hanterar förändringsprocesser i efterhand, samtidigt som de bortser från de ekonomiska aspekterna av besluten och inte främjar ett verkligt föregripande av sysselsättningsutvecklingen i företag eller förebyggande av risker.
(14) Hela denna politiska, ekonomiska, sociala och rättsliga utveckling gör det nödvändigt att anpassa den befintliga rättsliga ramen inom vilken de rättsliga och praktiska instrument som gör det möjligt att utöva rätten till information och samråd föreskrivs.
(15) Detta direktiv påverkar inte de nationella system inom vilkas ram det konkreta utövandet av denna rättighet förutsätter en kollektiv viljeyttring från rättsinnehavarnas sida.
(16) Detta direktiv påverkar inte de system som föreskriver direkt deltagande av arbetstagarna, under förutsättning att dessa fortfarande har möjlighet att utöva rätten till information och samråd genom sina representanter.
(17) Eftersom målen för den planerade åtgärden, såsom den beskrivs ovan, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna, eftersom syftet är att inrätta en ram för information till och samråd med arbetstagare, vilken är anpassad till de nya europeiska förutsättningar som beskrivs ovan, och därför på grund av den planerade åtgärdens omfattning och verkningar bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
(18) Denna allmänna ram har till syfte att fastställa minimiföreskrifter som skall tillämpas i hela gemenskapen men den hindrar inte medlemsstaterna från att anta bestämmelser som är förmånligare för arbetstagarna.
(19) Denna allmänna ram bör också syfta till att undvika sådana administrativa, ekonomiska och rättsliga förpliktelser som kan motverka etableringen och utvecklingen av små och medelstora företag. Det förefaller därför rimligt att enligt medlemsstaternas val begränsa tillämpningsområdet för detta direktiv till företag med minst 50 arbetstagare eller till driftställen med minst 20 arbetstagare.
(20) Detta tar hänsyn till och påverkar inte andra nationella åtgärder och förfaranden som syftar till att främja en social dialog inom företag som inte omfattas av detta direktiv, och inom den offentliga förvaltningen
(21) Emellertid bör medlemsstater där det inte finns något lagstadgat system för information till och samråd med arbetstagare eller arbetstagarrepresentanter ha möjlighet att under en övergångsperiod ytterligare begränsa tillämpningsområdet för detta direktiv vad gäller antalet anställda.
(22) Gemenskapsramen för information till och samråd med arbetstagare bör i så hög grad som möjligt begränsa de bördor som läggs på företagen eller driftsställena men likväl säkerställa ett effektivt utövande av rättigheterna.
(23) Målet i detta direktiv uppnås genom inrättandet av en allmän ram med principer, definitioner och villkor för informationen och samrådet, som medlemsstaterna skall respektera och anpassa i förhållande till sina nationella förutsättningar, där det vid behov säkerställs att arbetsmarknadens parter får en ledande roll genom att de får rätt att genom avtal fritt fastställa de arrangemang för information och samråd som bäst överensstämmer med deras behov och önskemål.
(24) Man bör undvika att påverka vissa specifika regler om information till och samråd med arbetstagare i vissa nationella lagstiftningar, vilka gäller företag och driftställen som ägnar sig åt politik, yrkessammanslutningars verksamhet, religiös verksamhet, välgörenhet, utbildning, vetenskap, konst, information eller opinionsbildning.
(25) Företagen och driftställena bör skyddas mot att viss särskilt känslig information lämnas ut.
(26) Arbetsgivaren bör ges möjlighet att underlåta att informera och samråda, när detta skulle innebära allvarlig skada för företaget eller driftstället eller när han omedelbart måste hörsamma en anvisning som en övervaknings- eller tillsynsmyndighet givit honom.
(27) Information och samråd innebär rättigheter och skyldigheter för arbetsmarknadens parter på företags- eller driftställenivå.
(28) Administrativa eller rättsliga förfaranden och sanktioner som är effektiva och avskräckande samt står i proportion till hur allvarlig övertädelsen är bör tillämpas när skyldigheterna i detta direktiv inte uppfylls.
(29) Detta direktiv bör inte påverka andra mer specifika bestämmelser i rådets direktiv 98/59/EG av den 20 juli 1998 om tillnärmning av medlemsstaternas lagstiftning om kollektiva uppsägningar(5) och i rådets direktiv 2001/23/EG av den 12 mars 2001 om tillnärmning av medlemsstaternas lagstiftning om skydd för arbetstagares rättigheter vid överlåtelse av företag, verksamheter eller delar av företag eller verksamheter(6).
(30) Övriga rättigheter till information och samråd, inklusive de rättigheter som följer av rådets direktiv 94/45/EG av den 22 september 1994 om inrättandet av ett europeiskt företagsråd eller ett förfarande i gemenskapsföretag och grupper av gemenskapsföretag för information till och samråd med arbetstagare(7), bör inte påverkas av detta direktiv.
(31) Genomförandet av detta direktiv bör inte anses vara ett tillräckligt skäl för att rättfärdiga en sänkning av arbetstagarnas allmänna skyddsnivå på det område som omfattas av direktivet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte och principer
1. Detta direktiv syftar till att inrätta en allmän ram med minimikrav avseende arbetstagarnas rätt till information och samråd i företag eller driftställen inom gemenskapen.
2. Formerna för information och samråd skall fastställas och genomföras i enlighet med nationell lagstiftning och den praxis för relationerna mellan arbetsmarknadens parter som finns i de enskilda medlemsstaterna på ett sådant sätt att ändamålet med desamma säkerställs.
3. När formerna för information eller samråd fastställs och genomförs, skall arbetsgivaren och arbetstagarrepresentanterna arbeta i samförståndsanda med respekt för varandras ömsesidiga rättigheter och skyldigheter samt med beaktande av såväl företagets eller driftställets intressen som arbetstagarnas intressen.
Artikel 2
Definitioner
I detta direktiv avses med
a) företag: offentligt eller privat företag som bedriver ekonomisk verksamhet med eller utan vinstsyfte och som är beläget inom medlemsstaternas territorium,
b) driftställe: en verksamhetsenhet som definieras enligt nationell lagstiftning och nationell praxis där ekonomisk verksamhet som inbegriper mänskliga och materiella resurser bedrivs kontinuerligt och som är belägen inom en medlemsstats territorium,
c) arbetsgivare: en fysisk eller juridisk person som är part i ett anställningsavtal eller anställningsförhållande gentemot en arbetstagare i enlighet med nationell lagstiftning och nationell praxis,
d) arbetstagare: varje person som i den berörda medlemsstaten åtnjuter skydd som arbetstagare inom ramen för den nationella arbetslagstiftningen och enligt nationell praxis,
e) arbetstagarrepresentanter: företrädare för arbetstagare enligt definitionen i nationell lagstiftning och/eller nationell praxis,
f) information: arbetsgivarens överlämnande av uppgifter till arbetstagarrepresentanterna som gör det möjligt för dem att sätta sig in i vad den behandlade frågan avser och att granska densamma,
g) samråd: diskussion och upprättande av en dialog mellan arbetstagarrepresentanterna och arbetsgivaren.
Artikel 3
Räckvidd
1. I enlighet med medlemsstaternas val skall detta direktiv tillämpas på
a) företag som i en medlemsstat sysselsätter minst 50 arbetstagare, eller
b) driftställen som i en medlemsstat sysselsätter minst 20 arbetstagare.
Medlemsstaterna skall själva besluta om hur tröskelvärdena för anställda arbetstagare skall beräknas.
2. I enlighet med principerna och målen i detta direktiv får medlemsstaterna fastställa särskilda bestämmelser, som skall tillämpas på företag eller driftställen som direkt och huvudsakligen ägnar sig åt politik, yrkessammanslutningars verksamhet, religiös verksamhet, välgörenhet, utbildning, vetenskap, konst, information eller opinionsbildning, under förutsättning att sådana bestämmelser redan förekommer i nationell lagstiftning vid det datum då detta direktiv träder i kraft.
3. Medlemsstaterna får göra undantag från detta direktiv genom särskilda bestämmelser för besättningar på fartyg som trafikerar öppet hav.
Artikel 4
Former för information och samråd
1. I enlighet med principerna i artikel 1 och utan att det påverkar tillämpningen av gällande bestämmelser och/eller praxis som är mer gynnsamma för arbetstagarna, skall medlemsstaterna besluta om formerna för rätt till information och samråd på lämplig nivå i enlighet med denna artikel.
2. Information och samråd skall omfatta följande:
a) Information om den senaste och den förväntade utvecklingen av företagets eller driftställets verksamhet och ekonomiska situation.
b) Information och samråd om situationen, strukturen och den förväntade utvecklingen när det gäller sysselsättningen i företaget eller driftstället samt om eventuella föregripande åtgärder som planeras, bland annat vid hot mot sysselsättningen.
c) Information och samråd om beslut som kan medföra väsentliga förändringar i arbetsorganisationen eller anställningsavtalen, inklusive de beslut som avses i de gemenskapsbestämmelser som anges i artikel 9.1.
3. Informationen skall överlämnas vid ett sådant tillfälle, på ett sådant sätt och med ett sådant innehåll som gör det möjligt för särskilt arbetstagarrepresentanterna att granska informationen på ett adekvat sätt och vid behov förbereda samråd.
4. Samråd skall äga rum
a) med säkerställande av att tillfället, sättet och innehållet är lämpligt,
b) på den lednings- och representationsnivå som är relevant med hänsyn till den fråga som behandlas,
c) på grundval av de uppgifter som arbetsgivaren lämnat i enlighet med artikel 2 f) och det yttrande som arbetstagarrepresentanterna har rätt att avge,
d) på ett sådant sätt som gör det möjligt för arbetstagarrepresentanterna att sammanträda med arbetsgivaren och få motiverade svar på eventuella yttranden,
e) i syfte att söka nå en överenskommelse när det gäller de beslut som omfattas av arbetsgivarens befogenheter och som avses i punkt 2 c).
Artikel 5
Avtalsreglerad information och avtalsreglerat samråd
Medlemsstaterna får ge arbetsmarknadens parter tillåtelse att på lämplig nivå, inbegripet på företags- eller driftställesnivå, fritt och när som helst genom avtal fastställa formerna för information till och samråd med arbetstagare. Dessa avtal och de avtal som redan finns vid den tidpunkt som anges i artikel 11 samt alla därpå följande förnyelser av sådana avtal får på de villkor och med de begränsningar som fastställs av medlemsstaterna innehålla bestämmelser som avviker från bestämmelserna i artikel 4, om de överensstämmer med principerna i artikel 1.
Artikel 6
Konfidentiell information
1. Medlemsstaterna skall på de villkor och med de begränsningar som fastställs i nationell lagstiftning föreskriva att de arbetstagarrepresentanter och experter som eventuellt biträder dem inte har rätt att för arbetstagare eller tredje man röja information som de i företagets eller driftställets legitima intresse uttryckligen fått i förtroende. Denna förpliktelse skall fortsätta att gälla oavsett var experterna eller företrädarna befinner sig, även efter det att deras mandatperiod har löpt ut. En medlemsstat kan emellertid tillåta arbetstagarrepresentanter eller någon som biträder dem att vidarebefordra konfidentiell information till arbetstagare eller tredje man som är bundna av tystnadsplikt.
2. I särskilda fall och på de villkor och med de begränsningar som fastställs i nationell lagstiftning skall medlemsstaterna föreskriva att arbetsgivaren inte är skyldig att lämna ut sådan information eller inleda sådant samråd som utifrån objektiva kriterier skulle skada företaget eller driftstället eller vara till allvarligt förfång för dess verksamhet.
3. Utan att det påverkar befintliga nationella förfaranden skall medlemsstaterna säkerställa att det finns tillgång till rättsligt eller administrativt överklagandeförfarande i de fall arbetsgivaren hävdar att informationen är konfidentiell eller inte lämnar ut information i enlighet med punkt 1 och 2. De får dessutom införa förfaranden som säkerställer att den berörda informationen förblir konfidentiell.
Artikel 7
Skydd för arbetstagarrepresentanterna
Medlemsstaterna skall se till att arbetstagarrepresentanterna, när de utför sina uppdrag, får tillräckligt skydd och tillräckliga garantier, så att de på ett adekvat sätt kan utföra sina uppgifter.
Artikel 8
Tillvaratagande av rättigheterna
1. Medlemsstaterna skall föreskriva lämpliga åtgärder för de fall då arbetsgivaren eller arbetstagarrepresentanterna inte följer detta direktiv. De skall särskilt se till att det finns administrativa eller rättsliga förfaranden för att säkerställa att de skyldigheter som följer av detta direktiv iakttas.
2. Medlemsstaterna skall föreskriva lämpliga påföljder, som skall tillämpas när arbetsgivaren eller arbetstagarrepresentanterna överträder bestämmelserna i detta direktiv. Dessa påföljder skall vara effektiva, proportionella och avskräckande.
Artikel 9
Förhållandet mellan detta direktiv och andra bestämmelser på gemenskapsnivå och nationell nivå
1. Detta direktiv skall inte påverka tillämpningen av de särskilda förfaranden för information och samråd som avses i artikel 2 i direktiv 98/59/EG och i artikel 7 i direktiv 2001/23/EG.
2. Detta direktiv skall inte påverka de bestämmelser som antagits i enlighet med direktiv 94/45/EG och direktiv 97/74/EG.
3. Detta direktiv skall inte påverka övriga gällande rättigheter till information, samråd och medverkan enligt nationell lagstiftning.
4. Genomförandet av detta direktiv skall inte utgöra något tillräckligt skäl för tillbakagång i förhållande till den nuvarande situationen i medlemsstaterna och i förhållande till arbetstagarnas allmänna skyddsnivå på det område som omfattas av direktivet.
Artikel 10
Övergångsbestämmelser
Om det i en medlemsstat, vid den tidpunkt då detta direktiv träder i kraft, varken finns något allmänt, varaktigt och lagstadgat system för information till och samråd med arbetstagare eller något allmänt, varaktigt och lagstadgat system för arbetstagarrepresentation på arbetsplatsen, genom vilket de anställda kan företrädas, får denna medlemsstat, trots vad som sägs i artikel 3, såvitt avser detta ändamål begränsa tillämpningen av de nationella genomförandebestämmelserna för direktivet till
a) företag med minst 150 anställda eller driftställen med minst 100 anställda till och med den 23 mars 2007, och
b) företag med minst 100 anställda eller driftställen med minst 50 anställda under det år som följer efter den tidpunkt som anges i a).
Artikel 11
Genomförande av direktivet
1. Medlemsstaterna skall anta de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 23 mars 2005 eller se till att arbetsmarknadens parter inför de nödvändiga bestämmelserna genom avtal, varvid medlemsstaterna skall var skyldiga att vidta alla nödvändiga åtgärder för att alltid kunna garantera de resultat som införs genom detta direktiv. De skall genast underrätta kommissionen om detta.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 12
Översyn av kommissionen
Senast den 23 mars 2007 skall kommissionen i samråd med medlemsstaterna och arbetsmarknadens parter på gemenskapsnivå se över tillämpningen av detta direktiv och vid behov föreslå nödvändiga ändringar.
Artikel 13
Ikraftträdande
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Artikel 14
Adressater
Detta direktiv riktar sig till medlemsstaterna.
Europaparlamentets och rådets direktiv 2002/61/EG
av den 19 juli 2002
om ändring för nittonde gången av rådets direktiv 76/769/EEG om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar) (azofärger)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 95 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Arbetet med att upprätta den inre marknaden bör stegvis förbättra livskvaliteten samt hälso- och konsumentskyddet. Åtgärderna i detta direktiv säkerställer en hög hälso- och konsumentskyddsnivå.
(2) Textilier och läderartiklar som innehåller vissa azofärgämnen kan avge arylaminer som kan innebära risk för cancer.
(3) Fullbordandet av den inre marknaden och dess funktion påverkas av att vissa medlemsstater redan har begränsat eller planerat att begränsa användningen av azofärgade textilier och läderartiklar. Det är därför nödvändigt att tillnärma medlemsstaternas lagstiftning på detta område, och bilaga I till rådets direktiv 76/769/EEG av den 27 juli 1976 om tillnärmning av medlemsstaternas lagar och andra författningar om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar)(4) måste därför ändras.
(4) Vetenskapliga kommittén för toxicitet, ekotoxicitet och miljö har efter det att kommissionen samrått med den bekräftat att cancerrisken som orsakas av textilier och läderartiklar som färgats med vissa azofärgämnen ger anledning till oro.
(5) För att skydda människors hälsa bör användning av farliga azofärgämnen och utsläppande på marknaden av vissa artiklar som färgats med sådana färgämnen förbjudas.
(6) För textilier som framställts av återanvända fibrer bör en maximikoncentration på 70 ppm tillämpas för de aminer som är förtecknade i punkt 43 i tillägget till direktiv 76/769/EEG. Detta bör gälla under en övergångsperiod fram till den 1 januari 2005 om aminerna avges via rester från tidigare färgning av samma fibrer. Detta kommer att möjliggöra återanvändning av textilier, vilket generellt sett är gynnsamt för miljön.
(7) Tillämpningen av detta direktiv kräver harmoniserade analysmetoder. Kommissionen bör fastställa sådana metoder i enlighet med artikel 2a i direktiv 76/769/EEG. Analysmetoderna bör företrädesvis utarbetas på europeisk nivå, om så är lämpligt av Europeiska standardiseringskommittén (CEN).
(8) Mot bakgrund av nya vetenskapliga rön bör analysmetoderna ses över, inbegripet metoder för att analysera 4-aminoazobensen.
(9) Mot bakgrund av nya vetenskapliga rön bör bestämmelserna om vissa azofärger ses över, särskilt när det gäller behovet av att inbegripa andra material som inte omfattas av detta direktiv och andra aromatiska aminer. Särskild uppmärksamhet bör ägnas eventuella risker för barn.
(10) Detta direktiv påverkar inte tillämpningen av gemenskapens lagstiftning om minimikrav för arbetarskydd i rådets direktiv 89/391/EEG(5) och i särdirektiv som grundas på det direktivet, i synnerhet rådets direktiv 90/394/EEG(6) och Europaparlamentets och rådets direktiv 98/24/EG(7).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till direktiv 76/769/EEG ändras härmed i enlighet med bilagan till det här direktivet.
Artikel 2
Kommissionen skall i enlighet med förfarandet i artikel 2a i direktiv 76/769/EEG anta analysmetoder för tillämpning av punkt 43 i bilaga I till det direktivet.
De skall tillämpa dessa bestämmelser från och med 11 september 2003.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 4
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
Europaparlamentets och rådets direktiv 2002/85/EG
av den 5 november 2002
om ändring av rådets direktiv 92/6/EEG om montering och användning av hastighetsbegränsande anordningar i vissa kategorier av motorfordon inom gemenskapen
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 71 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Säkerheten vid transporter samt miljöfrågor i samband med transporter är mycket viktiga för en hållbar rörlighet.
(2) Användningen av hastighetsbegränsande anordningar för de tyngsta motorfordonskategorierna har haft en gynnsam inverkan på trafiksäkerheten. Den har också bidragit till miljöskyddet.
(3) I rådets direktiv 92/6/EEG(4) anges att kraven på montering och användning av hastighetsbegränsande anordningar senare kan utvidgas till att omfatta lättare nyttofordon, beroende på de tekniska möjligheterna och erfarenheterna i medlemsstaterna.
(4) Utvidgningen av tillämpningsområdet för direktiv 92/6/EEG till att omfatta fordon på över 3,5 ton avsedda för godstransport eller personbefordran var en av de åtgärder som rådet förordade i sin resolution av den 26 juni 2000 om ökad vägtrafiksäkerhet(5), i enlighet med kommissionens meddelande av den 20 mars 2000 om prioriteringar när det gäller vägtrafiksäkerheten inom Europeiska unionen.
(5) Tillämpningsområdet för direktiv 92/6/EEG bör utvidgas till att omfatta motorfordon i kategori M2, fordon i kategori M3 med en totalvikt på över 5 ton men högst 10 ton samt till fordon i kategori N2.
(6) Eftersom målen för den föreslagna åtgärden, nämligen att ändra gemenskapsbestämmelserna om montering och användning av hastighetsbegränsande anordningar i vissa tunga motorfordonskategorier, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför på grund av åtgärdens omfattning och verkningar bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
(7) Direktiv 92/6/EEG bör ändras i enlighet härmed.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 92/6/EEG ändras på följande sätt:
1. Artiklarna 1-5 skall ersättas med följande:
"Artikel 1
I detta direktiv avses med motorfordon sådana motordrivna fordon som tillhör någon av kategorierna M2, M3, N2 eller N3, är avsedda att användas på väg, har minst fyra hjul och är konstruerade för en högsta hastighet som överstiger 25 km/h.
Med kategori M2, M3, N2 och N3 avses de kategorier som anges i bilaga II till direktiv 70/156/EEG(6).
Artikel 2
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att de motorfordon i kategorierna M2 och M3 som avses i artikel 1 används på väg endast om de är utrustade med en hastighetsbegränsande anordning som ställts in så att fordonens hastighet inte kan överskrida 100 km/h.
Fordon i kategori M3 vars totalvikt överstiger 10 ton och som registrerades före den 1 januari 2005 får även i fortsättningen vara utrustade med anordningar där den högsta hastigheten ställts in på 100 km/h.
Artikel 3
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att motorfordon i kategorierna N2 och N3 används på väg endast om de är utrustade med en hastighetsbegränsande anordning som ställts in så att fordonens hastighet inte kan överskrida 90 km/h.
2. När det gäller den hastighetsbegränsande anordningen i fordon som är registrerade inom medlemsstaternas territorium och som endast används för transport av farligt gods har medlemsstaterna rätt att kräva att denna är inställd så att dessa fordon inte kan överskrida en högsta hastighet som understiger 90 km/h.
Artikel 4
1. När det gäller motorfordon i kategori M3 med en totalvikt på över 10 ton och motorfordon i kategori N3, skall artiklarna 2 och 3 tillämpas på
a) fordon som registrerats den 1 januari 1994 eller senare, från och med den 1 januari 1994,
b) fordon som registrerats mellan den 1 januari 1988 och den 1 januari 1994,
i) från och med den 1 januari 1995 om det rör sig om fordon som används för såväl nationella som internationella transporter,
ii) från och med den 1 januari 1996 om det rör sig om fordon som endast används för nationella transporter.
2. När det gäller motorfordon i kategori M2, fordon i kategori M3 med en totalvikt på över 5 ton men högst 10 ton samt fordon i kategori N2, skall artiklarna 2 och 3 senast tillämpas på
a) fordon som registrerats den 1 januari 2005 eller senare, från och med den 1 januari 2005,
b) fordon som uppfyller de gränsvärden som anges i direktiv 88/77/EEG(7) och registrerats mellan den 1 oktober 2001 och den 1 januari 2005,
i) från och med den 1 januari 2006, om det rör sig om fordon som används för såväl nationella som internationella transporter,
ii) från och med den 1 januari 2007, om det rör sig om fordon som endast används för nationella transporter.
3. Varje medlemsstat får bevilja undantag från tillämpningen av artiklarna 2 och 3 under högst tre år från och med den 1 januari 2005 för fordon som tillhör kategori M2 eller som tillhör kategori N2 med en totalvikt på över 3,5 ton men högst 7,5 ton, är registrerade i det nationella fordonsregistret och inte används på en annan medlemsstats territorium.
Artikel 5
1. De hastighetsbegränsande anordningar som avses i artiklarna 2 och 3 skall uppfylla de tekniska krav som fastställs i bilagan till direktiv 92/24/EEG(8). Alla fordon som omfattas av det här direktivet och registrerats före den 1 januari 2005 får dock även i fortsättningen vara utrustade med sådana hastighetsbegränsande anordningar som uppfyller de tekniska krav som fastställts av de behöriga nationella myndigheterna.
2. Hastighetsbegränsande anordningar skall monteras av sådana verkstäder eller organ som är godkända av medlemsstaterna.".
2. Följande artikel skall läggas till:
"Artikel 6a
Kommissionen skall i samband med åtgärdsprogrammet om trafiksäkerhet för perioden 2002-2010 utvärdera återverkningarna på trafiksäkerheten och vägtrafiken av att de hastighetsbegränsande anordningar som föreskrivs i detta direktiv används i fordon i kategori M2 och fordon i kategori N2 med en totalvikt av högst 7,5 ton.
Kommissionen skall vid behov lägga fram lämpliga förslag.".
Artikel 2
Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 2005. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 3
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
Europaparlamentets och rådets direktiv 2002/87/EG
av den 16 december 2002
om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat och om ändring av rådets direktiv 73/239/EEG, 79/267/EEG, 92/49/EEG, 92/96/EEG, 93/6/EEG och 93/22/EEG samt Europaparlamentets och rådets direktiv 98/78/EG och 2000/12/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 47.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
med beaktande av Europeiska centralbankens yttrande(3),
i enlighet med förfarandet i artikel 251 i fördraget(4), och
av följande skäl:
(1) Den nuvarande gemenskapslagstiftningen innehåller ett omfattande regelverk om tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag på enskild nivå samt över kreditinstitut, försäkringsföretag och värdepappersföretag som utgör en del av en bank- eller investeringsgrupp respektive en försäkringsgrupp, det vill säga grupper med en homogen finansiell verksamhet.
(2) Den senaste utvecklingen på finansmarknaderna har lett till skapandet av finansiella grupper som tillhandahåller tjänster och produkter inom olika sektorer av finansmarknaderna - så kallade finansiella konglomerat. Hittills har det inte förekommit någon form av tillsyn på gruppnivå över kreditinstitut, försäkringsföretag och värdepappersföretag som ingår i ett sådant konglomerat, särskilt vad gäller solvensställning och riskkoncentration på konglomeratnivå, transaktioner inom det finansiella konglomeratet, processer för intern riskhantering på konglomeratnivå och ledningens lämplighet. Några av dessa konglomerat är bland de största finansiella grupper som verkar på finansmarknaderna, och de tillhandahåller tjänster i en global omfattning. Om sådana konglomerat, och särskilt kreditinstitut, försäkringsföretag och värdepappersföretag som ingår i ett sådana konglomerat, skulle stöta på finansiella problem kan de allvarligt destabilisera det finansiella systemet och påverka enskilda insättare, försäkringstagare och investerare.
(3) I kommissionens handlingsplan för finansiella tjänster utpekas en rad åtgärder som krävs för att fullborda den inre marknaden för finansiella tjänster, och det aviseras att det skall utarbetas lagstiftning om extra tillsyn för finansiella konglomerat i syfte att eliminera kryphål i den nuvarande särlagstiftningen och hantera ytterligare stabilitetsrisker för att på så sätt säkra sunda arrangemang för tillsyn över finansiella grupper med sektorsöverskridande finansiell verksamhet. Ett så ambitiöst mål kan bara uppnås stegvis. Införandet av extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat utgör ett sådant steg.
(4) Även inom andra internationella forum har behovet av att utveckla lämpliga tillsynsformer för finansiella konglomerat slagits fast.
(5) För att den extra tillsynen över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat skall bli effektiv bör den tillämpas på alla sådana konglomerat, vars sektorsöverskridande finansiella verksamhet är betydande, vilket är fallet när vissa trösklar har uppnåtts oavsett hur de är strukturerade. Denna extra tillsyn bör täcka all finansiell verksamhet som anges i den finansiella särlagstiftningen och alla enheter som huvudsakligen ägnar sig åt sådan verksamhet bör omfattas av den extra tillsynen, inklusive kapitalförvaltningsbolagen.
(6) Beslut att inte låta en viss enhet omfattas av räckvidden för den extra tillsynen bör fattas med beaktande bl.a. av om en sådan enhet omfattas av tillsynen på gruppnivå enligt särreglerna.
(7) De behöriga myndigheterna bör kunna bedöma den finansiella ställningen på gruppnivå för kreditinstitut, försäkringsföretag och värdepappersföretag som ingår i ett finansiellt konglomerat, särskilt vad gäller solvens (inbegripet att eliminera dubbelt utnyttjande av poster i kapitalbasen), riskkoncentration och transaktioner inom det finansiella konglomeratet.
(8) Finansiella konglomerat leds ofta utifrån affärsområden som inte helt motsvarar konglomeratets juridiska strukturer. För att beakta denna tendens bör kraven på ledningen utvidgas ytterligare, särskilt när det gäller ledningen av blandade finansiella holdingföretag.
(9) Samtliga finansiella konglomerat som omfattas av den extra tillsynen bör ha en samordnare som utses bland berörda behöriga myndigheter.
(10) Samordnarens uppgifter bör inte påverka de behöriga myndigheternas uppgifter och ansvar enligt särreglerna.
(11) De berörda behöriga myndigheterna och särskilt samordnaren bör ha de erforderliga medlen för att från enheterna i ett finansiellt konglomerat eller från andra behöriga myndigheter kunna erhålla de upplysningar som krävs för att utöva sin extra tillsyn.
(12) Det finns ett trängande behov av ett ökat samarbete mellan de myndigheter som ansvarar för tillsynen över kreditinstitut, försäkringsföretag och värdepappersföretag, inbegripet att utveckla särskilda arrangemang för samarbete mellan de myndigheter som är delaktiga i tillsynen över enheter som ingår i samma finansiella konglomerat.
(13) Kreditinstitut, försäkringsföretag och värdepappersföretag som har sitt huvudkontor i gemenskapen kan ingå i ett finansiellt konglomerat vars ledande enhet ligger utanför gemenskapen. Dessa reglerade enheter bör också vara föremål för sådana likvärdiga och lämpliga ordningar för extra tillsyn som medför att liknande mål och resultat som de som anges i bestämmelserna i detta direktiv uppnås. Insyn i bestämmelserna och informationsutbyte med myndigheter i tredje land om alla viktiga omständigheter är här av stor vikt.
(14) Det kan antas att det finns en likvärdig och lämplig ordning för extra tillsyn endast om tillsynsmyndigheterna i tredje land har samtyckt till att samarbeta med de berörda behöriga myndigheterna om metoderna och målen för att utöva extra tillsyn över reglerade enheter i ett finansiellt konglomerat.
(15) Av detta direktiv följer inte att de behöriga myndigheterna till Kommittén för finansiella konglomerat skall lämna ut information som är belagd med sekretess enligt detta direktiv eller andra sektorsdirektiv.
(16) Eftersom målet för den föreslagna åtgärden, nämligen att fastställa regler för extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och därför, på grund av den planerade åtgärdens omfattning eller verkningar, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå detta mål. Eftersom det i direktivet anges minimistandarder, kan medlemsstaterna införa strängare regler.
(17) I detta direktiv iakttas de grundläggande rättigheter och principer som erkänns särskilt i Europeiska unionens stadga om grundläggande rättigheter.
(18) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(5).
(19) Teknisk vägledning och genomförandeåtgärder för de bestämmelser som fastställs i detta direktiv kan ibland vara nödvändiga med hänsyn till ny utveckling på finansmarknaderna. Kommissionen bör följaktligen bemyndigas att anta genomförandeåtgärder, förutsatt att dessa inte ändrar det väsentliga innehållet i detta direktiv.
(20) De befintliga särreglerna för kreditinstitut, försäkringsföretag och värdepappersföretag bör kompletteras upp till en miniminivå, särskilt för att undvika tillsynsarbitrage mellan särreglerna och reglerna för finansiella konglomerat. Rådets första direktiv 73/239/EEG av den 24 juli 1973 om samordning av lagar och andra författningar angående rätten att etablera och driva verksamhet med annan direkt försäkring än livförsäkring(6), rådets första direktiv 79/267/EEG av den 5 mars 1979 om samordning av lagar och andra författningar om rätten att starta och driva direkt livförsäkringsrörelse(7), rådets direktiv 92/49/EEG av den 18 juni 1992 om samordning av lagar och andra författningar som avser annan direkt försäkring än livförsäkring (tredje direktivet om annan direkt försäkring än livförsäkring)(8), rådets direktiv 92/96/EEG av den 10 november 1992 om samordning av lagar och andra författningar som avser direkt livförsäkring (tredje livförsäkringsdirektivet)(9), rådets direktiv 93/6/EEG av den 15 mars 1993 om kapitalkrav för värdepappersföretag och kreditinstitut(10) och rådets direktiv 93/22/EEG av den 10 maj 1993 om investeringstjänster inom värdepappersområdet(11) samt Europaparlamentets och rådets direktiv 98/78/EG av den 27 oktober 1998 om extra tillsyn över försäkringsföretag som ingår i en försäkringsgrupp(12) och Europaparlamentets och rådets direktiv 2000/12/EG av den 20 mars 2000 om rätten att starta och driva verksamhet i kreditinstitut(13) bör därför ändras på motsvarande sätt. Målet om ytterligare harmonisering kan dock bara uppnås stegvis och måste baseras på en grundlig analys.
(21) För att man skall kunna bedöma behovet av ytterligare harmonisering av behandlingen av kapitalförvaltningsbolag som omfattas av särregler och förbereda denna harmonisering bör kommissionen rapportera om medlemsstaternas praxis på detta område.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
MÅL OCH DEFINITIONER
Artikel 1
Mål
I detta direktiv fastställs regler för extra tillsyn över reglerade enheter som har erhållit auktorisation enligt artikel 6 i direktiv 73/239/EEG, artikel 6 i direktiv 79/267/EEG, artikel 3.1 i direktiv 93/22/EEG eller artikel 4 i direktiv 2000/12/EG och som ingår i ett finansiellt konglomerat. Genom direktivet ändras också berörda särregler för enheter som regleras av ovannämnda direktiv.
Artikel 2
Definitioner
I detta direktiv används följande beteckningar med de betydelser som här anges:
1. kreditinstitut: ett kreditinstitut i den mening som avses i artikel 1.1 andra stycket i direktiv 2000/12/EG.
2. försäkringsföretag: ett försäkringsföretag i den mening som avses i artikel 6 i direktiv 73/239/EEG, artikel 6 i direktiv 79/267/EEG eller artikel 1 b i direktiv 98/78/EG.
3. värdepappersföretag: ett värdepappersföretag i den mening som avses i artikel 1.2 i direktiv 93/22/EEG, inbegripet företag som avses i artikel 2.4 i direktiv 93/6/EEG.
4. reglerad enhet: ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag.
5. kapitalförvaltningsbolag: ett förvaltningsbolag i den mening som avses i artikel 1a.2 i rådets direktiv 85/611/EEG av den 20 december 1985 om samordning av lagar och andra författningar som avser företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag)(14), samt ett företag vars säte är beläget utanför gemenskapen, vilket, om det hade sitt säte i gemenskapen, skulle behöva auktorisation i enlighet med artikel 5.1 i det direktivet.
6. återförsäkringsföretag: ett återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG.
7. särregler: gemenskapslagstiftning som rör tillsynen över reglerade enheter, särskilt den som fastställs i direktiv 73/239/EEG, 79/267/EEG, 98/78/EG, 93/6/EEG, 93/22/EEG och 2000/12/EG.
8. finansiell sektor: en sektor som består av en eller flera av följande enheter:
a) Ett kreditinstitut, ett finansiellt institut eller ett företag som tillhandahåller tjänster anknutna till bankverksamhet enligt artikel 1.5 och 1.23 i direktiv 2000/12/EG (banksektorn).
b) Ett försäkringsföretag, ett återförsäkringsföretag eller ett försäkringsholdingbolag enligt artikel 1 led i i direktiv 98/78/EG (försäkringssektorn).
c) Ett värdepappersföretag eller ett finansiellt institut enligt artikel 2.7 i direktiv 93/6/EEG (sektorn för investeringstjänster).
d) Ett blandat finansiellt holdingföretag.
9. moderföretag:ett moderföretag i den mening som avses i artikel 1 i rådets sjunde direktiv 83/349/EEG av den 13 juni 1983 om sammanställd redovisning(15) och varje företag som enligt de behöriga myndigheterna i praktiken utövar ett bestämmande inflytande över ett annat företag.
10. dotterföretag: ett dotterföretag i den mening som avses i artikel 1 i direktiv 83/349/EEG och varje företag över vilket ett moderföretag enligt de behöriga myndigheterna i praktiken utövar ett bestämmande inflytande. Alla dotterföretag till dotterföretag skall också betraktas som dotterföretag till det moderföretag som är överordnat dessa företag.
11. ägarintresse: ett ägarintresse i den mening som avses i artikel 17 första meningen i rådets fjärde direktiv 78/660/EEG av den 25 juli 1978 om årsbokslut i vissa typer av bolag(16) eller direkt eller indirekt ägande av 20 % eller mer av rösterna eller kapitalet i ett företag.
12. grupp: en grupp av företag som består av ett moderföretag, dess dotterföretag och enheter i vilka moderföretaget och dess dotterföretag har ägarintressen samt företag som är knutna till varandra genom ett sådant förhållande som avses i artikel 12.1 i direktiv 83/349/EEG.
13. nära förbindelser: en situation där två eller flera fysiska eller juridiska personer är förenade genom
a) ägarintresse, innebärande ett innehav, direkt eller genom kontroll av 20 % eller mer av rösterna eller kapitalet i ett företag, eller
b) kontroll, innebärande förbindelse mellan ett moderföretag och ett dotterföretag i alla de fall som omfattas av artikel 1.1 och 1.2 i direktiv 83/349/EEG, eller en likartad förbindelse mellan någon fysisk eller juridisk person och ett företag. Varje dotterföretag till ett dotterföretag skall också anses som dotterföretag till moderföretaget vilket står över dessa företag.
Som nära förbindelse skall även anses en situation där två eller flera fysiska eller juridiska personer kontrolleras genom en varaktig förbindelse till en och samma person.
14. finansiellt konglomerat: en grupp som uppfyller följande villkor, om inte annat följer av artikel 3:
a) En reglerad enhet i den mening som avses i artikel 1 finns i toppen av gruppen eller minst ett av dotterföretagen i gruppen är en reglerad enhet i den mening som avses i artikel 1.
b) Om en reglerad enhet i den mening som avses i artikel 1 finns i toppen av gruppen, är den antingen ett moderföretag till en enhet i den finansiella sektorn, en enhet med ägarintresse i en enhet i den finansiella sektorn eller en enhet som har ett sådant samband med en enhet i den finansiella sektorn som avses i artikel 12.1 i direktiv 83/349/EEG.
c) Om ingen reglerad enhet i den mening som avses i artikel 1 finns i toppen av gruppen, bedrivs gruppens verksamhet huvudsakligen inom den finansiella sektorn i den mening som avses i artikel 3.1.
d) Minst en av gruppens enheter ingår i försäkringssektorn och minst en i bank- eller värdepapperssektorn.
e) Den konsoliderade och/eller aggregerade verksamheten i gruppens enheter inom försäkringssektorn och den konsoliderade och/eller aggregerade verksamheten i gruppens enheter inom bank- och värdepapperssektorn är betydande enligt artikel 3.2 eller 3.3.
Varje undergrupp till en grupp enligt punkt 12 som uppfyller kriterierna i denna punkt skall anses vara ett finansiellt konglomerat.
15. blandat finansiellt holdingföretag: ett moderföretag som inte utgör en reglerad enhet men som tillsammans med sina dotterföretag, varav minst ett är en reglerad enhet med huvudkontor inom gemenskapen, och andra enheter utgör ett finansiellt konglomerat.
16. behöriga myndigheter: de nationella myndigheter i medlemsstaterna som enligt lag eller annan författning har behörighet att utöva tillsyn över kreditinstitut, försäkringsföretag och/eller värdepappersföretag såväl enskilt som på gruppnivå.
17. relevanta behöriga myndigheter:
a) de behöriga myndigheter i medlemsstaterna som har ansvar för den sektoriella tillsynen på gruppnivå över de reglerade enheterna i ett finansiellt konglomerat,
b) samordnaren som utsetts i enlighet med artikel 10, om annan än de myndigheter som anges under a,
c) andra berörda behöriga myndigheter, om de myndigheter som anges under a och b anser detta vara relevant. Vid en sådan bedömning skall särskilt beaktas den marknadsandel de reglerade enheterna i konglomeratet har i andra medlemsstater, i synnerhet om den överstiger 5 %, och den betydelse varje reglerad enhet som är etablerad i en annan medlemsstat har inom konglomeratet.
18. transaktioner inom det finansiella konglomeratet: alla transaktioner genom vilka reglerade enheter inom ett finansiellt konglomerat direkt eller indirekt anlitar andra företag inom samma grupp eller en fysisk eller juridisk person som har "nära förbindelser" med företagen i den gruppen, för att uppfylla en skyldighet, oavsett om den är avtalsenlig eller ej och om den sker mot betalning eller ej.
19. riskkoncentration: alla exponeringar med förlustpotential som bärs av enheter inom ett finansiellt konglomerat, vilka är tillräckligt stora för att hota dessa reglerade enheters solvens eller deras finansiella ställning i allmänhet; sådana exponeringar kan orsakas av motpartsrisk/kreditrisk, investeringsrisk, försäkringsrisk, marknadsrisk eller andra risker, eller en kombination av eller samverkan mellan dessa risker.
Artikel 3
Tröskelvärden för identifiering av ett finansiellt konglomerat
1. För att en grupp skall bedömas bedriva verksamhet huvudsakligen inom den finansiella sektorn i den mening som avses i artikel 2.14 c, skall balansomslutningen inom gruppens reglerade och icke reglerade enheter inom den finansiella sektorn utgöra mer än 40 % av hela gruppens balansomslutning.
2. För att verksamheten inom olika finansiella sektorer skall bedömas som betydande i den mening som avses i artikel 2.14 e, skall för varje finansiell sektor genomsnittet av kvoten mellan denna finansiella sektors balansomslutning och den totala balansomslutningen för gruppens enheter inom finansiella sektorer och kvoten mellan solvenskraven för denna finansiella sektor och de totala solvenskraven för gruppens enheter inom finansiella sektorer överstiga 10 %.
I detta direktiv är den minsta finansiella sektorn i ett finansiellt konglomerat den sektor som har det lägsta genomsnittet och den mest betydande finansiella sektorn i ett finansiellt konglomerat den sektor som har det högsta genomsnittet. Vid beräkningen av genomsnittet för den minsta finansiella sektorn och den mest betydande finansiella sektorn skall banksektorn och värdepapperssektorn beaktas tillsammans.
3. Sektorsövergripande verksamhet skall också bedömas som betydande i den mening som avses i artikel 2.14 e, om balansomslutningen för den minsta finansiella sektorn i gruppen överstiger 6 miljarder euro. Om gruppen inte uppnår det tröskelvärde som anges i punkt 2, får de relevanta behöriga myndigheterna i samförstånd besluta sig för att inte betrakta gruppen som ett finansiellt konglomerat eller att inte tillämpa bestämmelserna i artiklarna 7, 8 eller 9, om de anser att det inte är nödvändigt eller att det vore olämpligt eller vilseledande att låta gruppen omfattas av detta direktivs räckvidd eller att tillämpa sådana bestämmelser med hänsyn till de mål som skall uppnås genom extra tillsyn, till exempel med beaktande av följande:
a) Den relativa storleken på dess minsta finansiella sektor överstiger inte 5 %, mätt antingen i termer av det genomsnitt som anges i punkt 2 eller i termer av balansomslutningen eller solvenskraven för en sådan finansiell sektor.
b) Marknadsandelen överstiger inte 5 % i någon medlemsstat, mätt i termer av balansomslutningen för bank- och värdepapperssektorerna och i termer av tecknade bruttopremier inom försäkringssektorn.
Beslut som fattas i överensstämmelse med denna punkt skall anmälas till övriga berörda behöriga myndigheter.
4. För tillämpningen av punkterna 1, 2 och 3 får de relevanta behöriga myndigheterna i samförstånd
a) undanta en enhet från beräkningen av procentsatserna i de fall som avses i artikel 6.5,
b) beakta att de trösklar som anges i punkterna 1 och 2 har iakttagits under tre år i följd, så att plötsliga byten av det tillämpliga regelverket kan undvikas, och bortse ifrån att så har skett, om väsentliga förändringar i gruppens struktur uppstår.
När ett finansiellt konglomerat har identifierats enligt punkterna 1, 2 och 3 skall de beslut som avses i första stycket och detta stycke fattas på grundval av ett förslag från samordnaren för detta finansiella konglomerat.
5. Vid tillämpningen av punkterna 1 och 2 får de relevanta behöriga myndigheterna, i exceptionella fall och i samförstånd, ersätta balansomslutningen som kriterium med en av följande parametrar eller båda eller lägga till en eller båda av dessa parametrar, om de anser att de är av särskild relevans för den extra tillsynen enligt detta direktiv: intäktsstruktur, poster utanför balansräkningen.
6. Om de procentsatser som avses i punkterna 1 och 2 hamnar under 40 % respektive 10 % för konglomerat som redan är föremål för extra tillsyn, skall vid tillämpningen av dessa punkter en lägre procentsats på 35 % respektive 8 % tillämpas under de tre följande åren, för att plötsliga byten av tillämpligt regelverk skall undvikas.
Vid tillämpningen av punkt 3 skall, om balansomslutningen för den minsta finansiella sektorn inom gruppen understiger 6 miljarder euro för konglomerat som redan är föremål för extra tillsyn, även ett lägre belopp om 5 miljarder euro tillämpas under de tre följande åren, för att plötsliga byten av tillämpligt regelverk skall kunna undvikas.
Under den period som avses i denna punkt får samordnaren, med medgivande från de övriga relevanta behöriga myndigheterna, besluta att de lägre procentsatser eller det lägre belopp som anges i denna punkt inte längre skall tillämpas.
7. De beräkningar som anges i denna artikel och som rör balansräkningen skall utföras på grundval av den aggregerade balansomslutningen för gruppens enheter enligt deras årsbokslut. Vid denna beräkning skall företag som är föremål för ett ägarintresse ingå till det belopp i deras balansomslutning som motsvarar den aggregerade proportionella andel som gruppen innehar. Om sammanställd redovisning emellertid finns tillgänglig, skall denna användas i stället för aggregerad redovisning.
De solvenskrav som avses i punkterna 2 och 3 skall beräknas enligt bestämmelserna i de relevanta särreglerna.
Artikel 4
Identifiering av ett finansiellt konglomerat
1. De behöriga myndigheter som har auktoriserat reglerade enheter skall på grundval av artiklarna 2, 3 och 5 identifiera varje grupp som omfattas av detta direktivs räckvidd.
För detta ändamål
- skall de behöriga myndigheter som har auktoriserat reglerade enheter i denna grupp, om så är nödvändigt, ha ett nära samarbete,
- skall en behörig myndighet som anser att en av denna myndighet auktoriserad reglerad enhet tillhör en grupp som kan vara ett finansiellt konglomerat, som inte redan har identifierats enligt detta direktiv, underrätta de andra berörda behöriga myndigheterna om sin inställning.
2. Den samordnare som utsetts enligt artikel 10 skall informera det moderföretag som finns i toppen av en grupp eller, i avsaknad av moderföretag, den reglerade enhet som har den största balansomslutningen inom den största finansiella sektorn i en grupp, om att gruppen har identifierats som ett finansiellt konglomerat och om utnämningen av samordnare. Samordnaren skall också informera de behöriga myndigheter som har auktoriserat reglerade enheter i gruppen och de behöriga myndigheterna i den medlemsstat i vilken det blandade finansiella holdingföretaget har sitt huvudkontor samt kommissionen.
KAPITEL II
EXTRA TILLSYN
AVSNITT I
RÄCKVIDD
Artikel 5
Räckvidd för den extra tillsynen över de reglerade enheter som avses i artikel 1
1. Utan att det påverkar särreglernas bestämmelser om tillsyn skall medlemsstaterna ombesörja extra tillsyn över de reglerade enheter som avses i artikel 1, i den omfattning och på det sätt som föreskrivs i detta direktiv.
2. Följande reglerade enheter skall underkastas extra tillsyn på nivån finansiella konglomerat i enlighet med artiklarna 6-17:
a) Varje reglerad enhet i toppen av ett finansiellt konglomerat.
b) Varje reglerad enhet vars moderföretag är ett blandat finansiellt holdingföretag med huvudkontor inom gemenskapen.
c) Varje reglerad enhet som har ett sådant samband med en annan enhet i den finansiella sektorn som avses i artikel 12.1 i direktiv 83/349/EEG.
Om ett finansiellt konglomerat är en undergrupp till ett annat finansiellt konglomerat som uppfyller kraven i första stycket, får medlemsstaterna tillämpa artiklarna 6-17 enbart på reglerade enheter i den senare gruppen, och alla hänvisningar i direktivet till begreppen grupp och finansiellt konglomerat skall då anses syfta på denna.
3. Varje reglerad enhet som inte är föremål för extra tillsyn enligt punkt 2 och vars moderföretag är en reglerad enhet eller ett blandat finansiellt holdingföretag med huvudkontor utanför gemenskapen skall vara föremål för extra tillsyn på nivån finansiellt konglomerat i den omfattning och på det sätt som föreskrivs i artikel 18.
4. Om personer har ägarintresse i eller kapitalförbindelser med en eller flera reglerade enheter eller utövar ett betydande inflytande över sådana enheter utan att ha ägarintresse eller kapitalförbindelser utöver de fall som avses i punkterna 2 och 3, skall de relevanta behöriga myndigheterna i samförstånd och i enlighet med den nationella lagstiftningen avgöra huruvida och i vilken omfattning extra tillsyn skall utövas över dessa reglerade enheter som om de utgjorde ett finansiellt konglomerat.
För att sådan extra tillsyn skall kunna utövas, skall minst en av enheterna vara en reglerad enhet enligt artikel 1 och de villkor som anges i artikel 2.14 d och e skall vara uppfyllda. De relevanta behöriga myndigheterna skall fatta sitt beslut med beaktande av de mål för extra tillsyn som anges i detta direktiv.
Vid tillämpning av det första stycket på "kooperativa grupper" skall de behöriga myndigheterna beakta de offentliga finansieringsåtaganden som dessa grupper har gentemot andra finansiella enheter.
5. Utan att det påverkar tillämpningen av artikel 13 skall utövandet av extra tillsyn på nivån finansiellt konglomerat inte på något sätt anses innebära att de behöriga myndigheterna är skyldiga att utöva tillsyn över blandade finansiella holdingföretag, över reglerade enheter i tredje land som tillhör ett finansiellt konglomerat eller över enskilda icke reglerade enheter i ett finansiellt konglomerat.
AVSNITT 2
FINANSIELL STÄLLNING
Artikel 6
Kapitaltäckning
1. Utan att särreglerna åsidosätts skall extra tillsyn över kapitaltäckningen i de reglerade enheterna i ett finansiellt konglomerat utövas enligt de regler som anges i punkterna 2-5, i artikel 9, i avsnitt 3 i detta kapitel och i bilaga I.
2. Medlemsstaterna skall kräva att reglerade enheter i ett finansiellt konglomerat säkerställer att det finns en tillgänglig kapitalbas på nivån finansiellt konglomerat som alltid minst motsvarar de kapitaltäckningskrav som beräknas enligt bilaga I.
Medlemsstaterna skall också kräva att reglerade enheter följer en adekvat kapitaltäckningsstrategi på nivån finansiellt konglomerat.
De krav som avses i första och andra stycket skall vara föremål för samordnarens tillsyn enligt avsnitt 3.
Samordnaren skall se till att den beräkning som avses i första stycket utförs minst en gång per år, antingen av de reglerade enheterna eller av det blandade finansiella holdingföretaget.
Resultatet av beräkningen och relevanta uppgifter för beräkningen skall överlämnas till samordnaren av den reglerade enhet i den mening som avses i artikel 1 som finns i toppen av det finansiella konglomeratet eller, när det finansiella konglomeratet inte har en reglerad enhet i den mening som avses i artikel 1 i toppen, av det blandade finansiella holdingföretaget eller av den reglerade enhet i det finansiella konglomeratet som identifierats av samordnaren efter samråd med de övriga relevanta behöriga myndigheterna och med det finansiella konglomeratet.
3. För den beräkning av kapitaltäckningskraven som avses i punkt 2 första stycket skall följande enheter omfattas av extra tillsyn i den form och utsträckning som fastställs i bilaga I:
a) Kreditinstitut, finansiella institut eller företag som tillhandahåller tjänster anknutna till bankverksamhet i den mening som avses i artikel 1.5 och 1.23 i direktiv 2000/12/EG.
b) Försäkringsföretag, återförsäkringsföretag eller försäkringsholdingbolag i den mening som avses i artikel 1 i i direktiv 98/78/EG.
c) Värdepappersföretag eller finansiella institut i den mening som avses i artikel 2.7 i direktiv 93/6/EEG.
d) Blandade finansiella holdingföretag.
4. Vid beräkning av de extra kapitaltäckningskraven avseende ett finansiellt konglomerat genom tillämpning av metod 1 (metod baserad på sammanställd redovisning) som avses i bilaga I skall kapitalbas och solvenskrav för enheterna i gruppen beräknas genom tillämpning av de motsvarande särregler för sammanställningens form och omfattning som fastställs framför allt i artikel 54 i direktiv 2000/12/EG och i punkt 1 B i bilaga I till direktiv 98/78/EG.
Vid tillämpning av metod 2 eller 3 (Avräknings- och totalmetoden respektive Metod för kravavräkning eller avräkning av bokfört värde) vilka avses i bilaga I skall hänsyn tas till den proportionella andel som moderföretaget eller företaget med ägarintresse innehar i en annan enhet i gruppen. Med "proportionell andel" avses den del av det tecknade kapitalet som direkt eller indirekt innehas av detta företag.
5. Samordnaren kan besluta att inte inbegripa en viss enhet vid beräkningen av den extra kapitaltäckningskraven i följande fall:
a) Om enheten finns i ett tredje land där det finns rättsliga hinder för att överföra erforderliga upplysningar, utan att detta påverkar tillämpningen av särreglernas bestämmelser om de behöriga myndigheternas skyldighet att vägra auktorisation när de är förhindrade att effektivt utöva sin tillsyn.
b) Om enheten är av försumbar betydelse i förhållande till målen för den extra tillsynen över reglerade enheter i ett finansiellt konglomerat.
c) Om det skulle vara olämpligt eller missvisande att inbegripa enheten med hänsyn till målen för den extra tillsynen.
Om flera enheter utesluts till följd av b i första stycket, måste de dock inkluderas om de tillsammans inte är av försumbar betydelse.
I det fall som nämns i c i första stycket skall samordnaren, utom i brådskande fall, samråda med de andra relevanta behöriga myndigheterna innan beslut fattas.
Om samordnaren inte inkluderar en reglerad enhet i tillämpningsområdet med stöd av ett av de fall som anges i b och c i första stycket, får de behöriga myndigheterna i den medlemsstat där denna enhet är belägen begära att den enhet som finns i toppen av det finansiella konglomeratet lämnar upplysningar som underlättar tillsynen över den reglerade enheten.
Artikel 7
Riskkoncentration
1. Utan att särreglerna åsidosätts skall extra tillsyn över riskkoncentrationen i de reglerade enheterna i ett finansiellt konglomerat utövas enligt reglerna i artikel 9.2-9.4 i avsnitt 3 i detta kapitel och i bilaga II.
2. Medlemsstaterna skall kräva att reglerade enheter eller blandade finansiella holdingföretag regelbundet och minst en gång per år till samordnaren rapporterar varje betydande riskkoncentration på nivån finansiellt konglomerat enligt reglerna i denna artikel och i bilaga II. Den nödvändiga informationen skall överlämnas till samordnaren av den reglerade enhet i den mening som avses i artikel 1 som finns i toppen av det finansiella konglomeratet eller, när det finansiella konglomeratet inte leds av en reglerad enhet i den mening som avses i artikel 1, av det blandade finansiella holdingföretaget eller av den reglerade enhet i det finansiella konglomeratet som identifierats av samordnaren efter samråd med de övriga relevanta behöriga myndigheterna och med det finansiella konglomeratet.
Samordnaren skall övervaka dessa riskkoncentrationer i enlighet med avsnitt 3.
3. Till dess att gemenskapens lagstiftning har samordnats ytterligare får medlemsstaterna fastställa kvantitativa gränser eller tillåta sina behöriga myndigheter att fastställa kvantitativa gränser eller vidta andra tillsynsåtgärder som skulle kunna uppfylla målen för extra tillsyn när det gäller riskkoncentration på nivån finansiellt konglomerat.
4. När ett finansiellt konglomerat leds av ett blandat finansiellt holdingföretag, skall eventuella särregler om riskkoncentration i den största finansiella sektorn i det finansiella konglomeratet gälla för hela den sektorn, inklusive det blandade finansiella holdingföretaget.
Artikel 8
Transaktioner inom det finansiella konglomeratet
1. Utan att särreglerna åsidosätts skall extra tillsyn över reglerade enheters transaktioner inom det finansiella konglomeratet, utövas enligt reglerna i artikel 9.2-9.4 i avsnitt 3 i detta kapitel och bilaga II.
2. Medlemsstaterna skall kräva att reglerade enheter eller blandade finansiella holdingföretag regelbundet och minst en gång per år till samordnaren rapporterar samtliga transaktioner inom det finansiella konglomeratet enligt reglerna i denna artikel och i bilaga II. I den mån de tröskelvärden som anges i sista meningen i första stycket i bilaga II inte har fastställts, skall en transaktion inom det finansiella konglomeratet åtminstone anses som betydande, om beloppet överstiger 5 % av det totala belopp som kapitaltäckningskraven uppgår till på nivån finansiellt konglomerat.
Den nödvändiga informationen skall överlämnas till samordnaren av den reglerade enhet i den mening som avses i artikel 1 som finns i toppen av det finansiella konglomeratet eller, när det finansiella konglomeratet inte leds av en reglerad enhet i den mening som avses i artikel 1, av det blandade finansiella holdingföretaget eller av den reglerade enhet i det finansiella konglomeratet som identifierats av samordnaren efter samråd med de övriga relevanta behöriga myndigheterna och med det finansiella konglomeratet.
Samordnaren skall övervaka dessa transaktioner inom det finansiella konglomeratet.
3. Till dess att gemenskapens lagstiftning har samordnats ytterligare får medlemsstaterna fastställa kvantitativa gränser och kvalitativa krav eller tillåta sina behöriga myndigheter att fastställa kvantitativa gränser och kvalitativa krav eller vidta andra tillsynsåtgärder som skulle kunna uppfylla målen för extra tillsyn när det gäller transaktioner inom det finansiella konglomeratet av reglerade enheter i ett finansiellt konglomerat.
4. När ett finansiellt konglomerat leds av ett blandat finansiellt holdingföretag, skall särregler om transaktioner inom det finansiella konglomeratet i den största finansiella sektorn i det finansiella konglomeratet tillämpas för hela den sektorn, inklusive det blandade finansiella holdingföretaget.
Artikel 9
Rutiner för intern kontroll och metoder för riskhantering
1. Medlemsstaterna skall kräva att det hos reglerade enheter på nivån finansiellt konglomerat finns erforderliga metoder för riskhantering och rutiner för intern kontroll, inbegripet sunda rapporterings- och redovisningsförfaranden.
2. Metoderna för riskhantering skall inbegripa följande:
a) Ett sunt styre och en sund förvaltning, varvid lämpliga ledande organ på nivån finansiellt konglomerat skall godkänna och regelbundet övervaka strategier och inriktningar med beaktande av alla risker de tar.
b) En adekvat kapitaltäckningsstrategi för att kunna förutse den inverkan som deras affärsstrategi har på riskprofilen och kapitalkraven, så som de fastställts i enlighet med artikel 6 och bilaga I.
c) Lämpliga förfaranden för att säkerställa att systemen för övervakning av risker är väl integrerade i organisationen och att alla åtgärder har vidtagits för att se till att de system som genomförts i alla de företag som omfattas av extra tillsyn är samstämmiga, så att riskerna kan mätas, övervakas och kontrolleras på nivån finansiellt konglomerat.
3. Rutinerna för intern kontroll skall innehålla följande:
a) Adekvata mekanismer för kapitaltäckning för att identifiera och mäta samtliga materiella risker och på ett lämpligt sätt ställa kapitalbasen i relation till riskerna.
b) Sunda rapporterings- och redovisningsförfaranden, för att identifiera, mäta, övervaka och kontrollera transaktionerna inom det finansiella konglomeratet och riskkoncentrationen.
4. Medlemsstaterna skall se till att det i alla företag som omfattas av extra tillsyn enligt artikel 5 finns erforderliga rutiner för intern kontroll för att ta fram de uppgifter och upplysningar som kan vara av betydelse för den extra tillsynen.
5. De metoder och mekanismer som avses i punkterna 1-4 skall övervakas av samordnaren.
AVSNITT 3
ÅTGÄRDER FÖR ATT UNDERLÄTTA EXTRA TILLSYN
Artikel 10
Behörig myndighet ansvarig för utövandet av extra tillsyn (samordnaren)
1. För att säkerställa korrekt extra tillsyn över de reglerade enheterna i ett finansiellt konglomerat skall en enda samordnare med ansvar för samordning och utövande av den extra tillsynen utses bland de berörda medlemsstaternas behöriga myndigheter, inbegripet dem som finns i den medlemsstat i vilken det blandade finansiella holdingföretaget har sitt huvudkontor.
2. Utnämningen skall grunda sig på följande kriterier:
a) Om ett finansiellt konglomerat leds av en reglerad enhet, skall samordningen utövas av den behöriga myndighet som har auktoriserat denna reglerade enhet enligt gällande särregler.
b) Om ett finansiellt konglomerat inte leds av en reglerad enhet, skall den behöriga myndighet som identifieras enligt följande principer fungera som samordnare:
i) Om moderföretaget till en reglerad enhet är ett blandat finansiellt holdingföretag, skall samordningen utövas av den behöriga myndighet som har auktoriserat denna reglerade enhet enligt gällande särregler.
ii) Om två eller flera reglerade enheter med huvudkontor inom gemenskapen har samma blandade finansiella holdingföretag som moderföretag och en av dessa enheter har auktoriserats i den medlemsstat där det blandade finansiella holdingföretaget har sitt huvudkontor, skall samordningen utövas av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som auktoriserats i denna medlemsstat.
Om två eller flera reglerade enheter som verkar inom olika finansiella sektorer har auktoriserats i den medlemsstat där det blandade finansiella holdingföretaget har sitt huvudkontor, skall samordningen utövas av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som verkar inom den största finansiella sektorn.
Om det finansiella konglomeratet leds av två eller flera blandade finansiella holdingföretag vilka har huvudkontor i olika medlemsstater och det finns en reglerad enhet i var och en av dessa medlemsstater, skall samordningen utövas av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som har den största balansomslutningen, om dessa enheter verkar inom samma finansiella sektor, eller av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som verkar inom den största finansiella sektorn.
iii) Om två eller flera reglerade enheter med huvudkontor inom gemenskapen har samma blandade finansiella holdingföretag som moderföretag och ingen av dessa enheter har auktoriserats i den medlemsstat där det blandade finansiella holdingföretaget har sitt huvudkontor, skall samordningen utövas av den behöriga myndighet som har auktoriserat den reglerade enhet som har den största balansomslutningen inom den största finansiella sektorn.
iv) Om det finansiella konglomeratet utgör en grupp utan något moderföretag i toppen, eller i övriga fall, skall samordningen utövas av den behöriga myndighet som har auktoriserat den reglerade enhet som har den största balansomslutningen inom den största finansiella sektorn.
3. I särskilda fall får de relevanta behöriga myndigheterna i samförstånd bevilja undantag från de kriterier som anges i punkt 2, om det skulle vara olämpligt att tillämpa dessa kriterier, med beaktande av konglomeratets struktur och den relativa betydelsen av dess verksamhet i olika länder, och utse en annan behörig myndighet till samordnare. I dessa fall skall de behöriga myndigheterna innan de fattar sitt beslut ge konglomeratet möjlighet att yttra sig om detta beslut.
Artikel 11
Samordnarens uppgifter
1. De uppgifter som samordnaren skall utföra inom ramen för den extra tillsynen skall omfatta följande:
a) Samordning av insamling och spridning av relevanta eller väsentliga uppgifter, såväl löpande som i krissituationer, inbegripet spridning av uppgifter som är av betydelse för en behörig myndighets tillsynsuppgifter enligt särreglerna.
b) Övervakning av och bedömning av ett finansiellt konglomerats finansiella ställning.
c) Bedömning av huruvida reglerna om kapitaltäckning, riskkoncentration och transaktioner inom det finansiella konglomeratet enligt artiklarna 6, 7 och 8 följs.
d) Bedömning av det finansiella konglomeratets struktur, organisation och system för intern kontroll enligt artikel 9.
e) Planering och samordning av tillsynen, såväl löpande som i krissituationer, i samarbete med de berörda behöriga myndigheterna.
f) Andra uppgifter, åtgärder och beslut som har tilldelats samordnaren genom detta direktiv eller som följer av detta direktivs tillämpning.
För att den extra tillsynen skall kunna underlättas och få en bred rättslig grund, skall samordnaren, de andra relevanta behöriga myndigheterna och vid behov andra berörda behöriga myndigheter införa samordningsåtgärder. Genom dessa kan samordnaren anförtros ytterligare uppgifter och förfaranden specificeras för de relevanta behöriga myndigheternas beslutsprocesser enligt artiklarna 3 och 4, artikel 5.4, artikel 6, artikel 12.2 samt artiklarna 16 och 18, samt för samarbetet med andra behöriga myndigheter.
2. Samordnaren bör, när den behöver uppgifter som redan överlämnats till en annan behörig myndighet i enlighet med särreglerna, vända sig till denna myndighet närhelst detta är möjligt i syfte att undvika dubblering av rapporteringen till de olika myndigheter som utövar tillsyn.
3. Utan att det påverkar möjligheten att delegera specifika tillsynsbefogenheter och specifikt tillsynsansvar enligt gemenskapslagstiftningen, skall förekomsten av en samordnare som anförtrotts specifika uppgifter i samband med den extra tillsynen över reglerade enheter i ett finansiellt konglomerat inte påverka de behöriga myndigheternas uppgifter och ansvar enligt särreglerna.
Artikel 12
Samarbete och utbyte av uppgifter mellan behöriga myndigheter
1. De behöriga myndigheter som ansvarar för tillsynen över reglerade enheter i ett finansiellt konglomerat och den behöriga myndighet som utses till samordnare för detta skall ha ett nära samarbete med varandra. Utan att det påverkar dessa myndigheters respektive ansvar enligt särreglerna skall de, oavsett om de är inrättade i samma medlemsstat, till varandra överlämna alla uppgifter som är väsentliga eller relevanta för de övriga behöriga myndigheternas utövande av tillsynsuppgifter enligt särreglerna och detta direktiv. Härvid skall de behöriga myndigheterna och samordnaren på begäran överlämna alla relevanta uppgifter och på eget initiativ överlämna alla väsentliga uppgifter.
Detta samarbete skall åtminstone omfatta insamling och utbyte av uppgifter avseende följande punkter:
a) Identifiering av hur alla större enheter som tillhör det finansiella konglomeratet är grupperade och av de behöriga myndigheter som ansvarar för tillsynen över de reglerade enheterna i gruppen.
b) Det finansiella konglomeratets strategier.
c) Det finansiella konglomeratets finansiella ställning, särskilt när det gäller kapitaltäckning, transaktioner inom det finansiella konglomeratet, riskkoncentration och lönsamhet.
d) Det finansiella konglomeratets största aktieägare och ledning.
e) Organisation, riskhantering och system för intern kontroll på det finansiella konglomeratets nivå.
f) Förfaranden för insamling av uppgifter från enheterna i ett finansiellt konglomerat samt kontroll av de uppgifterna.
g) Negativ utveckling i reglerade enheter eller i andra enheter i det finansiella konglomeratet som skulle kunna påverka de reglerade enheterna allvarligt.
h) Större sanktioner och exceptionella åtgärder som de behöriga myndigheterna vidtar i enlighet med särreglerna eller detta direktiv.
När det är nödvändigt för utförandet av deras respektive uppgifter, kan de behöriga myndigheterna också utbyta uppgifter om reglerade enheter i ett finansiellt konglomerat med följande myndigheter i enlighet med bestämmelserna i särreglerna: centralbanker, Europeiska centralbankssystemet och Europeiska centralbanken.
2. Utan att det påverkar dessa myndigheters respektive ansvar enligt särreglerna skall de berörda behöriga myndigheterna innan de fattar beslut samråda med varandra i följande fall, om deras beslut är av betydelse för andra behöriga myndigheters tillsynsuppgifter:
a) Sådana förändringar av aktieägar-, organisations- eller ledningsstrukturen i reglerade enheter i ett finansiellt konglomerat som kräver de behöriga myndigheternas godkännande eller auktorisation.
b) Större sanktioner eller exceptionella åtgärder som de behöriga myndigheterna vidtar.
En behörig myndighet får besluta att inte samråda i brådskande situationer eller när ett sådant samråd kan äventyra effektiviteten i besluten. Den behöriga myndigheten skall i detta fall utan dröjsmål informera de andra behöriga myndigheterna.
3. När de behöriga myndigheterna i den medlemsstat där ett moderföretag har sitt huvudkontor inte själva utövar den extra tillsynen enligt artikel 10, kan samordnaren begära att de av moderföretaget inhämtar alla uppgifter som kan vara relevanta för utövandet av samordningsuppgifterna enligt artikel 11 samt att de överlämnar dessa uppgifter till samordnaren.
Om de uppgifter som avses i artikel 14.2 redan har lämnats till en behörig myndighet enligt särreglerna, kan de behöriga myndigheter som ansvarar för att utöva extra tillsyn vända sig till den förstnämnda myndigheten för att erhålla dessa uppgifter.
4. Medlemsstaterna skall godkänna att deras behöriga myndigheter utbyter de uppgifter som avses i punkterna 1, 2 och 3 med varandra och med andra myndigheter. Insamling eller innehav av uppgifter om en enhet inom ett finansiellt konglomerat vilken inte är en reglerad enhet skall inte på något sätt anses innebära att de behöriga myndigheterna är skyldiga att utöva någon tillsynsfunktion i förhållande till den enskilda enheten.
Uppgifter som erhålls inom ramen för den extra tillsynen och särskilt varje utbyte av uppgifter mellan behöriga myndigheter eller mellan behöriga myndigheter och andra myndigheter enligt detta direktiv omfattas av särreglernas bestämmelser om tystnadsplikt och överlämnande av förtrolig information.
Artikel 13
Ledningsorgan för blandade finansiella holdingföretag
Medlemsstaterna skall kräva att de personer som faktiskt leder affärsverksamheten i ett blandat finansiellt holdingföretag har ett tillräckligt gott anseende och tillräcklig erfarenhet för att kunna fullgöra sina åligganden.
Artikel 14
Tillgång till uppgifter
1. Medlemsstaterna skall säkerställa att det inte finns några rättsliga hinder inom deras jurisdiktion för att de fysiska och juridiska personer, vare sig dessa är reglerade enheter eller ej, som omfattas av extra tillsyn inbördes utbyter uppgifter som kan vara relevanta för den extra tillsynen.
2. Medlemsstaterna skall föreskriva att deras behöriga myndigheter med ansvar för att utöva extra tillsyn skall få tillgång till alla uppgifter som kan vara relevanta för den extra tillsynen, genom att direkt eller indirekt vända sig till enheterna i ett finansiellt konglomerat, vare sig dessa är reglerade enheter eller ej.
Artikel 15
Kontroll
Om de behöriga myndigheterna vid tillämpningen av detta direktiv i specifika fall önskar kontrollera uppgifter om en reglerad eller icke reglerad enhet i en annan medlemsstat vilken ingår i ett finansiellt konglomerat, skall de begära att de behöriga myndigheterna i denna medlemsstat låter utföra kontrollen.
De myndigheter som får en sådan begäran skall inom ramen för sin behörighet tillgodose begäran, antingen genom att själva utföra kontrollen, genom att låta en revisor eller expert utföra den eller genom att låta den begärande myndigheten själv utföra den.
Den behöriga myndighet som har framställt begäran får om den så önskar delta i kontrollen, om den inte själv utför den.
Artikel 16
Verkställande åtgärder
Om de reglerade enheterna i ett finansiellt konglomerat inte uppfyller de krav som anges i artiklarna 6-9 eller om kraven är uppfyllda men enheternas solvens ändå kan vara hotad eller om transaktionerna inom det finansiella konglomeratet eller riskkoncentrationerna utgör ett hot mot de reglerade enheternas finansiella ställning, skall nödvändiga åtgärder vidtas för att avhjälpa situationen så snart som möjligt
- av samordnaren när det gäller det blandade finansiella holdingföretaget,
- av de behöriga myndigheterna när det gäller reglerade enheter. I detta syfte skall samordnaren underrätta de behöriga myndigheterna om sina upptäckter.
Utan att det påverkar tillämpningen av artikel 17.2 får medlemsstaterna bestämma vilka åtgärder som deras behöriga myndigheter får vidta när det gäller blandade finansiella holdingföretag.
Då så krävs skall de berörda behöriga myndigheterna, inklusive samordnaren, samordna sina tillsynsåtgärder.
Artikel 17
De behöriga myndigheternas ytterligare befogenheter
1. I avvaktan på ytterligare harmonisering av särreglerna skall medlemsstaterna se till att de behöriga myndigheterna har befogenhet att vidta alla tillsynsåtgärder som anses nödvändiga för att undvika eller bemöta att reglerade enheter i ett finansiellt konglomerat kringgår särreglerna.
2. Utan att det påverkar tillämpningen av nationella straffrättsliga bestämmelser skall medlemsstaterna se till att påföljder eller åtgärder, vars syfte är att konstaterade överträdelser eller orsakerna till desamma skall upphöra, kan utdömas respektive vidtas gentemot blandade finansiella holdingföretag eller deras faktiska ledare, när dessa bryter mot lagar och andra författningar som antagits för att genomföra bestämmelserna i detta direktiv. I vissa fall kan sådana åtgärder kräva domstols medverkan. De behöriga myndigheterna skall ha ett nära samarbete för att se till att dessa påföljder och åtgärder får avsedd effekt.
AVSNITT 4
TREDJE LÄNDER
Artikel 18
Moderföretag utanför gemenskapen
1. Utan att detta påverkar särreglerna skall de behöriga myndigheterna i det fall som avses i artikel 5.3 kontrollera huruvida reglerade enheter, vilkas moderföretag har huvudkontor utanför gemenskapen, är föremål för sådan tillsyn som utövas av en behörig myndighet i tredje land som är likvärdig med den extra tillsyn som föreskrivs i detta direktiv beträffande sådana reglerade enheter som avses i artikel 5.2. Kontrollen skall utföras av den behöriga myndighet som skulle vara samordnare om kriterierna i artikel 10.2 hade varit tillämpliga, på begäran av moderföretaget eller av någon av de reglerade enheter som auktoriserats i gemenskapen eller på egen begäran. Den behöriga myndigheten skall samråda med de andra relevanta behöriga myndigheterna och beakta varje tillämplig vägledning som Kommittén för finansiella konglomerat har utarbetat enligt artikel 21.5. Den behöriga myndigheten skall med anledning därav rådfråga kommittén innan beslut fattas.
2. I brist på sådan likvärdig tillsyn som avses i punkt 1 skall de behöriga myndigheterna på dessa reglerade myndigheter analogt tillämpa de bestämmelser om extra tillsyn över reglerade enheter som avses i artikel 5.2. Alternativt får de behöriga myndigheterna tillämpa en av de metoder som anges i punkt 3.
3. Medlemsstaterna skall tillåta sina behöriga myndigheter att tillämpa andra metoder som säkerställer lämplig extra tillsyn över reglerade enheter i ett finansiellt konglomerat. Metoderna måste godkännas av samordnaren, efter samråd med de andra relevanta behöriga myndigheterna. De behöriga myndigheterna kan särskilt kräva att det inrättas ett blandat finansiellt holdingföretag med huvudkontor inom gemenskapen och tillämpa detta direktiv på de reglerade enheterna i det finansiella konglomerat som leds av detta holdingföretag. Metoderna skall uppfylla de mål för den extra tillsynen som ställs upp i detta direktiv och skall rapporteras till de andra berörda behöriga myndigheterna och kommissionen.
Artikel 19
Samarbete med behöriga myndigheter i tredje land
1. Artikel 25.1 och 25.2 i direktiv 2000/12/EG och artikel 10a i direktiv 98/78/EG skall även tillämpas vid förhandlingar om avtal med ett eller flera tredje länder rörande metoder för utövande av extra tillsyn över reglerade enheter i ett finansiellt konglomerat.
2. Kommissionen, Rådgivande bankrörelsekommittén, Försäkringskommittén och Kommittén för finansiella konglomerat skall granska resultatet av de förhandlingar som avses i punkt 1 och den därigenom uppkomna situationen.
KAPITEL III
KOMMISSIONENS BEFOGENHETER OCH KOMMITTÉFÖRFARANDE
Artikel 20
Kommissionens befogenheter
1. Kommissionen skall, i enlighet med det förfarande som avses i artikel 21.2, anta tekniska ändringar av detta direktiv på följande områden:
a) En mer precis formulering av definitionerna i artikel 2 i syfte att beakta utvecklingen på finansmarknaderna vid tillämpningen av detta direktiv.
b) En mer precis formulering av definitionerna i artikel 2 i syfte att säkerställa en enhetlig tillämpning av detta direktiv i gemenskapen.
c) Harmonisering av terminologin och ramarna för definitionerna i direktivet i överensstämmelse med framtida gemenskapsrättsakter om reglerade enheter och närliggande frågor.
d) En mer precis definition av beräkningsmetoderna i bilaga I för att beakta utvecklingen på finansmarknaderna och av tillsynsmetoderna.
e) Samordning av bestämmelserna enligt artiklarna 7 och 8 och bilaga II, så att enhetlig tillämpning inom gemenskapen uppmuntras.
2. Kommissionen skall underrätta allmänheten om alla förslag som läggs fram i enlighet med denna artikel och kommer att samråda med de berörda parterna, innan den överlämnar utkastet till åtgärder till den kommitté för finansiella konglomerat som anges i artikel 21.
Artikel 21
Kommitté
1. Kommissionen skall bistås av en kommitté för finansiella konglomerat, nedan kallad "kommittén".
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning.
4. Utan att det påverkar redan antagna genomförandeåtgärder, skall tillämpningen av de bestämmelser i detta direktiv i vilka föreskrivs att tekniska regler och beslut skall antas i enlighet med förfarandet i punkt 2 upphöra fyra år efter det att detta direktiv har trätt i kraft. Europaparlamentet och rådet kan på förslag av kommissionen förnya bestämmelserna i fråga i enlighet med förfarandet i artikel 251 i fördraget och skall därvid granska dem före utgången av ovannämnda period.
5. Kommittén får ge allmän vägledning om huruvida det är sannolikt att de system för extra tillsyn som tillämpas av behöriga myndigheter i tredje land kommer att uppfylla det mål för den extra tillsynen som ställs upp i detta direktiv, när det gäller reglerade enheter i ett finansiellt konglomerat vars ledande enhet har sitt huvudkontor utanför gemenskapen. Kommittén skall fortlöpande se över all sådan vägledning och beakta varje förändring i den extra tillsyn som utförs av sådana behöriga myndigheter.
6. Kommittén skall hållas underrättad av medlemsstaterna om de principer som de tillämpar för tillsynen över transaktioner inom det finansiella konglomeratet och riskkoncentration.
KAPITEL IV
ÄNDRINGAR AV NUVARANDE DIREKTIV
Artikel 22
Ändringar av direktiv 73/239/EEG
Direktiv 73/239/EEG ändras på följande sätt:
1. Följande artikel skall läggas till:
"Artikel 12a
1. Samråd med behöriga myndigheter i den andra berörda medlemsstaten skall genomföras innan auktorisation beviljas för ett försäkringsföretag som
a) är dotterföretag till ett försäkringsföretag som är auktoriserat i en annan medlemsstat,
b) är dotterföretag till moderföretaget till ett försäkringsföretag som är auktoriserat i en annan medlemsstat, eller
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett försäkringsföretag som är auktoriserat i en annan medlemsstat.
2. Samråd med den behöriga myndigheten i en berörd medlemsstat som ansvarar för tillsynen över kreditinstitut eller värdepappersföretag skall genomföras innan auktorisation beviljas för ett försäkringsföretag som
a) är dotterföretag till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen,
b) är dotterföretag till moderföretaget till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen, eller
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen.
3. De relevanta behöriga myndigheter som avses i punkterna 1 och 2 skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla de uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet som är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
2. I artikel 16.2 skall följande stycken läggas till:
"Från den disponibla solvensmarginalen skall även följande dras:
a) Ägarintressen som försäkringsföretaget har i
- försäkringsföretag i den mening som avses i artikel 6 i detta direktiv, artikel 6 i första direktivet 79/267/EEG av den 5 mars 1979 om samordning av lagar och andra författningar om rätten att starta och driva direkt livförsäkringsrörelse(17) eller artikel 1 b i Europaparlamentets och rådets direktiv 98/78/EG(18),
- återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG,
- försäkringsholdingbolag i den mening som avses i artikel 1 led i i direktiv 98/78/EG,
- kreditinstitut och finansiella institut i den mening som avses i artiklarna 1.1 och 1.5 i Europaparlamentets och rådets direktiv 2000/12/EG(19),
- värdepappersföretag och finansiella institut i den mening som avses i artikel 1.2 i direktiv 93/22/EEG(20) och i artiklarna 2.4 och 2.7 i rådets direktiv 93/6/EEG(21).
b) Var och en av följande poster som ett försäkringsföretag innehar i de enheter som definierats i a i vilka det har ägarintresse:
- De instrument som avses i punkt 3.
- De instrument som avses i artikel 18.3 i direktiv 79/267/EEG.
- Fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 i direktiv 2000/12/EG.
Om aktier i ett annat kreditinstitut, värdepappersföretag, finansiellt institut, försäkringsföretag, återförsäkringsföretag eller försäkringsholdingbolag innehas tillfälligt i syfte att ge finansiellt bistånd för att rekonstruera och rädda denna enhet, får den behöriga myndigheten bevilja undantag från bestämmelserna om avdrag enligt a och b i fjärde stycket.
Som ett alternativ till avdrag av de poster enligt a och b i fjärde stycket som försäkringsföretag innehar i kreditinstitut, värdepappersföretag och finansiella institut, får medlemsstaterna tillåta att deras försäkringsföretag också tillämpar metoderna 1, 2 eller 3 i bilaga I till Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(22). Metod 1 (metod baserad på sammanställd redovisning) skall tillämpas endast om den behöriga myndigheten är säker på graden av samordnad förvaltning och intern kontroll avseende de enheter som skall inbegripas i tillämpningsområdet för sammanställningen. Den valda metoden skall tillämpas konsekvent över tiden.
För beräkningen av solvensmarginalen enligt detta direktiv får medlemsstaterna föreskriva att försäkringsföretag som är föremål för extra tillsyn enligt direktiv 98/78/EG eller direktiv 2002/87/EG inte behöver dra ifrån poster enligt a och b i fjärde stycket i de kreditinstitut, värdepappersföretag, finansiella institut, försäkrings- eller återförsäkringsföretag eller försäkringsholdingbolag som ingår i den extra tillsynen.
Med det avdrag av ägarintresse som anges i detta stycke menas här ägarintresse i den mening som avses i artikel 1 f i direktiv 98/78/EG.".
Artikel 23
Ändringar av direktiv 79/267/EEG
Direktiv 79/267/EEG ändras på följande sätt:
1. Följande artikel skall läggas till:
"Artikel 12a
1. Samråd med behöriga myndigheter i den andra berörda medlemsstaten skall genomföras innan auktorisation beviljas för ett livförsäkringsföretag som
a) är dotterföretag till ett försäkringsföretag som är auktoriserat i en annan medlemsstat,
b) är dotterföretag till moderföretaget till ett försäkringsföretag som är auktoriserat i en annan medlemsstat, eller
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett försäkringsföretag som är auktoriserat i en annan medlemsstat.
2. Samråd med den behöriga myndighet som ansvarar för tillsynen över kreditinstitut eller värdepappersföretag skall genomföras innan auktorisation beviljas för ett livförsäkringsföretag som
a) är dotterföretag till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen,
b) är dotterföretag till moderföretaget till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen, eller
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen.
3. De relevanta behöriga myndigheter som avses i punkterna 1 och 2 skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla de uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet som är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
2. I artikel 18.2 skall följande stycken läggas till:
"Från den disponibla solvensmarginalen skall även följande avdrag göras:
a) Ägarintressen som försäkringsföretaget har i
- försäkringsföretag i den mening som avses i artikel 6 i detta direktiv, artikel 6 i direktiv 73/239/EEG(23)eller artikel 1 b i Europaparlamentets och rådets direktiv 98/78/EG(24),
- återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG,
- försäkringsholdingbolag i den mening som avses i artikel 1 led i i direktiv 98/78/EG,
- kreditinstitut och finansiella institut i den mening som avses i artiklarna 1.1 och 1.5 i Europaparlamentets och rådets direktiv 2000/12/EG(25),
- värdepappersföretag och finansiella institut i den mening som avses i artikel 1.2 i direktiv 93/22/EEG(26) och i artiklarna 2.4 och 2.7 i direktiv 93/6/EEG(27).
b) Var och en av följande poster som ett försäkringsföretag innehar i de enheter som definierats under a i vilka det har ägarintresse:
- De instrument som avses i punkt 3.
- De instrument som avses i artikel 16.3 i direktiv 73/239/EEG.
- Fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 i direktiv 2000/12/EG.
För beräkningen av solvensmarginalen enligt detta direktiv får medlemsstaterna föreskriva att försäkringsföretag som är föremål för extra tillsyn enligt direktiv 98/78/EG eller enligt direktiv 2002/87/EG inte behöver dra ifrån poster enligt a och b i tredje stycket i de kreditinstitut, värdepappersföretag, finansiella institut, försäkrings- eller återförsäkringsföretag eller försäkringsholdingbolag som ingår i den extra tillsynen.
Med det avdrag av ägarintresse som anges i denna punkt menas här ägarintresse i den mening som avses i artikel 1 f i direktiv 98/78/EG.".
Artikel 24
Ändring av direktiv 92/49/EEG
Direktiv 92/49/EEG ändras på följande sätt:
1. I artikel 15 skall följande punkt införas:
"1a. Om köparen av det innehav som avses i punkt 1 är ett försäkringsföretag, ett kreditinstitut eller ett värdepappersföretag med auktorisation i en annan medlemsstat eller moderföretag till en sådan enhet, eller en fysisk eller juridisk person som har ägarkontroll över en sådan enhet, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av ett sådant samråd som avses i artikel 12a i direktiv 73/239/EEG.".
2. Artikel 16.5c skall ersättas med följande:
"5c. Denna artikel skall inte hindra en behörig myndighet från att
- till centralbanker och andra organ med liknande funktion i egenskap av monetära myndigheter,
- i förekommande fall till andra myndigheter med ansvar för övervakning av betalningssystem,
överföra uppgifter för att dessa skall kunna utföra sina uppgifter, och den skall inte heller hindra sådana myndigheter eller organ från att vidarebefordra sådana uppgifter som de kan behöva enligt punkt 4. Uppgifter som erhålls i detta sammanhang skall omfattas av de bestämmelser om tystnadsplikt som fastställs i denna artikel.".
Artikel 25
Ändring av direktiv 92/96/EEG
Direktiv 92/96/EEG skall ändras på följande sätt:
1. I artikel 14 skall följande punkt införas:
"1a. Om köparen av det innehav som avses i punkt 1 är ett försäkringsföretag, ett kreditinstitut eller ett värdepappersföretag med auktorisation i en annan medlemsstat eller moderföretag till en sådan enhet, eller en fysisk eller juridisk person som har ägarkontroll över en sådan enhet, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av ett sådant samråd som avses i artikel 12a i direktiv 79/267/EEG.".
2. Artikel 15.5c skall ersättas med följande:
"5c. Denna artikel skall inte hindra en behörig myndighet från att
- till centralbanker och andra organ med liknande funktion i egenskap av monetära myndigheter,
- i förekommande fall till andra myndigheter med ansvar för övervakning av betalningssystem,
överföra uppgifter för att dessa skall kunna utföra sina uppgifter, och den skall inte heller hindra sådana myndigheter eller organ från att vidarebefordra sådana uppgifter som de kan behöva enligt punkt 4. Uppgifter som erhålls i detta sammanhang skall omfattas av de bestämmelser om tystnadsplikt som fastställs i denna artikel.".
Artikel 26
Ändring av direktiv 93/6/EEG
I artikel 7.3 i direktiv 93/6/EEG skall första och andra strecksatsen ersättas med följande text:
"- finansiellt holdingföretag: ett finansiellt institut vars dotterföretag antingen uteslutande eller huvudsakligen är värdepappersföretag eller andra finansiella institut av vilka åtminstone ett är ett värdepappersföretag, vilket inte är ett finansiellt holdingföretag med blandad verksamhet i den mening som avses i Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(29).
- holdingföretag med blandad verksamhet: ett moderföretag som inte utgör ett finansiellt holdingföretag, ett värdepappersföretag eller ett blandat finansiellt holdingföretag i den mening som avses i direktiv 2002/87/EG, bland vars dotterföretag det finns minst ett värdepappersföretag.".
Artikel 27
Ändringar av direktiv 93/22/EEG
Direktiv 93/22/EEG ändras på följande sätt:
1. I artikel 6 skall följande stycken läggas till:
"Samråd med den behöriga myndighet i en berörd medlemsstat som har ansvar för tillsynen över kreditinstitut eller försäkringsföretag skall genomföras innan auktorisation beviljas för ett värdepappersföretag som
a) är dotterföretag till ett kreditinstitut eller försäkringsföretag som är auktoriserat i gemenskapen,
b) är dotterföretag till moderföretaget till ett kreditinstitut eller försäkringsföretag som är auktoriserat i gemenskapen, eller
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett kreditinstitut eller ett försäkringsföretag som är auktoriserat i gemenskapen.
De relevanta behöriga myndigheter som avses i första och andra stycket skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla de uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet som är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
2. Artikel 9.2 skall ersättas med följande:
"2. Om förvärvaren av det innehav som avses i punkt 1 är ett värdepappersföretag, ett kreditinstitut eller ett försäkringsföretag med auktorisation i en annan medlemsstat eller moderföretag till ett värdepappersföretag, ett kreditinstitut eller ett försäkringsföretag med auktorisation i en annan medlemsstat, eller en fysisk eller juridisk person som har ägarkontroll över ett värdepappersföretag, ett kreditinstitut eller ett försäkringsföretag med auktorisation i en annan medlemsstat, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av sådant samråd som avses i artikel 6.".
Artikel 28
Ändringar i direktiv 98/78/EG
Direktiv 98/78/EG ändras på följande sätt:
1. I artikel 1 skall g, h, i och j ersättas med följande:
"g) företag med ägarintresse: ett företag som är antingen moderföretag eller ett annat företag som har ett ägarintresse eller ett företag som är knutet till ett annat företag genom ett sådant förhållande som avses i artikel 12.1 i direktiv 83/349/EEG.
h) anknutet företag: ett företag som är antingen ett dotterföretag eller ett annat företag som är föremål för ägarintresse eller ett företag som är knutet till ett annat företag genom ett sådant förhållande som avses i artikel 12.1 i direktiv 83/349/EEG.
i) försäkringsholdingbolag: ett moderföretag vars huvudsakliga verksamhet består i att förvärva och ha ägarintresse i dotterföretag, vilka enbart eller huvudsakligen är försäkringsföretag, återförsäkringsföretag eller försäkringsföretag i tredje land, där minst ett av dotterföretagen är ett försäkringsföretag, och vilket inte är ett blandat finansiellt holdingföretag i den mening som avses i Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(30).
j) försäkringsholdingföretag med blandad verksamhet: ett annat moderföretag än ett försäkringsföretag, ett försäkringsföretag i tredje land, ett återförsäkringsföretag, ett försäkringsholdingföretag eller ett blandat finansiellt holdingföretag i den mening som avses i direktiv 2002/87/EG, vilket har minst ett försäkringsföretag bland sina dotterföretag.".
2. I artikel 6.3 skall följande mening läggas till:
"Den behöriga myndighet som har framställt begäran får om den så önskar delta i kontrollen, om den inte själv utför den.".
3. I artikel 8.2 skall det första stycket ersättas med följande:
"Medlemsstaterna skall kräva att försäkringsföretagen följer adekvata metoder för riskhantering och rutiner för intern kontroll, inbegripet sunda rapporterings- och redovisningsförfaranden, för att på ett lämpligt sätt identifiera, mäta, övervaka och kontrollera transaktioner enligt bestämmelserna i punkt 1. Medlemsstaterna skall också kräva att försäkringsföretagen minst en gång om året rapporterar betydande transaktioner till de behöriga myndigheterna. Dessa förfaranden och betydande transaktioner skall övervakas av de behöriga myndigheterna.".
4. Följande artiklar skall läggas till:
"Artikel 10a
Samarbete med behöriga myndigheter i tredje land
1. Kommissionen kan antingen på begäran av en medlemsstat eller på eget initiativ ställa förslag till rådet i fråga om förhandlingar om avtal med ett eller flera tredje länder om metoderna för att utöva extra tillsyn över
a) försäkringsföretag bland vars delägare det finns företag i den mening som avses i artikel 2 med huvudkontor i tredje land, och
b) försäkringsföretag i ett icke-medlemsland bland vars delägare det finns företag i den mening som avses i artikel 2 med huvudkontor inom gemenskapen.
2. Av de avtal som avses i punkt 1 skall särskilt framgå både
a) att de behöriga myndigheterna i medlemsstaterna kan få fram den information som krävs för att utöva extra tillsyn över försäkringsföretag med huvudkontor inom gemenskapen och med dotterföretag eller ägarintressen i företag utanför gemenskapen, och
b) att de behöriga myndigheterna i tredje land kan få fram den information som krävs för att utöva extra tillsyn över försäkringsföretag med huvudkontor inom deras territorier och med dotterföretag eller ägarintressen i företag i en eller flera medlemsstater.
3. Kommissionen och Försäkringskommittén skall granska resultaten av de förhandlingar som avses i punkt 1 och den därigenom uppkomna situationen.
Artikel 10b
Ledningsorgan för holdingföretag med blandad verksamhet
Medlemsstaterna skall kräva att de personer som faktiskt leder affärsverksamheten i ett holdingföretag med blandad verksamhet har ett tillräckligt gott anseende och tillräcklig erfarenhet för att kunna fullgöra dessa åligganden.".
5. I punkt 1 B i bilaga I skall följande stycke läggas till:
"Om det inte finns några kapitalband mellan vissa av företagen i en försäkringsgrupp, skall den behöriga myndigheten fastställa vilken proportionell andel som det skall tas hänsyn till.".
6. I punkt 2 i bilaga I skall följande punkt läggas till:
"2.4a Berörda kreditinstitut, värdepappersföretag och finansiella institut
Reglerna om avdrag av ett sådant ägarintresse enligt artikel 16.1 i direktiv 73/239/EEG och artikel 18 i direktiv 79/267/EEG samt bestämmelserna om medlemsstaternas möjlighet att under vissa villkor tillåta alternativa metoder och att tillåta att ett sådant ägarintresse inte skall dras av, skall även tillämpas vid beräkningen av jämkad solvens hos ett försäkringsföretag som är ett företag med ägarintresse i ett kreditinstitut, ett värdepappersföretag eller ett finansiellt institut.".
Artikel 29
Ändringar av direktiv 2000/12/EG
Direktiv 2000/12/EG ändras på följande sätt:
1. Artikel 1 skall ändras på följande sätt:
a) Punkt 9 skall ersättas med följande:
"9. ägarintresse vid tillämpningen av gruppbaserad tillsyn och vid tillämpningen av artikel 34.2.15 och 34.2.16: ägarintresse i den mening som avses i artikel 17 första meningen i direktiv 78/660/EEG eller direkt eller indirekt innehav av 20 % eller mer av rösterna eller kapitalet i ett företag.".
b) Punkterna 21 och 22 skall ersättas med följande:
"21. finansiellt holdingföretag: ett finansiellt institut vars dotterföretag uteslutande eller huvudsakligen är kreditinstitut eller finansiella institut, varvid minst ett av dotterföretagen skall vara ett kreditinstitut, och som inte är ett blandat finansiellt holdingföretag i den mening som avses i Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(31).
22. holdingföretag med blandad verksamhet: ett moderföretag som inte är ett finansiellt holdingföretag, ett kreditinstitut eller ett blandat finansiellt holdingföretag i den mening som avses i direktiv 2002/87/EG, vilket har minst ett kreditinstitut bland sina dotterföretag.".
2. I artikel 12 skall följande stycken läggas till:
"Samråd med den behöriga myndighet som har ansvar för tillsynen över försäkringsföretag eller värdepappersföretag skall genomföras innan auktorisation beviljas för ett kreditinstitut som
a) är dotterföretag till ett försäkringsföretag som är auktoriserat i gemenskapen,
b) är dotterföretag till moderföretaget till ett försäkringsföretag som är auktoriserat i gemenskapen, eller
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett försäkringsföretag som är auktoriserat i gemenskapen.
De relevanta behöriga myndigheter som avses i första och andra stycket skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet vilka är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
3. Artikel 16.2 skall ersättas med följande:
"2. Om förvärvaren av det innehav som avses i punkt 1 är ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag med auktorisation i en annan medlemsstat eller moderföretag till ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag med auktorisation i en annan medlemsstat, eller en fysisk eller juridisk person som har ägarkontroll över ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag med auktorisation i en annan medlemsstat, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av sådant samråd som avses i artikel 12.".
4. Artikel 34.2 skall ändras på följande sätt:
a) I det första stycket skall punkterna 12 och 13 ersättas med följande:
"12. Sådana ägarposter i andra kreditinstitut och finansiella institut som motsvarar mer än 10 % av deras kapital.
13. Fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 som ett kreditinstitut innehar hos kreditinstitut och finansiella institut, i vilka kreditinstitutet har en ägarandel som i varje enskilt fall motsvarar mer än 10 % av kapitalet.
14. Ägarposter i andra kreditinstitut och finansiella institut, motsvarande högst 10 % av deras kapital, fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 som ett kreditinstitut innehar hos andra kreditinstitut och finansiella institut än de som anges i punkterna 12 och 13 i detta stycke, i den mån dessa ägarposter, fordringar och instrument tillsammans överstiger 10 % av kreditinstitutets kapitalbas beräknad före avdrag för posterna enligt punkterna 12-16 i detta stycke.
15. Ägarintresse av det slag som avses i artikel 1.9, vilket ett kreditinstitut innehar i
- försäkringsföretag i den mening som avses i artikel 6 i direktiv 73/239/EEG, artikel 6 i direktiv 79/267/EEG eller artikel 1 b i Europaparlamentets och rådets direktiv 98/78/EG(32),
- återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG,
- försäkringsholdingföretag i den mening som avses i artikel 1 led i i direktiv 98/78/EG.
16. Var och en av följande poster som ett kreditinstitut innehar i de enheter som definieras i punkt 15 i vilka det har ägarintresse
- de instrument som avses i artikel 16.3 i direktiv 73/239/EEG,
- de instrument som avses i artikel 18.3 i direktiv 79/267/EEG.".
b) Andra stycket skall ersättas med följande:
"Om aktier i ett annat kreditinstitut, finansiellt institut, försäkringsföretag, återförsäkringsföretag eller försäkringsholdingföretag innehas tillfälligt i syfte att ge finansiellt bistånd för att rekonstruera och rädda denna enhet, får den behöriga myndigheten bevilja undantag från bestämmelserna om avdrag i punkterna 12-16.
Som ett alternativ till avdrag av poster enligt punkterna 15 och 16 får medlemsstaterna tillåta att deras kreditinstitut också tillämpar metoderna 1, 2 eller 3 i bilaga I i direktiv 2002/87/EG. Metod 1 (metod baserad på sammanställd redovisning) skall endast tillämpas om den behöriga myndigheten är säker på graden av samordnad förvaltning och intern kontroll avseende de enheter som skall inbegripas i tillämpningsområdet för sammanställningen. Den valda metoden skall tillämpas konsekvent över tiden.
Medlemsstaterna får föreskriva att kreditinstitut som är föremål för gruppbaserad tillsyn enligt kapitel 3 eller extra tillsyn enligt ovan nämnda direktiv 2002/87/EG, vid beräkning av den egna icke gruppbaserade kapitalbasen inte behöver dra ifrån poster enligt punkterna 15 och 16 i de kreditinstitut, finansiella institut eller försäkrings- eller återförsäkringsföretag eller försäkringsholdingföretag som omfattas av den gruppbaserade tillsynen eller av den extra tillsynen.
Denna bestämmelse skall tillämpas på alla försiktighetsregler som är harmoniserade genom gemenskapsakten.".
5. Artikel 51.3 skall ersättas med följande:
"3. Medlemsstaterna behöver inte tillämpa begränsningarna enligt punkterna 1 och 2 för ägarposter i försäkringsföretag enligt definitionen i direktiv 73/239/EEG och direktiv 79/267/EEG eller i återförsäkringsföretag enligt definitionen i direktiv 98/78/EG.".
6. Artikel 52.2 sista meningen skall ersättas med följande:
"Utan att det påverkar tillämpningen av artikel 54a skall sammanställningen inte på något sätt anses innebära att de behöriga myndigheterna har skyldighet att utöva tillsyn i förhållande till det enskilda finansiella holdingföretaget.".
7. Artikel 54 skall ändras på följande sätt:
a) I punkt 1 skall följande stycke läggas till:
"Om företagen står i ett sådant samband som avses i artikel 12.1 i direktiv 83/349/EEG skall de behöriga myndigheterna bestämma hur sammanställningen skall ske.".
b) I punkt 4 första stycket skall tredje strecksatsen utgå.
8. Följande artikel skall införas:
"Artikel 54a
Ledningsorgan för finansiella holdingföretag
Medlemsstaterna skall kräva att de personer som faktiskt leder affärsverksamheten i ett finansiellt holdingföretag har ett tillräckligt gott anseende och tillräcklig erfarenhet för att kunna fullgöra dessa åligganden.".
9. Följande artikel skall läggas till:
"Artikel 55a
Transaktioner inom det finansiella konglomeratet med holdingföretag med blandad verksamhet
Utan att detta påverkar bestämmelserna i avdelning V kapitel 2 avsnitt 3 i detta direktiv skall medlemsstaterna, då moderföretaget till ett eller flera kreditinstitut är ett holdingföretag med blandad verksamhet, se till att de behöriga myndigheter som ansvarar för tillsynen över dessa kreditinstitut utövar allmän tillsyn över transaktioner mellan kreditinstitutet och holdingföretaget med blandad verksamhet samt dess dotterföretag.
De behöriga myndigheterna skall kräva att kreditinstituten följer adekvata metoder för riskhantering och rutiner för intern kontroll, inbegripet sunda rapporterings- och redovisningsförfaranden, för att på ett lämpligt sätt identifiera, mäta, övervaka och kontrollera transaktionerna med det holdingföretag med blandad verksamhet som är moderföretag och dess dotterföretag. De behöriga myndigheterna skall kräva att kreditinstituten rapporterar varje annan betydande transaktion med dessa enheter än den som avses i artikel 48. Dessa förfaranden och betydande transaktioner skall övervakas av de behöriga myndigheterna.
Om ovannämnda transaktioner inom det finansiella konglomeratet utgör ett hot mot kreditinstitutets finansiella ställning, skall den behöriga myndighet som ansvarar för tillsynen över institutet vidta lämpliga åtgärder.".
10. I artikel 56.7 skall följande mening läggas till:
"Den behöriga myndighet som har framställt begäran får om den så önskar delta i kontrollen, om den inte själv utför den.".
11. Följande artikel skall läggas till:
"Artikel 56a
Moderföretag i tredje land
Om ett kreditinstitut, vars moderföretag är ett kreditinstitut eller ett finansiellt holdingföretag med huvudkontor utanför gemenskapen, inte är föremål för gruppbaserad tillsyn enligt artikel 52, skall de behöriga myndigheterna kontrollera huruvida kreditinstitutet är föremål för gruppbaserad tillsyn av en behörig myndighet i tredje land, vilken är likvärdig med den som styrs av de principer som anges i artikel 52. Kontrollen skall utföras av den behöriga myndighet som skulle vara ansvarig för den extra tillsynen om fjärde stycket hade varit tillämpligt, på begäran av moderföretaget eller av någon av de reglerade enheter som auktoriserats i gemenskapen eller på eget initiativ. Denna behöriga myndighet skall samråda med de andra berörda behöriga myndigheterna.
Den rådgivande bankrörelsekommittén får ge allmän vägledning om huruvida det är sannolikt att de system för gruppbaserad tillsyn som tillämpas av behöriga myndigheter i tredje land kommer att uppfylla de mål för den gruppbaserade tillsynen som ställs upp i detta kapitel, när det gäller kreditinstitut vars moderföretag har sitt huvudkontor utanför gemenskapen. Kommittén skall fortsätta att se över all sådan vägledning och beakta varje förändring i de system för den gruppbaserade tillsynen som tillämpas av sådana behöriga myndigheter.
Alternativt skall medlemsstaterna tillåta sina behöriga myndigheter att använda andra lämpliga metoder för tillsyn vilka uppfyller målen för den gruppbaserade tillsynen över kreditinstitut. De myndigheter som skulle vara ansvariga för gruppbaserad tillsyn måste enas om dessa metoder efter att ha samrått med andra berörda behöriga myndigheter. De behöriga myndigheterna kan särskilt kräva att det inrättas ett finansiellt holdingföretag med huvudkontor inom gemenskapen och tillämpa bestämmelserna om gruppbaserad tillsyn på det finansiella holdingföretagets ställning på gruppnivå. Metoderna måste uppfylla de mål för den gruppbaserade tillsynen som ställs upp i detta kapitel och rapporteras till de andra berörda behöriga myndigheterna och kommissionen.".
KAPITEL V
KAPITALFÖRVALTNINGSBOLAG
Artikel 30
Kapitalförvaltningsbolag
Till dess att särreglerna har samordnats ytterligare skall medlemsstaterna föreskriva att kapitalförvaltningsbolag skall omfattas av
a) tillämpningsområdet för gruppbaserad tillsyn av kreditinstitut eller värdepappersföretag och/eller tillämpningsområdet för extra tillsyn över sådana försäkringsföretag som ingår i en försäkringsgrupp, och
b) tillämpningsområdet för extra tillsyn i den mening som avses i detta direktiv, om gruppen är ett finansiellt konglomerat.
För tillämpningen av det första stycket skall medlemsstaterna föreskriva eller ge sina behöriga myndigheter behörighet att besluta om enligt vilka särregler (för banksektorn, försäkringssektorn eller värdepapperssektorn) kapitalförvaltningsbolag skall omfattas av den gruppbaserade tillsyn och/eller den extra tillsyn som avses i första stycket a. I denna bestämmelse skall särreglerna om i vilken form och utsträckning finansiella institut (om kapitalförvaltningsbolag omfattas av tillämpningsområdet för gruppbaserad tillsyn över kreditinstitut och värdepappersföretag) och återförsäkringsföretag (om kapitalförvaltningsbolag omfattas av tillämpningsområdet för extra tillsyn över försäkringsföretag) skall omfattas också tillämpas på kapitalförvaltningsbolag. Vad avser den extra tillsyn som avses i första stycket b skall kapitalförvaltningsbolaget behandlas som en del av den sektor som det skall räknas till i enlighet med första stycket a.
Om ett kapitalförvaltningsbolag utgör en del av ett finansiellt konglomerat skall hänvisningar till begreppet reglerad enhet och till begreppet behöriga myndigheter och relevanta behöriga myndigheter i detta direktiv anses inbegripa kapitalförvaltningsbolag respektive de behöriga myndigheter som ansvarar för tillsynen över kapitalförvaltningsbolag. Detta skall också tillämpas på sådana grupper som avses i första stycket a.
KAPITEL VI
ÖVERGÅNGS- OCH SLUTBESTÄMMELSER
Artikel 31
Rapport från kommissionen
1. Senast 11 augusti 2007 skall kommissionen till den kommitté för finansiella konglomerat som avses i artikel 21 överlämna en rapport om medlemsstaternas praxis och i förekommande fall om behovet av ytterligare harmonisering i fråga om
- huruvida kapitalförvaltningsbolag bör omfattas av tillsynen på gruppnivå,
- vilka kapitaltäckningsmetoder i bilaga I som bör väljas och hur de bör tillämpas,
- hur betydande transaktioner inom det finansiella konglomeratet och betydande riskkoncentration bör definieras samt om tillsynen över transaktioner inom det finansiella konglomeratet och riskkoncentration som avses i bilaga II, särskilt i fråga om införandet av kvantitativa gränser och kvalitativa krav i detta syfte,
- hur ofta finansiella konglomerat skall beräkna kapitaltäckningskraven enligt artikel 6.2 och rapportera till samordnaren om betydande riskkoncentrationer enligt artikel 7.2.
Kommissionen skall samråda med kommittén innan den lägger fram sina förslag.
2. Inom ett år efter det att en överenskommelse träffats på internationell nivå om bestämmelserna om eliminering av dubbelt utnyttjande av poster i kapitalbasen i finansiella grupper skall kommissionen undersöka hur bestämmelserna i detta direktiv kan anpassas till dessa internationella överenskommelser och vid behov lägga fram lämpliga förslag.
Artikel 32
Införlivande
När medlemsstaterna antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare bestämmelser om hur denna hänvisning skall göras skall varje medlemsstat själv utfärda.
Artikel 33
Ikraftträdande
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska unionens officiella tidning.
Artikel 34
Adressater
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens direktiv 2002/97/EG
av den 16 december 2002
om ändring av bilagorna till rådets direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG beträffande fastställande av gränsvärden för bekämpningsmedelsrester (2,4-D, triasulfuron och tifensulfuronmetyl) i och på spannmål, livsmedel av animaliskt ursprung och vissa produkter av vegetabiliskt ursprung, inklusive frukt och grönsaker
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 86/362/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på spannmål(1), senast ändrat genom kommissionens direktiv 2002/79/EG(2), särskilt artikel 10 i detta,
med beaktande av rådets direktiv 86/363/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på livsmedel av animaliskt ursprung(3), senast ändrat genom direktiv 2002/79/EG, särskilt artikel 10 i detta,
med beaktande av rådets direktiv 90/642/EEG av den 27 november 1990 om fastställande av gränsvärden för bekämpningsmedelsrester i och på produkter av vegetabiliskt ursprung inklusive frukt och grönsaker(4), senast ändrat genom direktiv 2002/79/EG, särskilt artikel 7 i detta,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(5), senast ändrat genom kommissionens direktiv 2002/81/EG(6), särskilt artikel 4.1 f i detta, och
av följande skäl:
(1) Genom kommissionens direktiv 2001/103/EG(7), 2000/66/EG(8) respektive 2001/99/EG(9) infördes de befintliga verksamma ämnena 2,4-D, triasulfuron och tifensulfuronmetyl i bilaga I till direktiv 91/414/EEG för att användas som herbicider, utan att det angavs några särskilda förhållanden som skulle kunna inverka på grödor som eventuellt behandlades med växtskyddsmedel innehållande dessa verksamma ämnen.
(2) Nämnda införande i bilaga I till direktiv 91/414/EEG av dessa verksamma ämnen grundades på en utvärdering av de uppgifter som lämnats in om det föreslagna användningsområdet. Uppgifterna om användningen har lämnats in av vissa medlemsstater i enlighet med artikel 4.1 f i direktiv 91/414/EEG. Tillgängliga uppgifter har nu gåtts igenom, och de har befunnits vara tillräckliga för att vissa gränsvärden för bekämpningsmedelsrester skall kunna fastställas.
(3) Om det inte finns något permanent eller provisoriskt gränsvärde för bekämpningsmedelsrester på gemenskapsnivå måste medlemsstaterna fastställa ett provisoriskt nationellt gränsvärde i enlighet med artikel 4.1 f i direktiv 91/414/EEG innan växtskyddsmedel som innehåller detta verksamma ämne kan godkännas.
(4) I samband med införandet av de berörda verksamma ämnena i bilaga I till direktiv 91/414/EEG avslutades de tekniska och vetenskapliga utvärderingarna genom kommissionens granskningsrapport. Rapporten avslutades den 2 oktober 2001 för 2,4-D, den 13 juli 2000 för triasulfuron och den 29 juni 2001 för tifensulfuronmetyl. I rapporterna fastställs det acceptabla dagliga intaget (ADI) för 2,4-D till 0,05 mg per kg kroppsvikt och dag, för triasulfuron till 0,01 mg per kg kroppsvikt och dag och för tifensulfuronmetyl till 0,01 mg per kg kroppsvikt och dag. Konsumenternas livstidsexponering genom livsmedel som behandlats med de berörda verksamma ämnena har uppskattats och utvärderats med hjälp av de metoder som används inom gemenskapen. Hänsyn har också tagits till de riktlinjer som offentliggjorts av Världshälsoorganisationen(10) samt yttrandet om de använda metoderna från den Vetenskapliga kommittén för växter(11). Det har fastslagits att de föreslagna gränsvärdena inte leder till att de acceptabla dagliga intagen överskrids. Under de utvärderingar och diskussioner som föregick införandet av de berörda verksamma ämnena i bilaga I till direktiv 91/414/EEG noterades inga akuta toxiska effekter som skulle kräva att det fastställs en akut referensdos.
(5) För att konsumenterna skall kunna skyddas från exponering av bekämpningsmedelsrester i eller på produkter som inte har godkänts, bör de provisoriska gränsvärden som fastställs motsvara den lägsta analytiska bestämningsgränsen för samtliga produkter som omfattas av direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG.
(6) Även om gemenskapen fastställer sådana provisoriska gränsvärden hindrar detta inte att medlemsstaterna själva fastställer provisoriska gränsvärden enligt artikel 4.1 f i direktiv 91/414/EEG och bilaga VI till det direktivet. Fyra år anses vara en tillräckligt lång period för att utveckla ytterligare användningsområden för de berörda verksamma ämnena. De provisoriska gränsvärdena bör därefter bli permanenta.
(7) Bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG bör därför ändras.
(8) Kommissionen anmälde utkastet till detta direktiv till Världshandelsorganisationen (WTO), vars synpunkter beaktats vid den slutliga utformningen av direktivet. Möjligheten att för import fastställa gränsvärden för bekämpningsmedelsrester för vissa särskilda kombinationer av bekämpningsmedel och grödor kommer att undersökas av kommissionen, förutsatt att relevanta data lämnas in.
(9) Detta direktiv är förenligt med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande gränsvärde för bekämpningsmedelsrester skall läggas till i del A i bilaga II till direktiv 86/362/EEG:
">Plats för tabell>"
Artikel 2
Följande gränsvärden för bekämpningsmedelsrester skall läggas till i del B i bilaga II till direktiv 86/363/EEG:
">Plats för tabell>"
Artikel 3
Gränsvärdena för bekämpningsmedelsrester av de berörda verksamma ämnena i bilagan till detta direktiv skall läggas till i bilaga II till direktiv 90/642/EEG.
Artikel 4
Medlemsstaterna skall senast den 30 juni 2003 sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv. De skall omedelbart underrätta kommissionen om detta.
De skall tillämpa dessa bestämmelser från och med den 1 juli 2003.
När en medlemsstat antar dessa bestämmelser, skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 5
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 6
Detta beslut riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 204/2002
av den 19 december 2001
om ändring av rådets förordning (EEG) nr 3696/93 om den statistiska indelningen av produkter efter näringsgren (CPA) inom Europeiska ekonomiska gemenskapen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3696/93 av den 29 oktober 1993 om den statistiska indelningen av produkter efter näringsgren (CPA) inom Europeiska ekonomiska gemenskapen(1), ändrad genom kommissionens förordning (EG) nr 1232/98(2), särskilt artikel 5 b och artikel 6 i denna, och
av följande skäl:
(1) I förordning (EEG) nr 3696/93 fastställs en statistisk indelning av produkter efter näringsgren, nedan kallad CPA, för att tillgodose behovet av statistik inom gemenskapen.
(2) Med anledning av uppdateringen av den statistiska näringsgrensindelningen i gemenskapen (vanligen kallad NACE Rev. 1) är det nödvändigt att göra ändringar i CPA.
(3) Med anledning av revideringen av Harmoniserade systemet och Kombinerade nomenklaturen (HS/KN) enligt kommissionens förordning (EG) nr 2031/2001 av den 6 augusti 2001 om ändring av bilaga I till rådets förordning (EEG) nr 2658/87 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(3) är det nödvändigt att göra ändringar i CPA samt att anpassa och förtydliga texterna.
(4) Det är nödvändigt att ändra CPA, behålla det internationellt integrerade systemet och skapa konvergens globalt.
(5) Förordning (EEG) nr 3696/93 bör därför ändras.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för det statistiska programmet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (EEG) nr 3696/93 skall ersättas med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 315/2002
av den 20 februari 2002
om notering av priserna för färska och kylda slaktkroppar av får på gemenskapens representativa marknader
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2529/2001 av den 19 december 2001 om den gemensamma organisationen av marknaden för får- och getkött(1), särskilt artiklarna 20 och 24 i denna, och
av följande skäl:
(1) Genom förordning (EG) nr 2529/2001 införs ett nytt bidragssystem som ersätter det system som infördes genom rådets förordning (EG) nr 2467/98 av den 3 november 1998 om den gemensamma organisationen av marknaden för får- och getkött(2), ändrad genom förordning (EG) nr 1669/2000(3). För att ta hänsyn till de nya förfarandena och av tydlighetsskäl är det nödvändigt att införa nya regler som ersätter reglerna i kommissionens förordning (EEG) nr 1481/86 av den 15 maj 1986 om fastställande av priser på färska eller kylda slaktkroppar av lamm på gemenskapens representativa marknader och om registrering av priserna på vissa andra slaktkroppskvaliteter för får inom gemenskapen(4), senast ändrad genom förordning (EG) nr 2877/2000(5).
(2) Enligt artikel 20 i förordning (EG) nr 2529/2001 skall medlemsstaterna registrera priserna på får och fårkött. Närmare bestämmelser för prisrapporteringen bör fastställas.
(3) Priset skall vara det som noteras på den eller de representativa marknaderna i varje medlemsstat för de olika kategorierna av färska eller kylda slaktkroppar av får. I de medlemsstater som har mer än en representativ marknad bör det aritmetiska eller, om nödvändigt, det viktade genomsnittet av de priser som har noterats på dessa marknader användas.
(4) Det pris som noterats på marknaden skall grunda sig på priser på slaktkroppar exklusive mervärdeskatt men utan avdrag för andra pålagor. Marknadspriset skall noteras med avseende på "slaktkroppsvikten" enligt definitionen i kommissionens beslut 94/434/EG av den 30 maj 1994 om tillämpningsföreskrifter för rådets direktiv 93/25/EEG vad avser statistiska undersökningar av får- och getbestånd och får- och getproduktion(6), senast ändrad genom beslut 1999/47/EG(7). En avvikelse från denna definition bör dock tillåtas för slaktkroppar av unga lamm som väger mellan 9 och 16 kg av hänsyn till marknadspraxis som ger ett högre handelsvärde åt hela slaktkroppar med huvud och slaktbiprodukter.
(5) I vissa medlemsstater grundar sig dessa priser på priserna för levande djur. I de fallen bör priserna räknas om med hjälp av lämpliga koefficienter. I de områden där det görs en individuell värdering av levande djur för att uppskatta den slaktade vikten, kan dock omräkningen baseras på denna värdering.
(6) För att förklara de grunder på vilka medlemsstaterna genererar priserna skall de lämna uppgifter till kommissionen om den valda representativa marknaden och kategorierna av slaktkroppar samt vikten eller den relativa betydelsen av de uppgifter som används för att beräkna priserna.
(7) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för får och getter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Medlemsstater vars fårköttproduktion överstiger 200 ton per år skall senast varje torsdag meddela kommission priserna på färska eller kylda slaktkroppar av lamm och tackor.
2. Priserna skall vara de som noterats i de prisnoteringsområden som avses i artikel 12 i förordning (EG) nr 2529/2001 av medlemsstater som uppfyller kraven som infördes genom punkt 1. De skall vara grossistpriser som noteras av dessa medlemsstater på den eller de representativa marknaderna under den vecka som föregår den vecka då uppgifterna lämnas. Den eller de representativa marknaderna skall beslutas av medlemsstaterna som nämns ovan. Prisberäkningen skall grunda sig på marknadspriserna exklusive mervärdeskatt.
Artikel 2
1. Marknadspriserna skall noteras med avseende på "slaktvikt" enligt definitionen i beslut 94/434/EG.
Då priset är noterat enligt olika kategorier av slaktkroppar skall priset på den representativa marknaden vara lika med genomsnittet, viktat med koefficienter som har fastställts av medlemstaten för att avspegla den relativa betydelsen av varje kategori, av de priser som har noterats för dessa kategorier under en period på sju dagar i grossistled.
2. Priserna på slaktkroppar av lamm som väger mellan 9 och 16 kg kan dock noteras före borttagande av slaktbiprodukter och huvud i överensstämmelse med normal handelspraxis.
När priserna noteras på grundval av priserna för levande djur skall priset per kg levande vikt divideras med en omräkningskoefficient på högst 0,5. Om det är allmän praxis att sälja slaktkroppen med huvud och slaktbiprodukter kan medlemsstaten fastställa en högre koefficient för lamm med en levande vikt upp till 28 kg.
I de områden där priserna noteras på grundval av en individuell uppskattning av vikten på slaktkroppen av lammet skall omräkningen grundas på denna värdering.
Artikel 3
1. När det förekommer marknader mer än en gång under den period på sju dagar som anges i artikel 2.1 skall priset på varje kategori vara det aritmetiska genomsnittet av de priser som har noterats vid varje marknadstillfälle.
2. Priset i medlemsstaten skall vara genomsnittet av de priser som noteras på de aktuella marknaderna, viktat med koefficienter som avspeglar den relativa betydelsen av varje marknad eller av varje kategori.
3. Om det inte finns någon tillgänglig information skall dock priserna på medlemsstatens representativa marknader fastställas med hjälp särskilt av de senast noterade priserna.
Artikel 4
Senast den 1 mars år 2002 skall medlemsstaterna meddela kommissionen:
a) Varje prisnoteringsområdes representativa marknader.
b) Kategorierna av slaktkroppar av lamm.
c) De koefficienter för viktning och omräkning som avses i artiklarna 2 och 3.
Medlemsstaterna skall underrätta kommissionen om eventuella ändringar i förfarandena senast en månad efter det att ändringarna gjorts.
Artikel 5
Förordning (EEG) nr 1481/86 upphör att gälla.
Artikel 6
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 538/2002
av den 25 mars 2002
om komplettering av bilagan till förordning (EG) nr 2400/96 om upptagandet av vissa namn i "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar" som föreskrivs i rådets förordning (EEG) nr 2081/92 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel(1), senast ändrad genom kommissionens förordning (EG) nr 2796/2000(2), särskilt artikel 6.3 och 6.4 i denna, och
av följande skäl:
(1) Grekland har i enlighet med artikel 5 i förordning (EEG) nr 2081/92 till kommissionen översänt en ansökan om registrering av "Πατατα Κατω Νευροκοπιου" (Patata Kato Nevrokopiou) som geografisk beteckning.
(2) Det har i enlighet med artikel 6.1 i nämnda förordning konstaterats att ansökan är förenlig med den förordningen, särskilt eftersom den omfattar alla komponenter som avses i artikel 4.
(3) Inga invändningar enligt artikel 7 i förordning (EEG) nr 2081/92 har framställts till kommissionen till följd av offentliggörandet i Europeiska gemenskapernas officiella tidning(3) av det produktnamn som anges i bilagan till den här förordningen.
(4) Detta produktnamn kan därför tas upp i "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar" och därmed vara skyddat inom gemenskapen såsom skyddad geografisk beteckning.
(5) Bilagan till denna förordning kompletterar bilagan till kommissionens förordning (EG) nr 2400/96(4) senast ändrad genom förordning (EG) nr 245/2002(5).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (EG) nr 2400/96 skall kompletteras med det produktnamn som anges i bilagan till denna förordning och detta namn skall tas upp i "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar" såsom skyddad geografisk beteckning (SGB) i enlighet med artikel 6.3 i förordning (EEG) nr 2081/92.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 780/2002
av den 8 maj 2002
om ändring av förordning (EG) nr 3063/93 om tillämpningsföreskrifter för rådets förordning (EEG) nr 2019/93 angående stödordningen för produktion av kvalitetshonung
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2019/93 av den 19 juli 1993 om införandet av särskilda bestämmelser för de mindre Egeiska öarna rörande vissa jordbruksprodukter(1), senast ändrad genom förordning (EG) nr 442/2002(2), särskilt artikel 12.3 i denna, och
av följande skäl:
(1) Genom förordning (EEG) nr 2019/93 inrättades för de mindre Egeiska öarna en ordning med stöd för bikupor med produktion av kvalitetshonung. Eftersom artikel 12 i förordningen i dess ändrade lydelse enligt förordning (EG) nr 442/2002 numera hänvisar till "sammanslutningar av producenter" bör följaktligen terminologin i kommissionens förordning (EG) nr 3063/93(3) anpassas.
(2) I syfte att aktualisera förordning (EG) nr 3063/93 bör de undantag för år 1993 strykas som berör sista ansökningsdag, sista utbetalningsdag för stöd och sista datum för inlämnande av uppgifter till kommissionen om utbetalade stöd och andelen stödansökningar som omfattas av kontroll på plats. Dessutom bör hänvisningen till jordbruksomräkningskursen strykas.
(3) Förordning (EG) nr 3063/93 bör därför ändras.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fjäderfäkött och ägg.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. I artikel 2.2 skall den första meningen ersättas med följande: "Sammanslutningarna av biodlare skall förelägga den behöriga myndigheten sina program för godkännande.".
3. Artikel 3 skall ändras på följande sätt:
a) I punkt 1 skall andra stycket utgå.
b) I punkt 2 skall första strecksatsen ersättas med följande: "- Sammanslutningarnas eller biodlarens namn och adress,".
4. I artikel 4 skall andra stycket utgå.
5. Artikel 5 skall ändras på följande sätt:
a) I första stycket skall första och andra strecksatserna ersättas med följande: "- Antal sammanslutningar av biodlare och antal enskilda biodlare som inkommit med stödansökningar.
- Antal bikupor för vilka sammanslutningar av biodlare eller enskilda biodlare ansökt om och beviljats stöd."
b) Det andra stycket utgå.
6. I artikel 6.2 första stycket skall andra meningen utgå.
7. Artikel 8 skall utgå.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets förordning (EG) nr 1460/2002
av den 27 juni 2002
om inrättande av en europeisk sjösäkerhetsbyrå
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
med beaktande av Regionkommitténs yttrande(3),
i enlighet med det förfarande som anges i artikel 251 i fördraget(4), och
av följande skäl:
(1) Ett stort antal lagstiftningsåtgärder har antagits inom gemenskapen för att förbättra säkerheten och förhindra förorening i samband med sjötransporter. För att vara effektiv måste sådan lagstiftning tillämpas korrekt och enhetligt i hela gemenskapen. På så sätt säkerställs likvärdiga konkurrens- och marknadsvillkor, minskas den snedvridning av konkurrensen som följer av de ekonomiska fördelar som fartyg som inte uppfyller normerna åtnjuter och gynnas de rederier och andra som bedriver sjöfartsverksamhet på ett seriöst sätt.
(2) Vissa av de arbetsuppgifter som nu utförs på gemenskapsnivå eller nationell nivå skulle kunna utföras av ett specialiserat expertorgan. Det behövs tekniskt och vetenskapligt stöd och en fast engagerad sakkunskap på hög nivå för att gemenskapens lagstiftning på områdena för sjösäkerhet och förhindrande av förorening från fartyg skall tillämpas korrekt och för att tillämpningen av lagstiftningen skall kunna bevakas och befintliga åtgärders effektivitet utvärderas. Det finns därför ett behov av att inrätta en europeisk sjösäkerhetsbyrå (byrån) inom gemenskapens befintliga institutionsstruktur och befogenhetsfördelning.
(3) Byrån bör allmänt sett fungera som ett tekniskt organ, som gör det möjligt för gemenskapen att agera effektivt för att förbättra bestämmelserna om den övergripande sjösäkerheten och förhindrandet av förorening från fartyg. Byrån bör bistå kommissionen i det fortgående arbetet med att uppdatera och utveckla gemenskapens lagstiftning när det gäller området för sjösäkerhet och förhindrande av förorening från fartyg och tillhandahålla det stöd som behövs för att se till att lagstiftningen tillämpas enhetligt och effektivt i hela gemenskapen genom att bistå kommissionen i utförandet av de uppgifter som den tilldelats genom nuvarande och framtida gemenskapslagstiftning om sjösäkerhet och förhindrande av förorening från fartyg.
(4) För att målsättningarna med byråns inrättande skall uppnås bör byrån utföra ett antal andra viktiga arbetsuppgifter avsedda att höja sjösäkerheten och förhindra förorening från fartyg i de vatten som tillhör medlemsstaterna. I detta avseende bör byrån i samarbete med medlemsstaterna anordna lämplig utbildningsverksamhet beträffande frågor som gäller hamnstatskontroll och flaggstat och tillhandahålla tekniskt stöd i samband med genomförandet av gemenskapslagstiftningen. Den bör underlätta samarbete mellan medlemsstaterna och kommissionen enligt Europaparlamentets och rådets direktiv 2002/59/EG av den 27 juni 2002 om inrättandet av ett övervaknings- och informationssystem för sjötrafik i gemenskapen och om upphävande av rådets direktiv 93/75/EEG(5) genom att utveckla och sköta det informationssystem som behövs dels för att uppnå de mål som uppställs i direktivet, dels i verksamhet som gäller utredningar av allvarliga olyckor till sjöss. Den bör ge kommissionen och medlemsstaterna objektiva, tillförlitliga och jämförbara uppgifter och data om sjösäkerhet och förhindrande av förorening från fartyg, så att dessa kan vidta nödvändiga åtgärder för att förbättra befintliga åtgärder och utvärdera åtgärdernas effektivitet. Den bör se till att den kunskap om sjösäkerhet som finns inom gemenskapen står till förfogande för de stater som ansöker om anslutning. Dessa stater och andra tredjeländer som ingått avtal med Europeiska gemenskapen, genom vilka de antar och genomför gemenskapslagstiftningen inom området för sjösäkerhet och förhindrande av förorening från fartyg, bör ha möjlighet att delta i byråns verksamhet.
(5) Byrån bör arbeta för att förbättra samarbetet mellan medlemsstaterna och utarbeta bra metoder och sprida kunskap om dessa i gemenskapen. Detta bör i sin tur leda till att sjösäkerhetssystemet i gemenskapen blir bättre och att risken för olyckor, förorening och dödsfall till sjöss minskar.
(6) För att byrån skall kunna utföra sina arbetsuppgifter på vederbörligt sätt, bör dess tjänstemän besöka medlemsstaterna för att kontrollera att gemenskapens system för sjösäkerhet och förhindrande av förorening från fartyg fungerar. Besöken bör genomföras i enlighet med en praxis som byråns styrelse fastställer, och de bör underlättas av medlemsstaternas myndigheter.
(7) Byrån bör tillämpa den relevanta gemenskapslagstiftningen rörande allmänhetens tillgång till handlingar och skydd för enskilda vid databehandling av personuppgifter. Den bör ge allmänheten och alla berörda parter objektiv, tillförlitlig och lättbegriplig information om sin verksamhet.
(8) När det gäller byråns avtalsrättsliga ansvar, som regleras av den lagstiftning som är tillämplig på det avtal som byrån ingått, bör domstolen vara behörig att träffa avgöranden med stöd av en skiljedomsklausul i avtalet. Domstolen skall också vara behörig i tvister som gäller byråns utomobligatoriska ersättningsansvar.
(9) För att effektivt kunna se till att byrån fullgör sina uppgifter bör medlemsstaterna och kommissionen vara företrädda i en styrelse som har de befogenheter som är nödvändiga för att fastställa budgeten och kontrollera att den genomförs, anta lämpliga finansiella bestämmelser, utarbeta tydliga förfaranden för byråns beslutsfattande, godkänna dess arbetsprogram, behandla ansökningar från medlemsstater om tekniskt bistånd, fastställa riktlinjer för besök i medlemsstaterna samt utnämna den verkställande direktören. Med tanke på denna särskilda byrås synnerligen tekniska och vetenskapliga uppdrag och uppgifter bör styrelsen bestå av en företrädare för varje medlemsstat och fyra företrädare för kommissionen som är ledamöter med en hög nivå av sakkunskap. För att ytterligare säkerställa högsta möjliga nivå när det gäller sakkunskap och erfarenhet i styrelsen och för att de mest berörda branschsektorerna skall kunna delta aktivt i byråns verksamhet, bör kommissionen utnämna oberoende yrkesverksamma personer inom dessa sektorer som ledamöter i styrelsen, utan rösträtt, på grundval av personliga meriter och personlig erfarenhet inom området för sjösäkerhet och förhindrande av förorening från fartyg och inte som företrädare för särskilda branschorganisationer.
(10) För att byrån skall fungera väl måste den verkställande direktören vara utsedd på grundval av meriter och dokumenterad skicklighet i förvaltning och ledarskap samt kompetens och erfarenheter som är relevanta för sjösäkerhet och förhindrande av förorening från fartyg och han/hon måste vid utförandet av sina arbetsuppgifter vara helt oavhängig och flexibel när det gäller byråns inre organisation. Den verkställande direktören bör därför förbereda och vidta alla åtgärder som är nödvändiga för att se till att byråns arbetsprogram genomförs, varje år utarbeta ett utkast till allmän rapport och lägga fram det för styrelsen, göra beräkningar av byråns intäkter och utgifter samt genomföra budgeten.
(11) För att garantera byråns fullständiga oberoende och självständighet anses det nödvändigt att den har en egen budget, där intäkterna främst utgörs av ett bidrag från gemenskapen.
(12) I takt med att allt fler decentraliserade organ har inrättats på senare år har budgetmyndigheten de gångna åren försökt förbättra insynen i och kontrollen av förvaltningen av gemenskapsanslagen till organen, särskilt när det gäller budgetering av avgifter, finansiell kontroll, befogenheter att bevilja ansvarsfrihet, avsättning till pensionssystemet samt det interna budgetförfarandet (uppförandekodex). På liknande sätt bör Europaparlamentets och rådets förordning (EG) nr 1073/1999 av den 25 maj 1999 om utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF)(6) oinskränkt tillämpas när det gäller byrån, som bör ansluta sig till det interinstitutionella avtalet av den 25 maj 1999 mellan Europaparlamentet, Europeiska unionens råd och Europeiska gemenskapernas kommission om interna utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF)(7).
(13) Senast fem år från det att byrån inlett sin verksamhet bör styrelsen beställa en oberoende extern utvärdering för att bedöma i vilken utsträckning förordningen, byrån och dess arbetsmetoder bidragit till att etablera en hög sjösäkerhetsnivå och en hög nivå på förhindrandet av förorening från fartyg.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
MÅL OCH UPPGIFTER
Artikel 1
Mål
1. Genom denna förordning inrättas en europeisk sjösäkerhetsbyrå, (byrån), i syfte att skapa en hög, enhetlig och effektiv sjösäkerhetsnivå och en hög nivå på förhindrandet av förorening från fartyg inom gemenskapen.
2. Byrån skall ge medlemsstaterna och kommissionen tekniskt och vetenskapligt stöd och tillhandahålla sakkunskap på hög nivå för att hjälpa dem att på ett korrekt sätt tillämpa gemenskapslagstiftningen på området för sjösäkerhet och förhindrande av förorening från fartyg, att bevaka genomförandet av denna och att utvärdera befintliga åtgärders effektivitet.
Artikel 2
Uppgifter
För att säkerställa att de mål som anges i artikel 1 uppnås på ett lämpligt sätt skall byrån utföra följande uppgifter:
a) Den skall vid behov bistå kommissionen i det förberedande arbetet med att uppdatera och utveckla gemenskapslagstiftningen när det gäller sjösäkerhet och förhindrande av förorening från fartyg, särskilt med beaktande av den internationella lagstiftningens utveckling på området. I denna uppgift ingår att analysera forskningsprojekt som utförs inom området för sjösäkerhet och förhindrande av förorening från fartyg.
b) Den skall bistå kommissionen i arbetet med att effektivt genomföra gemenskapslagstiftningen om sjösäkerhet och förhindrande av förorening från fartyg i hela gemenskapen. Byrån skall särskilt
i) kontrollera att hela gemenskapssystemet för hamnstatskontroll fungerar, eventuellt genom besök i medlemsstaterna, och föreslå kommissionen förbättringar av systemet,
ii) ge kommissionen det tekniska stöd den behöver för att delta i arbetet i de tekniska arbetsgrupper som inrättats inom ramen för det i Paris ingångna samförståndsavtalet om hamnstatskontroll (the Paris Memorandum of Understanding on Port State Control),
iii) bistå kommissionen i genomförandet av de arbetsuppgifter som den har tilldelats av kommissionen genom befintlig och kommande gemenskapslagstiftning om sjösäkerhet och förhindrande av förorening från fartyg, särskilt lagstiftning om klassificeringssällskap, säkerheten på passagerarfartyg, säkerheten för fartygsbesättningar samt sjöfolks utbildning, certifiering och vakthållning.
c) Den skall i samarbete med medlemsstaterna
i) vid behov anordna relevant utbildningsverksamhet på områden som står under hamnstatens och flaggstatens ansvar,
ii) utveckla tekniska lösningar och ge tekniskt stöd avseende genomförandet av gemenskapslagstiftningen.
d) Den skall underlätta samarbetet mellan medlemsstaterna och kommissionen på det område som omfattas av direktiv 2002/59/EG. Den skall särskilt
i) främja samarbete mellan kuststater i de sjöfartsområden som omfattas av det direktivet,
ii) utveckla och sköta de informationssystem som är nödvändiga för att uppnå det direktivets syften.
e) Den skall underlätta samarbetet mellan medlemsstaterna och kommissionen vid utarbetandet, med beaktande av medlemsstaternas olika rättssystem, av en gemensam metod för utredning av sjöolyckor i enlighet med internationellt överenskomna principer, vid tillhandahållande av stöd till medlemsstaterna vid utredning av allvarliga sjöolyckor och vid analys av befintliga olycksrapporter.
f) Byrån skall förse kommissionen och medlemsstaterna med objektiva, tillförlitliga och jämförbara uppgifter och data om sjösäkerhet och förorening från fartyg, så att dessa kan vidta nödvändiga åtgärder för att förbättra sjösäkerheten [och förhindrandet av förorening från fartyg] och utvärdera befintliga åtgärders effektivitet. I dessa uppgifter ingår att samla in, registrera och utvärdera tekniska data om sjösäkerhet, sjöfart och marina föroreningar, oavsiktliga eller avsiktliga, att systematiskt utnyttja och samköra befintliga databaser och att vid behov skapa nya databaser. Byrån skall, på grundval av insamlade data, bistå kommissionen när den var sjätte månad offentliggör uppgifter om fartyg som vägrats tillträde till hamnar i gemenskapen med tillämpning av rådets direktiv 95/21/EG av den 19 juni 1995 om tillämpning av internationella normer för säkerhet på fartyg, förhindrande av förorening samt boende- och arbetsförhållanden ombord på fartyg som anlöper gemenskapens hamnar och framförs i medlemsstaternas territorialvatten (hamnstatskontroll)(8). Byrån skall också bistå kommissionen och medlemsstaterna i deras verksamhet för att förbättra identifiering och lagföring av fartyg som gjort sig skyldiga till olagliga utsläpp.
g) Under förhandlingarna med de stater som ansöker om anslutning får byrån tillhandahålla tekniskt stöd för genomförandet av gemenskapslagstiftningen om sjösäkerhet och förhindrande av förorening från fartyg. Denna uppgift skall samordnas med befintliga regionala samarbetsprogram och vid behov omfatta anordnande av relevant utbildningsverksamhet.
Artikel 3
Besök i medlemsstaterna
1. För att sköta sina uppgifter får byrån genomföra besök i medlemsstaterna i enlighet med de riktlinjer som styrelsen fastställt. Medlemsstaternas nationella myndigheter skall underlätta arbetet för byråns personal.
2. Byrån skall underrätta den berörda medlemsstaten om det planerade besöket, namnen på de bemyndigade tjänstemännen och vilken dag besöket skall inledas. De bemyndigade tjänstemännen skall genomföra besöket efter uppvisande av ett beslut från byråns verkställande direktör, där syftet och målet med besöket anges.
3. Efter varje besök skall byrån upprätta en rapport och skicka den till kommissionen och den berörda medlemsstaten.
Artikel 4
Öppenhet och skydd av information
1. Byrån skall tillämpa principerna i Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar(9), när den behandlar ansökningar om tillgång till de handlingar som den innehar.
2. Byrån får på eget initiativ kommunicera på de områden som ingår i dess uppdrag. Den skall särskilt se till att allmänheten och alla berörda parter snabbt får objektiv, tillförlitlig och lättbegriplig information om dess arbete.
3. Styrelsen skall fastställa de interna regler som är nödvändiga för tillämpningen av punkterna 1 och 2.
4. Den information som kommissionen och byrån samlar in i enlighet med denna förordning skall omfattas av Europaparlamentets och rådets förordning (EG) nr 45/2001 av den 18 december 2000 om skydd för enskilda då gemenskapsinstitutionerna och gemenskapsorganen behandlar personuppgifter och om den fria rörligheten för sådana uppgifter(10).
KAPITEL II
BYRÅNS ORGANISATION OCH VERKSAMHET
Artikel 5
Rättslig status, regionala centrum
1. Byrån skall vara ett gemenskapsorgan. Den skall vara en juridisk person.
2. Byrån skall i varje medlemsstat ha den mest vittgående rättskapacitet som tillerkänns juridiska personer enligt den nationella lagstiftningen. Den skall särskilt kunna förvärva och avyttra lös och fast egendom samt föra talan inför domstolar och andra myndigheter.
3. På begäran från kommissionen och med samtycke från de berörda medlemsstaterna får styrelsen besluta att inrätta de regionala centrum som byrån behöver för att kunna utföra de arbetsuppgifter avseende övervakning av navigation och sjötrafik som anges i direktiv 2002/59/EG.
4. Byrån skall företrädas av den verkställande direktören.
Artikel 6
Personal
1. Tjänsteföreskrifterna för tjänstemän i Europeiska gemenskaperna, anställningsvillkoren för övriga anställda i Europeiska gemenskaperna och bestämmelser som antagits gemensamt av Europeiska gemenskapernas institutioner för tillämpningen av tjänsteföreskrifterna och anställningsvillkoren skall gälla för byråns personal. Styrelsen skall i samförstånd med kommissionen utfärda nödvändiga tillämpningsföreskrifter.
2. Om inte annat föreskrivs i artikel 16, skall byrån, när det gäller dess egen personal, utöva de befogenheter som enligt tjänsteföreskrifterna och anställningsvillkoren för övriga anställda tillkommer tillsättningsmyndigheten.
3. Byråns personal skall bestå av tjänstemän som utsetts eller avdelats temporärt av kommissionen eller medlemsstaterna och av andra anställda som vid behov skall anställas av byrån för att fullgöra dess uppgifter.
Artikel 7
Privilegier och immunitet
Byrån och dess personal skall omfattas av protokollet om Europeiska gemenskapernas immunitet och privilegier.
Artikel 8
Ansvar
1. Byråns avtalsrättsliga ansvar skall regleras av den lagstiftning som är tillämplig på avtalet i fråga.
2. Domstolen skall vara behörig att träffa avgöranden på grundval av skiljedomsklausuler i de avtal som ingåtts av byrån.
3. Vad beträffar utomobligatoriskt ansvar skall byrån, i enlighet med de allmänna principer som är gemensamma för medlemsstaternas rättsordningar, ersätta skada som orsakats av dess enheter eller av dess anställda under tjänsteutövning.
4. Domstolen skall vara behörig att avgöra tvister om sådant skadestånd som avses i punkt 3.
5. De anställdas personliga ansvar gentemot byrån skall regleras av bestämmelserna i de tjänsteföreskrifter eller de anställningsvillkor som gäller för dem.
Artikel 9
Språk
1. Bestämmelserna i förordning nr 1 av den 15 april 1958 om vilka språk som skall användas i Europeiska ekonomiska gemenskapen(11) skall gälla för byrån.
2. De översättningar som krävs för byråns arbete skall utföras av Översättningscentrum för Europeiska unionens organ.
Artikel 10
Styrelsens inrättande och dess befogenheter
1. En styrelse inrättas härmed för byrån.
2. Styrelsen skall
a) utnämna den verkställande direktören i enlighet med artikel 16,
b) senast den 30 april varje år anta byråns allmänna rapport för föregående år och skicka den till medlemsstaterna, Europaparlamentet, rådet och kommissionen,
c) inom ramen för utarbetandet av arbetsprogrammet behandla ansökningar från medlemsstater om tekniskt stöd enligt artikel 2 c ii,
d) senast den 31 oktober varje år, efter att ha beaktat kommissionens yttrande, anta byråns arbetsprogram för det kommande året och skicka det till medlemsstaterna, Europaparlamentet, rådet och kommissionen.
Detta arbetsprogram skall antas utan att det påverkar gemenskapens årliga budgetförfarande. Om kommissionen inom 15 dagar från den tidpunkt då arbetsprogrammet antagits meddelar att den inte samtycker till det antagna arbetsprogrammet, skall styrelsen behandla det igen och inom två månader, vid den andra behandlingen, anta det eventuellt ändrade arbetsprogrammet, antingen med två tredjedels majoritet, inbegripet kommissionens företrädare, eller med enhällighet bland medlemsstaternas företrädare,
e) anta byråns slutliga budget innan räkenskapsåret börjar och vid behov anpassa den till gemenskapens bidrag och byråns övriga intäkter,
f) utarbeta förfaranden för de beslut som skall fattas av den verkställande direktören,
g) fastställa riktlinjer för de besök som skall genomföras enligt artikel 3,
h) utföra de av sina åligganden som hör samman med byråns budget i enlighet med artiklarna 18, 19 och 21,
i) ha disciplinär bestämmanderätt över den verkställande direktören och de enhetschefer som avses i artikel 15.3,
j) fastställa sin arbetsordning.
Artikel 11
Styrelsens sammansättning
1. Styrelsen skall bestå av en företrädare för varje medlemsstat och fyra företrädare för kommissionen samt av fyra yrkesverksamma personer som kommissionen utsett inom de mest berörda sektorerna, vilka personer inte skall ha rösträtt.
Styrelseledamöter skall utses på grundval av relevant erfarenhet och sakkunskap inom området för sjösäkerhet och förhindrande av förorening från fartyg.
2. Varje medlemsstat och kommissionen skall utse sina företrädare i styrelsen samt en suppleant, som skall företräda ledamoten i dennes frånvaro.
3. Mandatperioden skall vara fem år. Mandatet kan förnyas en gång.
4. I förekommande fall skall deltagande av företrädare för tredje land och villkoren för detta fastställas genom de förfaranden som avses i artikel 17.2.
Artikel 12
Styrelsens ordförande
1. Styrelsen skall utse en ordförande och en vice ordförande bland sina ledamöter. Vice ordföranden skall automatiskt ersätta ordföranden om denne är förhindrad att fullgöra sina åligganden.
2. Mandatperioden för ordföranden och vice ordföranden skall vara tre år och skall upphöra om uppdraget som styrelseledamot upphör. Mandatet skall kunna förnyas en gång.
Artikel 13
Sammanträden
1. Styrelsens ordförande skall sammankalla till styrelsens sammanträden.
2. Byråns verkställande direktör skall delta i överläggningarna.
3. Styrelsen skall hålla två ordinarie sammanträden per år. Den skall dessutom sammanträda på initiativ av ordföranden eller på begäran av kommissionen eller en tredjedel av medlemsstaterna.
4. Styrelsen får, om det är fråga om konfidentiella uppgifter eller intressekonflikter, besluta att ta upp särskilda frågor på sin dagordning utan närvaro av de ledamöter som har utsetts i sin egenskap av yrkesverksamma personer från de mest berörda sektorerna. Närmare regler för tillämpningen av denna bestämmelse får fastställas i arbetsordningen.
5. Styrelsen får bjuda in alla personer vars åsikter kan vara av intresse att delta som observatörer vid sammanträdena.
6. Styrelseledamöterna får, med förbehåll för bestämmelserna i arbetsordningen, biträdas av rådgivare eller experter.
7. Styrelsens sekretariat skall tillhandahållas av byrån.
Artikel 14
Röstning
1. Styrelsen skall fatta sina beslut med två tredjedelars majoritet av alla ledamöter som har rösträtt.
2. Varje ledamot skall ha en röst. Den verkställande direktören får inte rösta.
I en ledamots frånvaro skall suppleanten ha rätt att utöva dennes rösträtt.
3. Röstningsförfarandena skall fastställas utförligare i arbetsordningen, särskilt villkoren för en ledamot att agera på en annan ledamots vägnar.
Artikel 15
Den verkställande direktörens arbetsuppgifter och befogenheter
1. Byrån skall ledas av den verkställande direktören, som skall vara fullständigt oavhängig i sin tjänsteutövning, utan att det påverkar kommissionens och styrelsens respektive befogenheter.
2. Den verkställande direktören skall ha följande arbetsuppgifter och befogenheter:
a) Han/hon skall utarbeta arbetsprogrammet och lägga fram det för styrelsen efter samråd med kommissionen. Han/hon skall vidta nödvändiga åtgärder för att genomföra programmet. Han/hon skall besvara alla ansökningar om stöd från någon medlemsstat i enlighet med artikel 10.2 c eller från kommissionen.
b) Han/hon skall efter att ha hört kommissionen besluta om genomförandet av sådana besök som avses i artikel 3, i enlighet med de riktlinjer som fastställts av styrelsen i enlighet med artikel 10.2 g.
c) Han/hon skall vidta nödvändiga åtgärder för att se till att byrån fungerar i enlighet med bestämmelserna i denna förordning, bl.a. genom att anta anvisningar för den interna administrationen och offentliggöra meddelanden.
d) Han/hon skall organisera ett effektivt övervakningssystem för att kunna jämföra byråns resultat med verksamhetens mål. På grundval därav skall den verkställande direktören varje år utarbeta ett utkast till allmän rapport och lägga fram det för styrelsen. Han/hon skall fastställa förfaranden för regelbunden utvärdering baserade på erkända branschnormer.
e) Han/hon skall utöva de befogenheter i förhållande till personalen som anges i artikel 6.2.
f) Han/hon skall göra beräkningar av byråns intäkter och utgifter i enlighet med artikel 18 och genomföra budgeten i enlighet med artikel 19.
3. Den verkställande direktören får biträdas av en eller flera enhetschefer. Om den verkställande direktören är frånvarande eller har förhinder, skall han/hon ersättas av någon av enhetscheferna.
Artikel 16
Utnämning av verkställande direktör
1. Byråns verkställande direktör skall utnämnas av styrelsen på grundval av meriter, dokumenterad skicklighet i förvaltning och ledarskap samt kompetens och erfarenheter som är relevanta för sjösäkerhet och förhindrande av förorening från fartyg. Styrelsen skall fatta sitt beslut med fyra femtedels majoritet av alla ledamöter som har rösträtt. Kommissionen får föreslå en eller flera kandidater.
Den verkställande direktören kan avsättas av styrelsen enligt samma förfarande.
2. Den verkställande direktörens mandatperiod skall vara fem år. Mandatet får förnyas en gång.
Artikel 17
Tredje lands deltagande
1. Tredjeländer får delta i byråns arbete, om de genom avtal med Europeiska gemenskapen har antagit och tillämpar gemenskapslagstiftningen inom området för sjösäkerhet och förhindrande av förorening från fartyg.
2. Inom ramen för dessa avtal skall förfaranden utarbetas genom vilka bl.a. skall fastställas karaktären och omfattningen av de detaljerade bestämmelserna för dessa länders deltagande i byråns arbete, inbegripet bestämmelser om ekonomiska bidrag och personal.
KAPITEL III
FINANSIELLA KRAV
Artikel 18
Budget
1. Byråns intäkter skall bestå av
a) bidrag från gemenskapen,
b) eventuella bidrag från de tredjeländer som deltar i byråns arbete i enlighet med artikel 17,
c) avgifter för publikationer, utbildning och/eller andra tjänster som byrån tillhandahåller.
2. Byråns utgifter skall omfatta kostnader för personal, administration, infrastruktur och drift.
3. Den verkställande direktören skall göra en beräkning av byråns intäkter och utgifter för påföljande budgetår och överlämna denna till styrelsen tillsammans med en tjänsteförteckning.
4. Intäkter och utgifter skall balansera varandra.
5. Styrelsen skall senast den 30 april varje år anta ett budgetförslag, tillsammans med ett preliminärt arbetsprogram, och överlämna det till kommissionen och de tredjeländer som deltar i byråns arbete i enlighet med artikel 17.
På grundval av detta budgetförslag skall kommissionen fastställa motsvarande beräkningar i det preliminära förslag till Europeiska unionens allmänna budget som den skall förelägga rådet enligt artikel 272 i fördraget. Ramarna för gemenskapens godkända budgetprognos för de kommande åren måste iakttas.
6. När budgetmyndigheten har antagit Europeiska unionens allmänna budget, skall styrelsen anta byråns budget och slutliga arbetsprogram och vid behov anpassa dem till gemenskapens bidrag. Den skall utan dröjsmål överlämna dem till kommissionen, budgetmyndigheten och de tredjeländer som deltar i byråns arbete.
Artikel 19
Genomförande och kontroll av budgeten
1. Den verkställande direktören skall genomföra byråns budget.
2. Kontroll av byråns åtaganden, betalningar av alla utgifter samt kontroll av alla intäkters existens och inkassering av alla intäkter skall utföras av kommissionens styrekonom.
3. Den verkställande direktören skall senast den 31 mars varje år översända utförliga räkenskaper över intäkter och utgifter under föregående räkenskapsår till kommissionen, styrelsen och revisionsrätten.
Revisionsrätten skall granska räkenskaperna i enlighet med artikel 248 i fördraget. Den skall årligen offentliggöra en rapport om byråns verksamhet.
4. Europaparlamentet skall på styrelsens rekommendation bevilja byråns verkställande direktör ansvarsfrihet för genomförandet av budgeten.
Artikel 20
Bekämpning av bedrägeri
1. För bekämpning av bedrägeri, korruption och annan olaglig verksamhet skall bestämmelserna i Europaparlamentets och rådets förordning (EG) nr 1073/1999 tillämpas utan begränsning när det gäller byrån.
2. Byrån skall ansluta sig till det interinstitutionella avtalet av den 25 maj 1999 om interna utredningar som utförs av OLAF och skall utan dröjsmål utfärda lämpliga föreskrifter, som skall gälla all dess personal.
3. I beslut om finansiering samt i de avtal om och instrument för genomförande som ingåtts till följd av dessa beslut skall det uttryckligen föreskrivas att revisionsrätten och OLAF vid behov skall få utföra kontroller på plats hos dem som mottagit anslag från byrån och hos de ombud som fördelat dessa anslag.
Artikel 21
Finansiella bestämmelser
Styrelsen skall, efter att ha mottagit kommissionens godkännande och revisionsrättens yttrande, anta byråns budgetförordning. I denna budgetförordning skall det särskilt anges vilket förfarande som skall användas vid utarbetandet och genomförandet av byråns budget i enlighet med artikel 142 i budgetförordningen av den 21 december 1977 för Europeiska gemenskapernas allmänna budget(12).
KAPITEL IV
SLUTBESTÄMMELSER
Artikel 22
Utvärdering
1. Senast fem år efter det att byrån inlett sin verksamhet skall styrelsen beställa en oberoende extern utvärdering av förordningens tillämpning. Kommissionen skall tillhandahålla byrån all den information som denna anser sig behöva för att kunna genomföra denna utvärdering.
2. I utvärderingen skall det bedömas i vilken utsträckning förordningen, byrån och dess arbetsmetoder bidragit till att etablera en hög sjösäkerhetsnivå och en hög nivå på förhindrandet av förorening från fartyg. Styrelsen skall utarbeta särskilda riktlinjer i samförstånd med kommissionen och efter samråd med de berörda parterna.
3. Styrelsen skall ta emot utvärderingen och utfärda rekommendationer till kommissionen om hur förordningen, byrån och dess arbetsmetoder eventuellt bör ändras. Utvärderingsresultatet och rekommendationerna skall överlämnas av kommissionen till Europaparlamentet och rådet samt offentliggöras.
Artikel 23
Inledande av byråns verksamhet
Byrån skall vara verksam senast tolv månader efter det att förordningen trätt i kraft.
Artikel 24
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Europaparlamentets och rådets förordning (EG) nr 1774/2002
av den 3 oktober 2002
om hälsobestämmelser för animaliska biprodukter som inte är avsedda att användas som livsmedel
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 152.4 b i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
enligt förfarandet i artikel 251 i fördraget(3), mot bakgrund av det gemensamma utkast som förlikningskommittén godkände den 12 september 2002, och
av följande skäl:
(1) I rådets direktiv 90/667/EEG av den 27 november 1990 om fastställande av veterinära bestämmelser om bortskaffande och bearbetning av animaliskt avfall och dess utsläppande på marknaden samt om förhindrande av sjukdomsalstrande organismer i foder av animaliskt ursprung samt om ändring av direktiv 90/425/EEG(4) fastställs principen att alla typer av animaliskt avfall, oavsett källa, efter lämplig behandling får användas för produktion av foderråvaror.
(2) Den vetenskapliga styrkommittén har antagit flera yttranden i denna fråga sedan det direktivet antogs. Den viktigaste slutsatsen i dessa är att animaliska biprodukter från djur som vid en hälsobesiktning inte bedöms vara lämpliga för användning som livsmedel inte heller bör få komma in i näringskedjan för djur.
(3) Mot bakgrund av dessa vetenskapliga yttranden bör det göras skillnad mellan de åtgärder som skall vidtas beroende på vilken typ av animaliska biprodukter som används. De möjliga användningsområdena för vissa animalieprodukter bör begränsas. Regler bör fastställas för annan användning av animaliska biprodukter än i foder och för bortskaffandet av dessa.
(4) Mot bakgrund av de senaste årens erfarenheter är det lämpligt att klargöra förhållandet mellan direktiv 90/667/EEG och gemenskapens miljölagstiftning. Denna förordning bör inte påverka tillämpningen av gällande miljölagstiftning eller förhindra utarbetandet av nya regler om miljöskydd, särskilt inte när det gäller biologiskt nedbrytbart avfall. I detta avseende har kommissionen åtagit sig att i slutet av 2004 utarbeta ett direktiv om bioavfall, inklusive matavfall, och vars syfte kommer att vara dels att fastställa bestämmelser om användning, återvinning, återanvändning och omhändertagande av detta avfall, dels att kontrollera eventuella föroreningar.
(5) Genom den internationella vetenskapliga konferens om kött- och benmjöl som kommissionen och Europaparlamentet arrangerade i Bryssel den 1-2 juli 1997, inleddes en debatt om produktionen av kött- och benmjöl och om dess användning som foder. Det framhölls vid denna konferens att den framtida politiken på området behövde diskuteras ytterligare. För att kunna skapa så bred offentlig debatt som möjligt om gemenskapens framtida foderlagstiftning, färdigställde kommissionen i november 1997 ett samrådsdokument om kött- och benmjöl. Efter detta samråd verkar det råda samsyn kring behovet av att ändra direktiv 90/667/EEG så att dess bestämmelser anpassas till de nya vetenskapliga rönen.
(6) I Europaparlamentets resolution om BSE och säkert djurfoder av den 16 november 2000(5) krävde Europaparlamentet ett förbud mot användning av animaliskt protein i foder fram till dess att denna förordning träder i kraft.
(7) Vetenskapliga utlåtanden pekar på att utfodring av en djurart med protein som härrör från kroppar, eller delar av kroppar, från samma djurart medför risk för spridning av sjukdomar. Som en försiktighetsåtgärd bör sådan utfodring således förbjudas. Genomförandebestämmelser bör antas för att säkerställa nödvändigt avskiljande av animaliska biprodukter avsedda för användning i foder i alla bearbetnings-, lagrings- och transportstadier. Det bör emellertid finnas utrymme för undantag från detta allmänna förbud för fisk och pälsdjur, om vetenskapliga utlåtanden motiverar detta.
(8) Matavfall som innehåller produkter av animaliskt ursprung kan också vara en vektor för sjukdomsspridning. Allt matavfall från transportmedel i internationell trafik bör bortskaffas på ett säkert sätt. Matavfall som produceras inom gemenskapen bör inte användas för utfodring av produktionsdjur, med undantag av pälsdjur.
(9) Sedan oktober 1996 har kontoret för livsmedels- och vetrinärfrågor (FVO) genomfört ett antal inspektioner i medlemsstaterna för att ta reda på vilka de viktigaste riskfaktorerna är och hur dessa hanteras samt hur övervakningen av BSE sker. Bedömningen gällde bland annat systemen för kommersiell konvertering och andra metoder för att hantera animaliskt avfall. Dessa inspektioner har utmynnat i allmänna slutsatser och ett antal rekommendationer, särskilt beträffande möjligheten att spåra animaliska biprodukter.
(10) För att eliminera risken för att patogener och/eller restsubstanser av ämnen sprids bör animaliska biprodukter bearbetas, lagras och hållas avskilda i godkända och övervakade anläggningar som den berörda medlemsstaten utsett, eller bortskaffas på lämpligt sätt. I vissa fall kan en bearbetnings-, förbrännings- eller samförbränningsanläggning som ligger i en annan medlemsstat användas, särskilt när detta är motiverat på grund av avstånd, transporttid eller kapacitetsproblem.
(11) Europaparlamentets och rådets direktiv 2000/76/EG av den 4 december 2000 om förbränning av avfall(6) skall inte tillämpas på förbränningsanläggningar om det avfall som hanteras endast består av slaktkroppar av djur. Det är nödvändigt att fastställa minimikrav för sådana förbränningsanläggningar för att skydda djurs och människors hälsa. I väntan på att gemenskapen skall införa dessa krav får medlemsstaterna anta miljölagar för sådana anläggningar. Mindre strikta krav bör tillämpas på förbränningsanläggningar med låg kapacitet, exempelvis sådana som är belägna på jordbruksföretag och krematorier för sällskapsdjur, eftersom det material som hanteras där utgör en lägre risk och för att undvika onödiga transporter av animaliska biprodukter.
(12) Särskilda bestämmelser bör fastställas om kontroll av bearbetningsanläggningar, särskilt när det gäller detaljförfaranden för validering av bearbetningsmetoder och för egentillsyn av produktionen.
(13) Undantag från reglerna för användning av animaliska biprodukter kan vara lämpliga för att underlätta utfodring av djur som inte är avsedda att användas som livsmedel. De behöriga myndigheterna bör övervaka sådan användning.
(14) Undantag kan även vara lämpliga för att göra det möjligt att bortskaffa animaliska biprodukter på plats under övervakning. Kommissionen bör få den information som behövs för att kunna övervaka situationen och fastställa tillämpningsföreskrifter om så är lämpligt.
(15) För att säkerställa att hälsobestämmelserna genomförs på ett enhetligt sätt bör gemenskapsinspektioner utföras i medlemsstaterna. Sådana inspektioner bör också omfatta kontrollförfaranden.
(16) Gemenskapens hälsolagstiftning bygger på etablerade vetenskapliga rön. De behöriga vetenskapliga kommittéer som inrättats genom kommissionens beslut 97/404/EG(7) och 97/579/EG(8) bör därför alltid vid behov höras. I synnerhet behövs det ytterligare vetenskapliga utlåtanden om användning av produkter av animaliskt ursprung i organiska gödningsmedel och jordförbättringsmedel. I avvaktan på att gemenskapsregler antas mot bakgrund av dessa utlåtanden, får medlemsstaterna behålla eller anta nationella regler som är strängare än de som återfinns i denna förordning om dessa regler överensstämmer med annan tillämplig gemenskapslagstiftning.
(17) Medlemsstaterna använder sig av ett stort antal system för finansiellt stöd för bearbetning, insamling, lagring och bortskaffande av animaliska biprodukter. För att detta inte skall påverka konkurrensvillkoren för jordbruksprodukter, är det nödvändigt att genomföra en undersökning på området och, vid behov, vidta lämpliga åtgärder på gemenskapsnivå.
(18) Mot bakgrund av vad som angetts ovan verkar det vara nödvändigt att göra en genomgripande revidering av de av gemenskapens bestämmelser som gäller animaliska biprodukter.
(19) Animaliska biprodukter som inte är avsedda att användas som livsmedel (särskilt bearbetat animaliskt protein, utsmält fett, sällskapsdjursfoder, hudar, skinn och ull) finns upptagna i produktförteckningen i bilaga I till fördraget. För vissa delar av jordbruksbefolkningen utgör avyttringen av sådana produkter en viktig inkomstkälla. För att säkerställa att denna sektor utvecklas på ett ändamålsenligt sätt och kan öka sin produktion, bör det fastställas hälsobestämmelser för människor och djur för dessa produkter på gemenskapsnivå. Med tanke på att djur lätt smittas av olika sjukdomar bör särskilda krav gälla när animaliska biprodukter släpps ut på marknaden, särskilt i regioner med hög hälsostatus.
(20) För att säkerställa att produkter som importeras från tredje land uppfyller hälsokrav som är minst likvärdiga med eller motsvarande dem som tillämpas i gemenskapen, bör det inrättas ett system för godkännande av tredje länder och anläggningar i dessa, liksom bestämmelser om gemenskapsinspektioner för att se till att villkoren för godkännande efterlevs. Import från tredje land av sällskapsdjursfoder och råvaror för sådant foder får göras på villkor som avviker från dem som gäller samma typer av material som producerats i gemenskapen, särskilt när det gäller de garantier som krävs beträffande restsubstanser som är förbjudna enligt rådets direktiv 96/22/EG av den 29 april 1996 om förbud mot användning av vissa ämnen med hormonell och tyreostatisk verkan samt av B-agonister vid animalieproduktion och om upphävande av direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG(9). För att det skall vara möjligt att garantera att sådant sällskapsdjursfoder och sådana råvaror bara används i avsett syfte är det nödvändigt att fastställa kontrollåtgärder för import av sådant material som omfattas av dessa undantagsbestämmelser.
(21) Animaliska biprodukter som passerar gemenskapen i transit, eller som har sitt ursprung i gemenskapen och är avsedda för export, kan medföra risk för djurs och människors hälsa inom gemenskapen. Vissa krav som fastställs i denna förordning bör därför tillämpas på sådan befordran.
(22) Det lämpligaste sättet för den behöriga myndigheten på destinationsorten att få garantier för att en sändning med animaliska produkter uppfyller bestämmelserna i denna förordning är via det dokument som skall åtfölja en sådan sändning. Hälsointyget bör sparas för att det skall vara möjligt att kontrollera vart vissa importerade produkter sänds.
(23) Rådets direktiv 92/118/EEG av den 17 december 1992 om djurhälso- och hygienkrav för handel inom gemenskapen med produkter, som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A.I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG, samt för import till gemenskapen av sådana produkter(10) syftar till att uppfylla ovannämnda mål.
(24) Rådet och kommissionen har antagit flera beslut om genomförande av direktiven 90/667/EEG och 92/118/EEG. Direktiv 92/118/EEG har dessutom ändrats på ett genomgripande sätt, och ytterligare ändringar skall göras. Följaktligen finns det för närvarande ett stort antal gemenskapsrättsakter som reglerar sektorn för animaliska biprodukter och det finns behov av förenkling.
(25) En sådan förenkling kommer att leda till större öppenhet när det gäller vissa hälsobestämmelser om sådana animaliska produkter som inte är avsedda som livsmedel. En förenkling av detaljbestämmelserna i hälsolagstiftningen får dock inte leda till att området avregleras. Det är därför nödvändigt att behålla och, för att garantera människors och djurs hälsa, skärpa de detaljerade hälsobestämmelserna för animaliska produkter som inte är avsedda som livsmedel.
(26) De berörda produkterna bör omfattas av bestämmelserna om veterinära kontroller, inklusive kontroller av experter från kommissionen, och av de skyddsåtgärder som anges i rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att fullborda den inre marknaden(11).
(27) Produkter som importeras till gemenskapen bör genomgå noggranna kontroller. Detta kan uppnås genom tillämpning av de kontroller som fastställs i rådets direktiv 97/78/EG av den 18 december 1997 om principerna för organisering av veterinärkontroller av produkter från tredje land som förs in i gemenskapen(12).
(28) Direktiv 90/667/EEG, rådets beslut 95/348/EG av den 22 juni 1995 om fastställande av veterinära bestämmelser och djurhälsobestämmelser gällande Förenade kungariket och Irland för bearbetning av vissa typer av avfall avsedda att saluföras lokalt som foder för vissa kategorier av djur(13) och rådets beslut 1999/534/EG av den 19 juli 1999 om åtgärder för bearbetning av visst animaliskt avfall till skydd mot transmissibel spongiform encefalopati och om ändring av kommissionens beslut 97/735/EG(14) bör därför upphävas.
(29) För att kunna ta hänsyn till den tekniska och vetenskapliga utvecklingen bör ett nära och välfungerande samarbete mellan kommissionen och medlemsstaterna säkerställas inom ramen för den ständiga kommitté, som inrättats genom Europaparlamentets och rådets förordning (EG) nr 178/2002 av den 28 januari 2002 om allmänna principer och krav för livsmedelslagstiftning, om inrättande av Europeiska myndigheten för livsmedelssäkerhet och om förfaranden i frågor som gäller livsmedelssäkerhet(15).
(30) De åtgärder som krävs för att genomföra denna förordning bör antas enligt rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(16).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) insamling, transport, lagring, hantering, bearbetning och användning eller bortskaffande av animaliska biprodukter, så att dessa produkter inte innebär några risker för folk- eller djurhälsan,
b) utsläppande på marknaden samt, i vissa särskilda fall, export och transitering av animaliska biprodukter och därav framställda produkter enligt bilagorna VII och VIII.
2. Denna förordning skall inte tillämpas på följande:
a) Färskt sällskapsdjursfoder från detaljhandelsledet eller i anläggningar vid försäljningsställen, där styckning och lagring enbart sker i samband med försäljning direkt till konsumenten.
b) Flytande mjölk och råmjölk som bortskaffats eller använts på det ursprungliga jordbruksföretaget.
c) Hela kroppar eller delar från vilda djur som inte misstänks vara infekterade med sjukdomar som kan överföras till människor eller djur, med undantag av fisk som fiskas i kommersiellt syfte och kroppar eller delar av vilda djur som används för att tillverka jakttroféer.
d) Färskt sällskapsdjursfoder som skall användas inom det ursprungliga jordbruksföretaget, om detta foder framställts från djur som slaktats inom detta företag i syfte att användas enbart för jordbrukaren och dennes familj, i enlighet med nationell lagstiftning (husbehovsslakt).
e) Matavfall såvida inte detta
i) härrör från transportmedel i internationell trafik,
ii) är avsett som foder, eller
iii) är avsett att användas i en biogasanläggning eller för kompostering.
f) Ägg, embryon och sperma avsedda för avel.
g) Transitering med båt eller flyg.
3. Denna förordning skall inte påverka tillämpningen av sådan veterinärlagstiftning som syftar till att utrota och bekämpa vissa sjukdomar.
Artikel 2
Definitioner
1. I denna förordning avses med
a) animaliska biprodukter: hela kroppar eller delar från djur eller animaliska produkter som avses i artiklarna 4-6 som inte är avsedda att användas som livsmedel, inbegripet ägg, embryon och sperma.
b) kategori 1-material: animaliska biprodukter som avses i artikel 4.
c) kategori 2-material: animaliska biprodukter som avses i artikel 5.
d) kategori 3-material: animaliska biprodukter som avses i artikel 6.
e) djur: alla ryggradsdjur och ryggradslösa djur (inklusive fiskar, kräldjur och groddjur).
f) produktionsdjur: alla djur som hålls, göds eller föds upp av människor och används för framställning av livsmedel (bland annat kött, mjölk och ägg), ull, päls, fjädrar, skinn eller andra produkter av animaliskt ursprung.
g) vilda djur: djur som inte hålls av människor.
h) sällskapsdjur: djur av sådana arter som, utan att användas som livsmedel, i normala fall hålls och föds upp av människor i annat syfte än användning som produktionsdjur.
i) behörig myndighet: den centrala myndighet i en medlemsstat som har till uppgift att se till att kraven i denna förordning följs, eller någon annan myndighet till vilken denna centrala myndighet har delegerat denna befogenhet, särskilt när det gäller kontroll av djurfoder. Den skall även i tillämpliga fall inbegripa motsvarande myndighet i tredje land.
j) utsläppande på marknaden: all verksamhet som syftar till att sälja sådana animaliska biprodukter eller därav framställda produkter som omfattas av denna förordning till tredje man i gemenskapen eller varje annan form av överlåtelse mot betalning eller utan motprestation till sådan tredje man eller lagring för leverans till sådan tredje man.
k) handel: handel med varor mellan medlemsstaterna enligt artikel 23.2 i fördraget.
l) transitering: en befordran genom gemenskapen från ett tredje land till ett annat.
m) producent: alla producenter vars verksamhet genererar animaliska biprodukter.
n) transmissibel spongiform encefalopati (TSE): alla typer av transmissibel spongiform encefalopati, utom de som förekommer hos människor.
o) specificerat riskmaterial: det material som avses i bilaga V till Europaparlamentets och rådets förordning (EG) nr 999/2001 av den 22 maj 2001 om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati(17).
2. De särskilda definitionerna i bilaga I skall också gälla.
Artikel 3
Allmänna skyldigheter
1. Animaliska biprodukter och produkter som framställts av dessa skall samlas in, transporteras, lagras, hanteras, bearbetas, bortskaffas, släppas ut på marknaden, exporteras, transiteras och användas i enlighet med denna förordning.
2. Medlemsstaterna får dock reglera import och utsläppande på marknaden av produkter som inte anges i bilagorna VII och VIII i sin nationella lagstiftning i väntan på att ett beslut skall fattas i enlighet med det förfarande som avses i artikel 33.2. De skall omedelbart informera kommissionen om de använder sig av den möjligheten.
3. Medlemsstaterna skall, antingen var för sig eller i samarbete, se till att det finns ändamålsenliga arrangemang och tillräcklig infrastruktur för att säkerställa att kravet i punkt 1 uppfylls.
Artikel 4
a) Alla delar av kroppen, inklusive hudar och skinn, från följande djur:
i) Djur som misstänks vara infekterade med TSE enligt förordning (EG) nr 999/2001 eller som officiellt bekräftats vara infekterade med TSE.
ii) Djur som avlivats som ett led i utrotningen av TSE.
iii) Andra djur än produktionsdjur och vilda djur, särskilt inbegripet sällskapsdjur, djurparksdjur och cirkusdjur.
iv) Försöksdjur enligt definitionen i artikel 2 i rådets direktiv 86/609/EEG av den 24 november 1986 om tillnärmning av medlemsstaternas lagar och andra författningar om skydd av djur som används för försök och andra vetenskapliga ändamål(18).
v) Vilda djur som misstänks vara infekterade med sjukdomar som kan överföras till människor eller djur.
b) i) Specificerat riskmaterial.
ii) Hela kroppar från döda djur som innehåller specificerat riskmaterial om det specificerade riskmaterialet inte har avlägsnats vid tidpunkten för bortskaffandet.
c) Produkter framställda från djur som tillförts ämnen som är förbjudna enligt direktiv 96/22/EG samt produkter av animaliskt ursprung som innehåller rest av miljöföroreningar och andra ämnen som förtecknas i grupp B.3 i bilaga I till rådets direktiv 96/23/EG av den 29 april 1996 om införande av kontrollåtgärder för vissa ämnen och restsubstanser av dessa i levande djur och i produkter framställda därav och om upphävande av direktiv 85/358/EEG och 86/469/EEG samt beslut 89/187/EEG och 91/664/EEG(19), om restsubstanserna av dessa ämnen överskrider de gränsvärden som fastställs i gemenskapens lagstiftning eller, om gemenskapsgränsvärden saknas, i nationell lagstiftning.
d) Allt animaliskt material som samlas in vid rening av avloppsvatten från bearbetningsanläggningar för kategori 1-material samt från andra lokaler där specificerat riskmaterial avlägsnas, inbegripet material som avskiljts genom siktning eller i sandfång, fett- och oljeblandningar, slam och material som avlägsnats från dessa anläggningars avloppssystem, utom i de fall då detta material inte innehåller specificerat riskmaterial eller delar av sådant material.
e) Matavfall som härrör från transportmedel i internationell trafik.
f) Blandningar av kategori 1-material med antingen kategori 2-material eller kategori 3-material eller med båda, inbegripet allt material som är avsett för bearbetning i en bearbetningsanläggning för kategori 1-material.
2. Kategori 1-material skall utan onödigt dröjsmål samlas in, transporteras bort och identifieras i enlighet med artikel 7, och skall, om inte annat föreskrivs i artiklarna 23 och 24,
a) direkt bortskaffas som avfall genom förbränning i en förbränningsanläggning som godkänts i enlighet med artikel 12,
b) bearbetas enligt någon av metoderna 1-5 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, eller enligt metod 1 om den behöriga myndigheten kräver detta, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI och slutligen bortskaffas som avfall genom förbränning eller samförbränning i en förbrännings- eller samförbränningsanläggning som godkänts i enlighet med artikel 12,
c) med undantag av material som avses i punkt 1 a i och ii, bearbetas enligt bearbetningsmetod 1 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI och slutligen bortskaffas som avfall genom nedgrävning på en deponi som godkänts i enlighet med rådets direktiv 1999/31/EG av den 26 april 1999 om deponering av avfall(20),
d) när det gäller matavfall enligt punkt 1 e bortskaffas som avfall genom nedgrävning på en deponi som godkänts i enlighet med direktiv 1999/31/EG, eller
e) mot bakgrund av nya vetenskapliga rön bortskaffas med någon annan metod som godkänts i enlighet med förfarandet i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén. Denna metod kan antingen komplettera eller ersätta de metoder som föreskrivs i punkterna a-d.
3. Mellanhantering eller mellanlagring av kategori 1-material får bara genomföras på hanteringsställen för kategori 1 som godkänts enligt artikel 10.
4. Kategori 1-material får endast importeras eller exporteras i enlighet med denna förordning eller regler som fastställts i enlighet med förfarandet i artikel 33.2. Import eller export av specificerat riskmaterial får emellertid endast ske i enlighet med artikel 8.1 i förordning (EG) nr 999/2001.
Artikel 5
Kategori 2-material
1. Kategori 2-material skall omfatta animaliska biprodukter som motsvarar följande beskrivning och allt material som innehåller sådana biprodukter:
a) Naturgödsel och mag- och tarminnehåll.
b) Allt slags animaliskt material som samlats in vid rening av avloppssvatten från slakterier, utom sådana slakterier som omfattas av artikel 4.1 d, eller från bearbetningsanläggningar för kategori 2-material, inbegripet material som avskiljts genom siktning eller i sandfång, fett- och oljeblandningar, slam och material som avlägsnats från dessa anläggningars avloppssystem.
c) Produkter av animaliskt ursprung som innehåller restsubstanser av veterinärmedicinska läkemedel och föroreningar som förtecknas i grupperna B.1 och B.2 i bilaga I till direktiv 96/23/EG, om restsubstanserna av dessa ämnen överskrider gällande gränsvärden enligt gemenskapslagstiftningen.
d) Produkter av animaliskt ursprung utom, kategori 1-material, som importeras från tredje land och som under sådana inspektioner som föreskrivs i gemenskapslagstiftningen inte uppfyller veterinärmedicinska bestämmelser för import till gemenskapen, om de inte återsänds eller importen godtas med vissa förbehåll som fastställts i gemenskapslagstiftningen.
e) Djur och delar av djur, med undantag av dem som avses i artikel 4, som dött på annat sätt än genom slakt för användning som livsmedel, inbegripet djur som avlivats för att utrota någon epizootisk sjukdom.
f) Blandningar av kategori 2- och kategori 3-material, inbegripet allt material som är avsett för bearbetning i en bearbetningsanläggning för kategori 2-material.
g) Animaliska biprodukter som inte består av kategori 1- eller kategori 3-material.
2. Kategori 2-material skall utan onödigt dröjsmål samlas in, transporteras bort och identifieras i enlighet med artikel 7, och skall, om inte annat föreskrivs i artiklarna 23 och 24,
a) direkt bortskaffas som avfall genom förbränning i en förbränningsanläggning som godkänts i enlighet med artikel 12,
b) bearbetas enligt någon av metoderna 1-5 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, eller om den behöriga myndigheten kräver detta, enligt bearbetningsmetod 1, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI, och
i) omedelbart bortskaffas som avfall genom förbränning eller samförbränning i en förbrännings- eller samförbränningsanläggning som godkänts i enlighet med artikel 12, eller,
ii) när det gäller utsmält fett, bearbetas vidare till fettderivat för användning i organiska gödningsmedel eller jordförbättringsmedel eller för annan teknisk användning, förutom i kosmetika, läkemedel och medicintekniska produkter, i en kategori 2-oleokemisk anläggning som godkänts i enlighet med artikel 14,
c) bearbetas enligt bearbetningsmetod 1 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI, och
i) när det gäller uppkommet proteinhaltigt material, användas som organiskt gödningsmedel eller jordförbättringsmedel i enlighet med eventuella krav som har fastställts enligt förfarandet i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén,
ii) omvandlas i en biogas- eller komposteringsanläggning som godkänts i enlighet med artikel 15, eller
iii) bortskaffas som avfall genom nedgrävning på en deponi som godkänts i enlighet med direktiv 1999/31/EG,
d) när det gäller material som kommer från fisk, ensileras eller komposteras i enlighet med bestämmelser som har antagits enligt förfarandet i artikel 33.2,
e) när det gäller naturgödsel, från mag- och tarmsystemet avskilt mag- och tarminnehåll, mjölk och råmjölk om den behöriga myndigheten inte anser att det medför risk för spridning av allvarliga överförbara sjukdomar,
i) användas utan föregående bearbetning som råvara i en biogas- eller komposteringsanläggning som godkänts i enlighet med artikel 15 eller behandlas i en teknisk anläggning som godkänts för detta ändamål i enlighet med artikel 18,
ii) användas på mark i enlighet med denna förordning, eller
iii) omvandlas i en biogasanläggning eller komposteras i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2,
f) när det gäller hela kroppar eller delar från vilda djur som inte misstänks vara infekterade med sjukdomar som kan överföras till människor eller djur, användas för att tillverka jakttroféer i en teknisk anläggning som godkänts för detta ändamål i enlighet med artikel 18, eller
g) bortskaffas med någon annan metod, eller användas på något annat sätt, i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2 efter samråd med den berörda vetenskapliga kommittén. Denna metod eller detta sätt får antingen komplettera eller ersätta dem som föreskrivs i punkterna a-f.
3. Mellanhantering eller mellanlagring av kategori 2-material med undantag av naturgödsel får bara genomföras på hanteringsställen för kategori 2 som godkänts i enlighet med artikel 10.
4. Kategori 2-material får endast släppas ut på marknaden eller exporteras i enlighet med denna förordning eller enligt regler som fastställts i enlighet med förfarandet i artikel 33.2.
Artikel 6
Kategori 3-material
1. Kategori 3-material skall omfatta animaliska biprodukter som motsvarar följande beskrivning och allt material som innehåller sådana biprodukter:
a) Delar från slaktade djur som är tjänliga som livsmedel i enlighet med gemenskapslagstiftningen, men som av kommersiella skäl inte är avsedda som livsmedel.
b) Delar från slaktade djur som förklaras otjänliga som livsmedel trots att de inte visar några tecken på sjukdomar som kan överföras till människor eller djur, och som kommer från slaktkroppar som är tjänliga som livsmedel i enlighet med gemenskapslagstiftningen.
c) Hudar, skinn, hovar, horn, svinborst och fjädrar från djur som slaktas i ett slakteri och som har genomgått en före slaktbesiktning där de befunnits lämpade för slakt för att användas som livsmedel i enlighet med gemenskapslagstiftningen.
d) Blod från andra djur än idisslare som slaktas i ett slakteri och som har genomgått en före slaktbesiktning där de befunnits lämpade för slakt för att användas som livsmedel i enlighet med gemenskapslagstiftningen.
e) Animaliska biprodukter som erhållits vid framställning av produkter som är avsedda som livsmedel, exempelvis avfettade ben och fettgrevar.
f) Livsmedel av animaliskt ursprung eller som innehåller produkter av animaliskt ursprung, med undantag av matavfall, som inte längre är avsedda att användas som livsmedel av kommersiella skäl eller på grund av tillverkningsproblem eller förpackningsdefekter eller andra defekter som inte innebär någon risk för människor eller djur.
g) Färsk mjölk från djur som inte visar några kliniska tecken på sådana sjukdomar som kan överföras till människor eller djur via produkten i fråga.
h) Fisk och andra havslevande djur, utom havslevande däggdjur, som fångats på öppet hav för tillverkning av fiskmjöl.
i) Färska biprodukter från fisk från anläggningar som tillverkar fiskprodukter som är avsedda att användas som livsmedel.
j) Skal, biprodukter från kläckerier samt biprodukter i form av knäckägg från djur som inte visat några kliniska tecken på sådana sjukdomar som kan överföras till människor eller djur via produkten i fråga.
k) Blod, hudar, skinn, hovar, fjädrar, ull, horn, hår och päls från djur som inte visat några kliniska tecken på sådana sjukdomar som kan överföras till människor eller djur via produkten i fråga.
l) Matavfall, med undantag av matavfall enligt artikel 4.1 e.
2. Kategori 3-material skall utan onödigt dröjsmål samlas in, transporteras bort och identifieras i enlighet med artikel 7, och skall, om inte annat föreskrivs i artiklarna 23 och 24,
a) direkt bortskaffas som avfall genom förbränning i en förbränningsanläggning som godkänts i enlighet med artikel 12,
b) bearbetas i en bearbetningsanläggning som godkänts i enlighet med artikel 13 med tillämpning av någon av bearbetningsmetoderna 1-5, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI och bortskaffas som avfall, antingen genom förbränning eller samförbränning i en förbrännings- eller samförbränningsanläggning som godkänts i enlighet med artikel 12, eller på en deponi som godkänts i enlighet med direktiv 1999/31/EG,
c) bearbetas i en bearbetningsanläggning som godkänts i enlighet med artikel 17,
d) omvandlas i en teknisk anläggning som godkänts i enlighet med artikel 18,
e) användas som råvara i en anläggning för framställning av sällskapsdjursfoder som godkänts i enlighet med artikel 18,
f) omvandlas i en biogas- eller komposteringsanläggning som godkänts i enlighet med artikel 15,
g) när det gäller matavfall enligt punkt 1 l, omvandlas i en biogasanläggning eller komposteras i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2, eller i väntan på att sådana bestämmelser skall antas, i enlighet med nationell lagstiftning,
h) när det gäller material som kommer från fisk, ensileras eller komposteras i enlighet med bestämmelser som fastställts enligt förfarandet i artikel 33.2, eller
i) bortskaffas med någon annan metod, eller användas på något annat sätt, i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2, efter samråd med berörd vetenskaplig kommitté. Denna metod eller detta sätt får komplettera eller ersätta dem som föreskrivs i punkterna a-h.
3. Mellanhantering eller mellanlagring av kategori 3-material får bara genomföras på hanteringsställen för kategori 3 som godkänts i enlighet med artikel 10.
Artikel 7
Insamling, transport och lagring
1. Animaliska biprodukter och bearbetade produkter, med undantag för matavfall av kategori 3, skall samlas in, transporteras och identifieras i enlighet med bilaga II.
2. Under transporten skall ett handelsdokument, eller, när det krävs enligt denna förordning, ett hälsointyg åtfölja animaliska biprodukter och bearbetade produkter. Handelsdokument och hälsointyg skall uppfylla de krav och bevaras under den tid som anges i bilaga II. De skall särskilt innehålla uppgifter om mängden och en beskrivning av materialet och dess märkning.
3. Medlemsstaterna skall säkerställa ändamålsenliga arrangemang för att garantera att insamling och transport av kategori 1- och kategori 2-material genomförs i enlighet med bilaga II.
4. I enlighet med artikel 4 i rådets direktiv 75/442/EEG av den 15 juli 1975 om avfall(21) skall medlemsstaterna vidta nödvändiga åtgärder för att se till att matavfall av kategori 3 insamlas, transporteras och bortskaffas utan att människors hälsa äventyras eller miljön skadas.
5. Bearbetade produkter får endast lagras vid lagringsanläggningar som godkänts enligt artikel 11.
6. Medlemsstaterna får emellertid besluta att inte tillämpa bestämmelserna i denna artikel på naturgödsel som transporteras mellan två platser inom samma jordbruksföretag, eller mellan jordbruksföretag och användare som är etablerade i samma medlemsstat.
Artikel 8
Avsändande av animaliska biprodukter och bearbetade produkter till andra medlemsstater
1. Animaliska biprodukter och bearbetade produkter får sändas till andra medlemsstater endast på de villkor som anges i punkterna 2-6.
2. Mottagande medlemsstat skall ha godkänt att ta emot kategori 1-material, kategori 2-material, bearbetade produkter som härrör från kategori 1- eller kategori 2-material och bearbetat animaliskt protein. Medlemsstaten får ställa som krav för mottagandet att bearbetningsmetod 1 skall tillämpas före avsändandet.
3. Animaliska biprodukter och de bearbetade produkter som avses i punkt 2 skall
a) åtföljas av ett handelsdokument eller, när det krävs enligt denna förordning, ett hälsointyg, och
b) transporteras direkt till den mottagande anläggningen, som skall ha godkänts i enlighet med denna förordning.
4. När medlemsstater sänder kategori 1-material, kategori 2-material, bearbetade produkter som härrör från kategori 1- eller kategori 2-material och bearbetat animaliskt protein till andra medlemsstater skall den behöriga myndigheten på ursprungsorten underrätta den behöriga myndigheten på bestämmelseorten om varje avgående sändning via Animo-systemet, eller med hjälp av någon annan överenskommen metod. Meddelandet skall innehålla de upplysningar som anges i kapitel I.2 i bilaga II.
5. När den behöriga myndigheten på bestämmelseorten underrättats om en sändning i enlighet med punkt 4, skall den underrätta den behöriga myndigheten på ursprungsorten om varje sändnings ankomst via Animo-systemet, eller med hjälp av någon annan överenskommen metod.
6. Den mottagande medlemsstaten skall genom regelbundna kontroller se till att de berörda anläggningarna i det egna landet endast använder sändningarna för godkända ändamål och att de för ett fullständigt register som visar att denna förordning har följts.
Artikel 9
Register
1. Den som avsänder, transporterar eller tar emot animaliska biprodukter skall föra register över sändningarna. Registren skall innehålla de upplysningar och bevaras under den tid som anges i bilaga II.
Artikel 10
Godkännande av hanteringsställen
1. Hanteringsställen för material i kategori 1, 2 och 3 skall godkännas av den behöriga myndigheten.
2. För att kunna godkännas skall ett hanteringsställe för kategori 1- eller kategori 2-material
a) uppfylla kraven i kapitel I i bilaga III,
b) hantera och lagra kategori 1- eller kategori 2-material i enlighet med kapitel II del B i bilaga III,
c) genomgå hanteringsställets egenkontroll på det sätt som föreskrivs i artikel 25,
d) kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
3. För att kunna godkännas skall ett hanteringsställe för kategori 3-material
a) uppfylla kraven i kapitel I i bilaga III,
b) kunna hantera och lagra kategori 3-material i enlighet med kapitel II del A i bilaga III,
c) genomgå hanteringsställets egenkontroll på det sätt som föreskrivs i artikel 25,
d) kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
Artikel 11
Godkännande av lagringsanläggningar
1. Lagringsanläggningar skall godkännas av den behöriga myndigheten.
2. För att kunna godkännas skall en lagringsanläggning
a) uppfylla kraven i kapitel III i bilaga III,
b) ha kontrollerats av den behöriga myndigheten i enlighet med artikel 26.
Artikel 12
Godkännande av förbrännings- och samförbränningsanläggningar
1. Förbränning och samförbränning av bearbetade produkter skall genomföras i enlighet med bestämmelserna i direktiv 2000/76/EG. Förbränning och samförbränning av animaliska biprodukter skall antingen genomföras i enlighet med bestämmelserna i direktiv 2000/76/EG eller, då det direktivet inte är tillämpligt, i enlighet med bestämmelserna i denna förordning. Förbrännings- och samförbränningsanläggningar skall godkännas i enlighet med det direktivet eller i enlighet med punkt 2 eller 3.
2. För att godkännas av den behöriga myndigheten för bortskaffande av animaliska biprodukter, skall en förbränningsanläggning eller samförbränningsanläggning med hög kapacitet som inte omfattas av direktiv 2000/76/EG uppfylla
a) de allmänna kraven i kapitel I i bilaga IV,
b) villkoren för verksamheten i kapitel II i bilaga IV,
c) kraven i kapitel III i bilaga IV beträffande utsläpp i vattnet,
d) kraven i kapitel IV i bilaga IV beträffande restsubstanser,
e) temperaturmätningskraven i kapitel V i bilaga IV,
f) bestämmelserna för onormala driftsförhållanden i kapitel VI i bilaga IV.
3. För att godkännas av den behöriga myndigheten för bortskaffande av animaliska biprodukter, skall en förbränningsanläggning eller samförbränningsanläggning med låg kapacitet som inte omfattas av direktiv 2000/76/EG
a) användas endast för bortskaffande av döda sällskapsdjur och/eller kategori 2- och kategori 3-material,
b) när den ligger på ett jordbruksföretag endast användas för bortskaffande av material från det jordbruksföretaget,
c) uppfylla de allmänna villkoren i kapitel I i bilaga IV,
d) uppfylla de tillämpliga villkoren för verksamheten i kapitel II i bilaga IV,
e) uppfylla kraven i kapitel V i bilaga IV beträffande restsubstanser,
f) uppfylla de tillämpliga temperaturmätningskraven i kapitel V i bilaga IV, och
g) uppfylla kraven för onormala driftsförhållanden i kapitel VI i bilaga IV.
4. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
5. Kraven i punkterna 2 och 3 får ändras med beaktande av nya vetenskapliga rön i enlighet med förfarandet i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén.
Artikel 13
Godkännande av bearbetningsanläggningar för kategori 1- och kategori 2-material
1. Bearbetningsanläggningar för kategori 1- och kategori 2-material skall godkännas av den behöriga myndigheten.
2. För att kunna godkännas skall bearbetningsanläggningar för kategori 1- eller kategori 2-material
a) uppfylla kraven i kapitel I i bilaga V,
b) hantera, bearbeta och lagra kategori 1- eller kategori 2-material i enlighet med kapitel II i bilaga V samt kapitel I i bilaga VI,
c) valideras av den behöriga myndigheten i enlighet med kapitel V i bilaga V,
d) genomgå anläggningens egenkontroll på det sätt som föreskrivs i artikel 25,
e) kontrolleras av den behöriga myndigheten i enlighet med artikel 26,
f) kunna säkerställa att de bearbetade produkterna uppfyller kraven i kapitel I i bilaga VI.
3. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
Artikel 14
Godkännande av oleokemiska anläggningar för kategori 2- och kategori 3-material
1. Oleokemiska anläggningar skall godkännas av den behöriga myndigheten.
a) bearbeta utsmält fett som härrör från kategori 2-material i enlighet med kraven i kapitel III i bilaga VI,
b) införa och genomföra rutiner för övervakning och kontroll av kritiska kontrollpunkter i de processer som används,
c) föra register över de uppgifter som erhållits genom de åtgärder som anges i punkt b så att de kan läggas fram för den behöriga myndigheten,
d) kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
3. För att kunna godkännas skall en oleokemisk anläggning för kategori 3-material bearbeta utsmält fett som härrör endast från kategori 3-material och uppfylla de relevanta kraven i punkt 2.
4. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
Artikel 15
Godkännande av biogas- och komposteringsanläggningar
1. Biogas- och komposteringsanläggningar skall godkännas av den behöriga myndigheten.
2. För att kunna godkännas skall biogas- och komposteringsanläggningar
a) uppfylla kraven i kapitel II del A i bilaga VI,
b) hantera och bearbeta animaliska biprodukter i enlighet med kapitel II delarna B och C i bilaga VI,
c) kontrolleras av den behöriga myndigheten i enlighet med artikel 26,
d) införa och genomföra rutiner för övervakning och kontroll av kritiska kontrollpunkter,
e) säkerställa att rötrest och, om tillämpligt, kompost uppfyller de mikrobiologiska krav som anges i kapitel II del D i bilaga VI.
3. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
Artikel 16
Allmänna djurhälsobestämmelser
1. Medlemsstaterna skall vidta alla åtgärder som behövs för att säkerställa att de animaliska biprodukter, och därav framställda produkter som avses i bilagorna VII och VIII, inte avsänds från något jordbruksföretag som ligger i en zon som är föremål för restriktioner som införts sedan zonen drabbats av en sjukdom för vilken den djurart som produkterna härrör från är mottaglig, eller från någon anläggning eller zon från vilka förflyttning eller handel skulle medföra risker för den djurhälsostatus som berör medlemsstaterna eller vissa områden i medlemsstaterna, utom då produkterna hanteras i enlighet med denna förordning.
2. De åtgärder som avses i punkt 1 skall säkerställa att produkterna har framställts från djur som
a) kommer från ett jordbruksföretag, ett område, en del av ett område eller, när det gäller vattenbruksprodukter, från en fiskodling, en zon eller en del av en zon som inte är föremål för djurhälsorestriktioner som gäller de berörda djuren och produkterna; detta gäller särskilt restriktioner som införts i samband med åtgärder för sjukdomsbekämpning enligt gemenskapslagstiftningen eller restriktioner till följd av en allvarlig överförbar sjukdom som förtecknas i rådets direktiv 92/119/EEG av den 17 december 1992 om införande av allmänna gemenskapsåtgärder för bekämpning av vissa djursjukdomar och särskilda åtgärder mot vesikulär svinsjuka(22),
b) inte har slaktats i en anläggning där det vid tidpunkten för slakt fanns djur som var infekterade eller som misstänktes vara infekterade med någon av de sjukdomar som omfattas av de bestämmelser som avses i punkt a.
3. Förutsatt att de villkor som gäller sådana åtgärder för sjukdomsbekämpning som avses i punkt 2 a är uppfyllda, skall det vara tillåtet att på marknaden släppa ut animaliska biprodukter, och sådana därav framställda produkter som avses i bilagorna VII och VIII, som kommer från ett område eller en del av ett område som är föremål för djurhälsorestriktioner men som inte är infekterade eller misstänks vara infekterade, förutsatt att produkterna, allt efter omständigheterna
a) har framställts, hanterats, transporterats och lagrats avskilt från, eller vid andra tidpunkter än produkter som uppfyller alla djurhälsovillkor,
b) har genomgått en behandling som är tillräcklig för att eliminera de aktuella djurhälsoriskerna i enlighet med denna förordning vid en anläggning som har godkänts för detta ändamål av den medlemsstat där djurhälsoproblemet förekom,
c) har identifierats på ett korrekt sätt,
d) uppfyller de särskilda krav som anges i bilagorna VII och VIII, eller de närmare bestämmelser som skall fastställas i enlighet med förfarandet i artikel 33.2.
Andra villkor än de som anges i första stycket får fastställas i särskilda situationer genom beslut som antas i enlighet med det förfarande som avses i artikel 33.2. I sådana beslut skall de åtgärder som rör djuren eller de prov som djuren skall bli föremål för beaktas, liksom de egenskaper hos sjukdomen som är kännetecknande för arten i fråga, och alla åtgärder som krävs för att säkerställa skyddet av djurhälsan i gemenskapen skall specificeras.
Artikel 17
Godkännande av bearbetningsanläggningar för kategori 3-material
1. Bearbetningsanläggningar för kategori 3-material skall godkännas av den behöriga myndigheten.
2. För att kunna godkännas skall en bearbetningsanläggning för kategori 3-material
a) uppfylla kraven i kapitel I i bilaga V och kapitel I i bilaga VII,
b) hantera, bearbeta och lagra endast kategori 3-material i enlighet med kapitel II i bilaga V och bilaga VII,
c) valideras av den behöriga myndigheten i enlighet med kapitel V i bilaga V,
d) genomgå anläggningens egenkontroll på det sätt som föreskrivs i artikel 25,
e) kontrolleras av den behöriga myndigheten i enlighet med artikel 26,
f) kunna säkerställa att de bearbetade produkterna uppfyller kraven i kapitel I i bilaga VII.
3. Godkännandet skall omedelbart återkallas om villkoren för godkännandet inte längre uppfylls.
Artikel 18
Godkännande av anläggningar för tillverkning av sällskapsdjursfoder och av tekniska anläggningar
1. Anläggningar för tillverkning av sällskapsdjursfoder och tekniska anläggningar skall godkännas av den behöriga myndigheten.
2. För att en anläggning för tillverkning av sällskapsdjursfoder eller en teknisk anläggning skall kunna godkännas, skall följande krav vara uppfyllda:
a) I enlighet med de särskilda kraven i bilaga VIII för de produkter som anläggningen framställer skall den åta sig att
i) uppfylla de särskilda krav på produktionen som ställs i denna förordning,
ii) införa och genomföra rutiner för övervakning och kontroll av kritiska kontrollpunkter i de processer som används,
iii) beroende på vilken produkt det gäller, ta prover som sedan analyseras på ett laboratorium som godkänts av den behöriga myndigheten, så att det kan kontrolleras att kraven i denna förordning är uppfyllda,
iv) föra register över de uppgifter som erhållits i enlighet med ii och iii och hålla dem tillgängliga för den behöriga myndigheten. Resultaten från kontroller och tester skall sparas i minst två år,
v) underrätta den behöriga myndigheten om resultatet av den laboratorieanalys som avses i iii eller annan information som de ansvariga för anläggningen har tillgång till, visar att det föreligger allvarlig fara för djurs eller människors hälsa.
b) Anläggningen skall kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
3. Godkännandet skall omedelbart återkallas om villkoren för godkännandet inte längre uppfylls.
Artikel 19
Utsläppande på marknaden och export av bearbetat animaliskt protein och andra bearbetade produkter som skulle kunna användas som foderråvara
Medlemsstaterna skall se till att bearbetat animaliskt protein och andra bearbetade produkter som skulle kunna användas som foderråvara släpps ut på marknaden eller exporteras endast om de
a) har framställts i en bearbetningsanläggning för kategori 3-material som har godkänts och står under tillsyn i enlighet med artikel 17,
b) har framställts enbart av sådant kategori 3-material som förtecknas i bilaga VII,
c) har hanterats, bearbetats, lagrats och transporterats i enlighet med bilaga VII och på ett sådant sätt att det säkerställs att artikel 22 följs,
d) uppfyller de särskilda kraven i bilaga VII.
Artikel 20
Utsläppande på marknaden och export av sällskapsdjursfoder, tuggben och tekniska produkter
1. Medlemsstaterna skall se till att sällskapsdjursfoder, tuggben, tekniska produkter, med undantag av dem som avses i punkterna 2 och 3, samt de animaliska biprodukter som avses i bilaga VIII släpps ut på marknaden eller exporteras endast om de
a) antingen
i) uppfyller de särskilda kraven i bilaga VIII, eller
ii) om en produkt kan användas både som en teknisk produkt och som foderråvara och bilaga VIII inte innehåller några särskilda krav, uppfyller de särskilda kraven i det relevanta kapitlet i bilaga VII,
b) kommer från anläggningar som har godkänts och står under tillsyn i enlighet med artikel 18 eller, när det gäller de animaliska biprodukter som avses i bilaga VIII, från andra anläggningar som har godkänts i enlighet med gemenskapens veterinärlagstiftning.
2. Medlemsstaterna skall se till att organiska gödningsmedel och jordförbättringsmedel som är framställda av bearbetade produkter, såvida de inte framställts av naturgödsel och mag- och tarminnehåll, släpps ut på marknaden eller exporteras endast om de uppfyller eventuella krav som fastställts i enlighet med det förfarande som avses i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén.
3. Medlemsstaterna skall se till att fettderivat som är framställda av kategori 2-material släpps ut på marknaden eller exporteras endast om de
a) har framställts av utsmält fett som kommer från bearbetning av kategori 2-material i en bearbetningsanläggning för kategori 2-material som godkänts i enlighet med artikel 13 med tillämpning av någon av bearbetningsmetoderna 1-5 i en oleokemisk anläggning för kategori 2-material som har godkänts i enlighet med artikel 14,
b) har hanterats, bearbetats, lagrats och transporterats i enlighet med bilaga VI,
c) uppfyller eventuella särskilda krav i bilaga VIII.
Artikel 21
Skyddsåtgärder
Artikel 10 i direktiv 90/425/EEG skall tillämpas på de produkter som omfattas av bilagorna VII och VIII till denna förordning.
Artikel 22
Begränsningar i användningen
1. Följande användningar av animaliska biprodukter och bearbetade produkter skall vara förbjudna:
a) Utfodring av ett djurslag med animaliskt protein som härrör från djurkroppar eller delar av djur av samma art.
b) Utfodring av produktionsdjur, med undantag av pälsdjur, med matavfall eller foderråvara som innehåller eller framställts av matavfall.
c) Användning av andra typer av organiska gödningsmedel eller jordförbättringsmedel än naturgödsel på betesmark.
2. Genomförandebestämmelser till denna artikel, inbegripet bestämmelser som rör kontrollåtgärder, skall antas i enlighet med det förfarande som avses i artikel 33.2. Undantag från punkt 1 a får beviljas för fisk och pälsdjur i enlighet med samma förfarande, efter samråd med den berörda vetenskapliga kommittén.
Artikel 23
Undantag när det gäller användning av animaliska biprodukter
1. Medlemsstaterna får, under de behöriga myndigheternas tillsyn, godkänna följande:
a) Användning av animaliska biprodukter för diagnostisk verksamhet samt i undervisnings- och forskningssyfte.
b) Användning av animaliska biprodukter för taxidermiska ändamål i tekniska anläggningar som godkänts för detta syfte i enlighet med artikel 18.
2. a) Medlemsstaterna får även godkänna användning av de animaliska biprodukter som anges i stycke b för utfodring av de djur som anges i stycke c under de behöriga myndigheternas tillsyn och i enlighet med reglerna i bilaga IX.
b) De animaliska biprodukter som avses i stycke a är följande:
i) Kategori 2-material under förutsättning att det kommer från djur som inte avlivats eller dött till följd av bekräftad eller förmodad förekomst av en sjukdom som kan överföras till människor eller djur.
ii) Kategori 3-material som avses i artikel 6.1 a-6.1 j och, om inte annat följer av artikel 22, i artikel 6.1 l.
c) De djur som avses i stycke a är följande:
i) djurparksdjur,
ii) cirkusdjur,
iii) andra kräldjur och rovfåglar än djurparksdjur och cirkusdjur,
iv) pälsdjur,
v) vilda djur vars kött inte är avsett som livsmedel,
vi) hundar från etablerade kennlar eller grupper av sådana hundar som jakt- eller draghundar,
vii) fluglarver som skall användas som fiskagn.
d) Medlemsstaterna får dessutom, under de behöriga myndigheternas tillsyn, tillåta användning av sådant kategori 1-material som avses i artikel 4.1 b ii för utfodring av utrotningshotade eller skyddade arter av asätande fåglar enligt regler som har fastställts i enlighet med det förfarande som anges i artikel 33.2, efter samråd med Europeiska myndigheten för livsmedelssäkerhet.
3. Medlemsstaterna skall informera kommissionen om
a) användningen av de undantag som avses i punkt 2,
b) de kontroller som införs för att säkerställa att de animaliska biprodukterna i fråga endast används för godkända ändamål.
4. Varje medlemsstat skall upprätta en förteckning över de användare och uppsamlingscentraler i det egna landet som godkänts och registrerats i enlighet med punkt 2 c iv, vi och vii. Varje användare och uppsamlingscentral skall tilldelas ett officiellt nummer för kontrolländamål och för att produkterna i fråga skall kunna spåras till sitt ursprung.
Den behöriga myndigheten skall utöva tillsyn över de i föregående stycke omnämnda användarnas och uppsamlingscentralernas anläggningar och skall när som helst kunna få tillträde till alla delar av anläggningarna, för att kunna kontrollera att de krav som avses i punkt 2 har uppfyllts.
Om det vid en sådan inspektion visar sig att dessa krav inte har uppfyllts skall den behöriga myndigheten vidta lämpliga åtgärder.
5. Närmare bestämmelser om kontrollåtgärder får antas i enlighet med det förfarande som avses i artikel 33.2.
Artikel 24
Undantag i fråga om bortskaffande av animaliska biprodukter
1. Den behöriga myndigheten får vid behov besluta att
a) döda sällskapsdjur omedelbart får bortskaffas som avfall genom nedgrävning,
b) följande animaliska biprodukter med ursprung i avlägsna områden får bortskaffas som avfall genom förbränning eller nedgrävning på platsen:
i) kategori 1-material som avses i artikel 4.1 b ii,
ii) kategori 2-material,
iii) kategori 3-material,
c) animaliska biprodukter får bortskaffas som avfall genom förbränning eller nedgrävning på platsen vid utbrott av en sjukdom som anges i A-listan från Internationella byrån för epizootiska sjukdomar (OIE) om den behöriga myndigheten avvisar transport till närmaste förbrännings- eller bearbetningsanläggning på grund av risken för spridning av hälsorisker eller på grund av att ett omfattande utbrott av en epizootisk sjukdom leder till kapacitetsbrist på sådana anläggningar.
2. Inget undantag får beviljas för kategori 1-material som avses i artikel 4.1 a i.
3. När det gäller kategori 1-material som avses i artikel 4.1 b ii får förbränning och nedgrävning utföras i enlighet med punkt 1 b eller c endast om den behöriga myndigheten godkänner och övervakar den metod som används och är övertygad om att den utesluter varje risk för överföring av TSE.
4. Medlemsstaterna skall informera kommissionen om
a) huruvida de använder möjligheterna enligt punkt 1 b när det gäller kategori 1- och kategori 2-material,
b) vilka områden de kategoriserar som avlägsna områden vid tillämpning av punkt 1 b och skälen till denna kategorisering.
5. Den behöriga myndigheten skall vidta nödvändiga åtgärder för att
a) säkerställa att förbränningen eller nedgrävningen av animaliska biprodukter inte hotar djurs eller människors hälsa,
b) hindra att animaliska biprodukter överges, dumpas eller bortskaffas på ett okontrollerat sätt.
6. Närmare bestämmelser för genomförandet av denna artikel får fastställas i enlighet med förfarandet i artikel 33.2.
Artikel 25
Anläggningarnas egenkontroll
1. Ansvariga för eller ägare till hanteringsställen och bearbetningsanläggningar eller deras företrädare skall vidta alla nödvändiga åtgärder för att uppfylla kraven i denna förordning. De skall införa, genomföra och upprätthålla ett permanent förfarande som utarbetats i enlighet med principerna för systemet för riskbedömning och kritiska kontrollpunkter (HACCP). De skall särskilt
a) identifiera och kontrollera de kritiska kontrollpunkterna i anläggningarna,
b) införa och genomföra rutiner för övervakning och kontroll av sådana kritiska kontrollpunkter i processen,
c) när det gäller bearbetningsanläggningar, ta representativa prov för att kontrollera att
i) varje bearbetad sats uppfyller produktkraven enligt denna förordning, och
ii) ligger inom de gränsvärden för fysisk-kemiska restsubstanser som anges i gemenskapslagstiftningen,
d) föra register över resultaten av de kontroller och tester som avses i styckena b och c, och bevara dessa i minst två år, så att de behöriga myndigheterna kan ta del av dem,
e) införa ett system som säkerställer att varje avsänt parti kan spåras.
2. Om resultatet av ett test som utförts på ett prov som tagits enligt punkt 1 c inte uppfyller bestämmelserna i denna förordning skall den ansvarige för bearbetningsanläggningen
a) omedelbart ge den behöriga myndigheten all relevant information om typen av prov och om det parti från vilket det tagits,
b) fastställa orsakerna till att bestämmelserna inte uppfyllts,
c) under den behöriga myndighetens tillsyn bortskaffa den kontaminerade satsen eller låta den genomgå förnyad bearbetning,
d) se till att inget material som konstaterats eller misstänks vara smittat avlägsnas från anläggningen innan det genomgått förnyad bearbetning under den behöriga myndighetens tillsyn samt förnyad officiell provtagning, så att kraven i denna förordning uppfylls, såvida det inte skall bortskaffas,
e) göra fler provtagningar och kontroller av produktionen,
f) granska de register över obearbetade animaliska biprodukter som är av betydelse för det färdiga provet,
g) införa lämpliga dekontaminerings- och rengöringsmetoder på anläggningen.
3. Närmare bestämmelser för genomförandet av denna artikel, inbegripet regler om hur ofta kontroller skall ske och om referensmetoder för mikrobiologiska analyser, får fastställas i enlighet med förfarandet i artikel 33.2.
Artikel 26
Officiella kontroller och förteckningar över godkända anläggningar
1. Den behöriga myndigheten skall genomföra regelbundna inspektioner och utöva regelbunden tillsyn vid anläggningar som godkänts i enlighet med denna förordning. Inspektioner och tillsyn vid bearbetningsanläggningar skall utföras i enlighet med kapitel IV i bilaga V.
2. Hur ofta inspektioner och tillsyn skall genomföras beror på anläggningens storlek, vilken typ av produkter som tillverkas, vilka riskbedömningar som gjorts samt vilka garantier som lämnats i enlighet med principerna för systemet för riskbedömning och kritiska kontrollpunkter (HACCP).
3. Om de besiktningar som utförs av den behöriga myndigheten visar att ett eller flera krav i denna förordning inte har uppfyllts, skall den behöriga myndigheten vidta lämpliga åtgärder.
4. Varje medlemsstat skall upprätta en förteckning över de anläggningar på dess territorium som godkänts i enlighet med denna förordning. Varje anläggning skall av medlemsstaten tilldelas ett officiellt nummer som identifierar anläggningen med hänsyn till den typ av verksamhet som bedrivs. Medlemsstaten skall sända kopior av förteckningen samt uppdaterade versioner till kommissionen och övriga medlemsstater.
5. Närmare bestämmelser för genomförandet av denna artikel, inbegripet regler om hur ofta kontroller skall ske och om referensmetoder för mikrobiologiska analyser, får fastställas i enlighet med det förfarande som avses i artikel 33.2.
Artikel 27
Gemenskapens kontroller i medlemsstaterna
1. Experter från kommissionen får, när så krävs för en enhetlig tillämpning av denna förordning, i samarbete med de behöriga myndigheterna i medlemsstaterna genomföra kontroller på plats. Den medlemsstat på vars territorium en inspektion företas skall ge all nödvändig hjälp till experterna så att de kan fullgöra sina uppgifter. Kommissionen skall informera den behöriga myndigheten om resultaten av de genomförda kontrollerna.
Artikel 28
Allmänna bestämmelser
De bestämmelser som skall tillämpas vid import från tredje land av de produkter som avses i bilagorna VII och VIII får varken vara fördelaktigare eller mindre fördelaktiga än de som gäller för produktion och saluföring av motsvarande produkter i gemenskapen.
Det skall dock vara tillåtet att importera sällskapsdjursfoder och råvaror för produktion av sådant foder från tredje land även om detta foder och dessa råvaror kommer från djur som har behandlats med vissa ämnen som är förbjudna enligt direktiv 96/22/EG, under förutsättning att dessa råvaror är permanent märkta och i enlighet med vissa särskilda villkor, som fastställts i enlighet med förfarandet i artikel 33.2.
Artikel 29
Förbud och efterlevnad av gemenskapsbestämmelser
1. Det skall vara förbjudet att importera eller transitera animaliska biprodukter och bearbetade produkter om det inte sker i enlighet med denna förordning.
2. De produkter som avses i bilagorna VII och VIII får importeras till eller transiteras genom gemenskapen endast om de uppfyller kraven i punkterna 3-6.
3. De produkter som avses i bilagorna VII och VIII skall, om inte något annat anges i dessa bilagor, komma från ett tredje land eller en del av ett tredje land som återfinns på en sådan förteckning som skall upprättas och uppdateras i enlighet med förfarandet i artikel 33.2.
Förteckningen får samordnas med andra förteckningar som upprättats av folk- och djurhälsoskäl.
När förteckningen upprättas skall särskilt följande beaktas:
a) Det tredje landets lagstiftning.
b) Hur den behöriga myndigheten i det tredje landet och dess inspektörer är organiserade, vilka befogenheter som inspektörerna har, vilken tillsyn inspektörerna är underkastade, samt inspektörernas behörighet att effektivt övervaka hur landets lagstiftning tillämpas.
c) De faktiska hälsovillkor som tillämpas på produktion, framställning, hantering, lagring och avsändande av produkter av animaliskt ursprung som är avsedda för gemenskapen.
d) Vilka garantier det tredje landet kan ge för att gällande hygienkrav uppfylls.
e) Erfarenheter från saluföringen av produkten från det tredje landet samt resultaten av de införselkontroller som genomförts.
f) Resultatet från eventuella gemenskapsinspektioner i det tredje landet.
g) Hälsostatus för livsmedelsproducerande djur samt för andra tamdjur och vilda djur i det tredje landet, med särskilt beaktande av exotiska djursjukdomar och alla sådana aspekter av den allmänna hälsosituationen i landet som skulle kunna innebära en risk för folk- eller djurhälsan i gemenskapen.
h) Hur snabbt och regelbundet det tredje landet tillhandahåller uppgifter om förekomsten av infektiösa eller smittsamma djursjukdomar på dess territorium, särskilt de sjukdomar som anges i OIE:s A-lista och B-lista eller, beträffande sjukdomar hos vattenbruksdjur, de anmälningspliktiga sjukdomar som förtecknas i OIE:s hälsokodex för vattenlevande djur.
i) De bestämmelser om förebyggande och bekämpning av infektiösa eller smittsamma djursjukdomar som gäller i det tredje landet samt tillämpningen av dessa, inklusive bestämmelser om import från andra länder.
4. De produkter som avses i bilagorna VII och VIII, med undantag av tekniska produkter, skall komma från en anläggning som finns upptagen på en gemenskapsförteckning som upprättats i enlighet med det förfarande som avses i artikel 33.2, på grundval av ett meddelande till kommissionen från de behöriga myndigheterna i det tredje landet i vilket det intygas att anläggningen uppfyller gemenskapens krav och att officiella inspektörer i det tredje landet ansvarar för tillsynen av anläggningen.
Godkända förteckningar skall ändras enligt följande:
a) Kommissionen skall underrätta medlemsstaterna om det tredje landets förslag till ändringar av förteckningen över anläggningar inom fem arbetsdagar från det att förslaget till ändringar från det tredje landet tagits emot.
b) Medlemsstaterna skall, inom sju arbetsdagar från det att de tagit emot de förslag till ändringar av förteckningen över anläggningar som avses i punkt a, skriftligen meddela kommissionen sina synpunkter på dessa förslag.
c) Om minst en medlemsstat har lämnat skriftliga synpunkter skall kommissionen inom fem arbetsdagar underrätta övriga medlemsstater om detta samt föra upp ärendet som en punkt på dagordningen till Ständiga kommitténs för livsmedelskedjan och djurhälsa nästa sammanträde för avgörande, i enlighet med förfarandet i artikel 33.2.
d) Om kommissionen inte har erhållit några synpunkter från medlemsstaterna inom den tidsfrist som anges i punkt b, skall medlemsstaterna anses ha godtagit ändringarna i förteckningen. Kommissionen skall underrätta medlemsstaterna om dessa ändringar inom fem arbetsdagar, och import från de berörda anläggningarna skall vara tillåten fem arbetsdagar efter det att medlemsstaterna tagit emot denna underrättelse.
5. De tekniska produkter som avses i bilaga VIII skall komma från anläggningar som har godkänts och registrerats av de behöriga myndigheterna i det tredje landet.
6. Sändningar av de produkter som avses i bilagorna VII och VIII skall, om inte något annat anges i dessa bilagor, åtföljas av ett hälsointyg som utformats enligt förlagan i bilaga X och som bestyrker att produkterna uppfyller de villkor som avses i dessa bilagor samt att de kommer från anläggningar som säkerställer att dessa villkor uppfylls.
7. I väntan på att förteckningen enligt punkt 4 skall upprättas och att de förlagor till intyg som avses i punkt 6 skall antas, får medlemsstaterna behålla de kontroller som föreskrivs i direktiv 97/78/EG och de intyg som föreskrivs enligt gällande nationella bestämmelser.
Artikel 30
Likvärdighet
1. I enlighet med förfarandet i artikel 33.2 får det fattas ett beslut genom vilket det erkänns att de hälsobestämmelser som tillämpas av ett tredje land, en grupp av tredje länder eller en region i ett tredje land vid produktion, framställning, hantering, lagring och transport av en eller flera av de produktkategorier som avses i bilagorna VII och VIII, innebär garantier som är likvärdiga med dem som tillämpas i gemenskapen förutsatt att det tredje landet kan visa detta på ett objektivt sätt.
I beslutet skall fastställas vilka villkor som gäller för import och/eller transitering av animaliska biprodukter från denna region, detta land eller denna grupp av länder.
2. De villkor som avses i punkt 1 skall omfatta
a) vilken typ av hälsointyg som skall åtfölja produkten samt intygets innehåll,
b) vilka särskilda hälsokrav som skall gälla för import till och/eller transitering genom gemenskapen,
c) vid behov, förfaranden för att upprätta och ändra förteckningar över regioner eller anläggningar från vilka import och/eller transitering är tillåten.
3. Närmare bestämmelser för tillämpningen av denna artikel skall fastställas i enlighet med förfarandet i artikel 33.2.
Artikel 31
Gemenskapens inspektioner och granskningar
1. Experter från kommissionen får, när så är lämpligt, tillsammans med experter från medlemsstaterna genomföra kontroller på plats för att
a) upprätta en förteckning över tredje länder eller delar av tredje länder samt för att fastställa villkor för import och/eller transitering,
b) kontrollera efterlevnaden av
i) villkoren för införande i en gemenskapsförteckning över tredje länder,
ii) villkoren för import och/eller transitering,
iii) villkoren för erkännande av att åtgärder är likvärdiga,
iv) alla slags nödåtgärder som tillämpas med stöd av gemenskapslagstiftningen.
De experter från medlemsstaterna som ansvarar för kontrollerna skall utses av kommissionen.
2. De kontroller som avses i punkt 1 skall utföras på gemenskapens vägnar och på gemenskapens bekostnad.
3. Hur ofta samt på vilket sätt kontrollerna i punkt 1 skall utföras får fastställas i enlighet med förfarandet i artikel 33.2.
4. Om det vid en kontroll enligt punkt 1 uppdagas allvarliga överträdelser av hälsobestämmelserna, skall kommissionen omedelbart begära att det tredje landet vidtar lämpliga åtgärder eller tillfälligt stoppa sändningarna av produkter och genast underrätta medlemsstaterna.
Artikel 32
Ändring av bilagor samt övergångsbestämmelser
1. Efter samråd med berörd vetenskaplig kommitté i frågor som kan ha betydelse för djurs och människors hälsa får bilagorna ändras eller kompletteras och lämpliga övergångsbestämmelser antas i enlighet med förfarandet i artikel 33.2.
2. När det gäller förbudet mot utfodring med matavfall som fastställs i artikel 22 skall, i medlemsstater där lämpliga kontrollsystem finns innan denna förordning börjar tillämpas, övergångsåtgärder vidtas, i enlighet med första stycket, för att tillåta fortsatt användning av vissa typer av matavfall under noga kontrollerade förhållanden under en period på högst fyra år från och med den 1 november 2002. Genom åtgärderna skall det garanteras att det inte finns några onödiga risker för djurs hälsa eller folkhälsan under övergångsperioden.
Artikel 33
Föreskrivande förfarande
1. Kommissionen skall biträdas av Ständiga kommittén för livsmedelskedjan och djurhälsa, nedan kallad "kommittén".
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara 15 dagar.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 34
Samråd med vetenskapliga kommittéer
Samråd skall genomföras med de berörda vetenskapliga kommittéerna i alla frågor inom denna förordnings tillämpningsområde som kan påverka människors eller djurs hälsa.
Artikel 35
Nationella bestämmelser
1. Medlemsstaterna skall till kommissionen överlämna texterna till nationell lagstiftning som de antar inom det område som omfattas av denna förordning.
2. I synnerhet skall medlemsstaterna informera kommissionen om de åtgärder som vidtas för att se till att bestämmelserna i denna förordning iakttas senast ett år efter dess ikraftträdande. På grundval av den information som den erhåller skall kommissionen lägga fram en rapport för Europaparlamentet och rådet, i förekommande fall åtföljd av lagförslag.
3. Medlemsstaterna får anta eller bibehålla nationella bestämmelser som i större utsträckning än denna förordning begränsar användningen av organiska gödningsmedel och jordförbättringsmedel i väntan på att gemenskapsregler skall antas för användningen av dessa medel, i enlighet med artikel 20.2. Medlemsstaterna får anta eller bibehålla nationella bestämmelser som i större utsträckning än denna förordning begränsar användningen av fettderivat som framställts ur kategori 2-material i avvaktan på ett tillägg till bilaga VIII av gemenskapsregler för deras användning i enlighet med artikel 32.
Artikel 36
Finansiella arrangemang
Kommissionen skall utarbeta en rapport om hur medlemsstaterna finansierar bearbetning, insamling, lagring och bortskaffande av animaliska biprodukter, och rapporten skall åtföljas av lämpliga förslag.
Artikel 37
Upphävande
Direktiv 90/667/EEG samt besluten 95/348/EG och 1999/534/EG skall upphöra att gälla sex månader efter det att denna förordning trätt i kraft.
Hänvisningar till direktiv 90/667/EEG skall från den dagen förstås som hänvisningar till denna förordning.
Artikel 38
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1802/2002
av den 10 oktober 2002
om rättelse av förordning (EG) nr 1282/2002 om ändring av bilagorna till rådets direktiv 92/65/EEG om fastställande av djurhälsokrav i handeln inom och importen till gemenskapen av djur, sperma, ägg (ova) och embryon som inte faller under de krav som fastställs i de specifika gemenskapsregler som avses i bilaga A.I till direktiv 90/425/EEG
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING,
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 92/65/EEG av den 13 juli 1992 om fastställande av djurhälsokrav i handeln inom och importen till gemenskapen av djur, sperma, ägg (ova) och embryon som inte faller under de krav som fastställs i de specifika gemenskapsregler som avses i bilaga A.I till direktiv 90/425/EEG(1), senast ändrat genom kommissionens förordning (EG) nr 1282/2002(2), särskilt artikel 22 i detta, och
av följande skäl:
(1) Förordning (EG) nr 1282/2002 om ändring av direktiv 92/65/EEG antogs den 15 juli 2002.
(2) För att ge tillräckligt med tid för att de nya bestämmelserna skulle kunna införas i samtliga medlemsstater borde det ha fastställts ett datum då förordning (EG) nr 1282/2002 skulle börja att tillämpas.
(3) Under antagandeprocessen fastställdes emellertid inte något sådant datum.
(4) Förordning (EG) nr 1282/2002 bör därför rättas.
(5) Det är nödvändigt att rättelsen gäller från och med det datum då förordning (EG) nr 1282/2002 träder i kraft.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 2 i förordning (EG) nr 1282/2002 skall följande läggas till som andra stycke: "Den skall tillämpas från och med den 1 mars 2003."
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
Rådets förordning (EG) nr 1881/2002
av den 14 oktober 2002
om rättelse av förordning (EG) nr 2200/96 när det gäller startdatum för övergångsperioden för erkännande av producentorganisationer
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
av följande skäl:
(1) I enlighet med artikel 13.1 i rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(4) beviljades en övergångsperiod på två år, med början samma dag som ikraftträdandet, under vilken bestämmelserna i avdelning IV i ovannämnda förordning skulle gälla, till producentorganisationer som erkänts enligt förordning (EEG) nr 1035/72(5), men som inte uppfyllde kraven för erkännande enligt förordning (EG) nr 2200/96. Denna tvååriga övergångsperiod kan förlängas till fem år om medlemsstaten i fråga godkänner en handlingsplan som läggs fram av producentorganisationen över hur denna skall uppfylla kraven i förordning (EG) nr 2200/96 för att erkännas av den medlemsstaten.
(2) I artikel 13.1 i förordning (EG) nr 2200/96 fastställs att det datum då de två- och femåriga övergångsperioderna inleds skall vara det datum förordningen träder i kraft, dvs. den 21 november 1996. Detta är ett misstag; faktum är att det skulle ha varit meningslöst att låta övergångsåtgärder vara stödberättigande från och med datumet för ikraftträdande av förordning (EG) nr 2200/96, eftersom förordning (EEG) nr 1035/72 gällde fram till och med den 31 december 1996. Övergångsperioderna i fråga borde ha inletts i och med tillämpningsdatumet för förordning (EG) nr 2200/96.
(3) Således bör nämnda misstag i artikel 13.1 i förordning (EG) nr 2200/96 rättas. Eftersom effekterna av misstaget kan ha haft negativa effekter för producentorganisationer som har utnyttjat övergångsperioderna bör motsvarande bestämmelser tillämpas från och med tillämpningsdatumet för förordning (EG) nr 2200/96.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 13.1 i förordning (EG) nr 2200/96 skall ersättas med följande: "1. De producentorganisationer som före den här förordningens ikraftträdande har erkänts med stöd av förordning (EEG) nr 1035/72, och som inte utan en övergångsperiod kan erkännas med stöd av artikel 11 i den här förordningen, får fortsätta att verka inom ramen för avdelning IV under två år från och med den 1 januari 1997, om dessa organisationer uppfyller kraven i berörda artiklar i förordning (EEG) nr 1035/72."
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1921/2002
av den 28 oktober 2002
om ändring av förordning (EEG) nr 3149/92 om närmare bestämmelser för leverans av livsmedel från interventionslager till förmån för de sämst ställda i gemenskapen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3730/87 av den 10 december 1987 om allmänna bestämmelser för leverans av livsmedel från interventionslager till utsedda organisationer för utdelning till de sämst ställda i gemenskapen(1), ändrad genom förordning (EG) nr 2535/95(2), särskilt artikel 6 i denna, och
av följande skäl:
(1) Enligt artikel 3 i kommissionens förordning (EEG) nr 3149/92(3), senast ändrad genom förordning (EEG) nr 1098/2001(4), skall den årliga planen för utdelning av livsmedel till de sämst ställda genomföras under perioden 1 oktober-30 september följande år. För att interventionslagren skall kunna förvaltas på bästa sätt bör de produkter som skall delas ut tas ut ur lagren senast den 31 augusti under genomförandeåret.
(2) I artikel 5 i förordning (EEG) nr 3149/92 fastställs bokföringsvärdet för de produkter som ställs till förfogande. Denna bestämmelse bör ändras för att hänsyn skall kunna tas till de ändringar som gjorts i interventionssystemet inom den gemensamma organisationen av marknaden för nötkött.
(3) Artikel 8 i förordning (EEG) nr 3149/92, som inte längre tillämpas eftersom ersättning för transportkostnaderna betalas ut på basis av faktiska utgifter, bör utgå.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från berörda förvaltningskommittéer.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 3149/92 ändras på följande sätt:
1. I artikel 3.1 skall följande läggas till som andra stycke:"Uttag av produkter från interventionslagren skall ske från och med den 1 oktober till och med den 31 augusti följande år."
2. Artikel 5 skall ersättas med följande:
"Artikel 5
1. I EUGFJ:s (garantisektionen) bokföring, och utan att det påverkar tillämpningen av artikel 8 i förordning (EEG) nr 1883/78(5), skall bokföringsvärdet för de interventionsprodukter som ställs till förfogande enligt den här förordningen vara detsamma som gällande interventionspris den 1 oktober varje räkenskapsår.
För nötkött skall bokföringsvärdet vara detsamma som gällande interventionspris den 30 juni 2002. Detta pris skall multipliceras med den koefficient som anges i bilagan.
För de medlemsstater som inte har infört euron skall interventionsprodukternas bokföringsvärde omräknas till den nationella valutan med hjälp av den växelkurs som gällde den 1 oktober.
2. Om interventionsprodukter transporteras från en medlemsstat till en annan skall den levererande medlemsstaten bokföra den levererade produkten till ett värde av noll, och destinationsmedlemsstaten skall bokföra produkten som intäkt under uttagsmånaden, till det pris som fastställs enligt punkt 1."
3. Artikel 8 skall utgå.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 1947/2002
av den 31 oktober 2002
om ändring av förordning (EG) nr 3223/94 om tillämpningsföreskrifter till importsystemet för frukt och grönsaker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom förordning (EG) nr 545/2002(2), särskilt artikel 32.5 i denna, och
av följande skäl:
(1) De belgiska och italienska myndigheterna har meddelat kommissionen att marknaderna i Antwerpen och Bologna inte längre är representativa importmarknader för frukt och grönsaker. Dessa marknader bör därför strykas från förteckningen i artikel 3.1 i kommissionens förordning (EG) nr 3223/94(3), senast ändrad genom förordning (EG) nr 453/2002(4).
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för färsk frukt och färska grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"- Belgien och Luxemburg: Bryssel".
2. Åttonde strecksatsen skall ersättas med följande:
"- Italien: Milano".
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets förordning (EG) nr 2099/2002
av den 5 november 2002
om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS) och om ändring av förordningarna om sjösäkerhet och förhindrande av förorening från fartyg
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
med beaktande av Regionkommitténs yttrande(3),
i enlighet med förfarandet i artikel 251 i fördraget(4), och
av följande skäl:
(1) Genomförandeåtgärderna i gällande förordningar och direktiv inom sjösäkerhetsområdet har antagits genom ett föreskrivande förfarande inom ramen för den kommitté som inrättas genom rådets direktiv 93/75/EEG av den 13 september 1993 om minimikrav för fartyg som anlöper eller avgår från gemenskapens hamnar med farligt eller förorenande gods(5) och i vissa fall en ad hoc-kommitté. Dessa kommittéer har styrts av reglerna i rådets beslut 87/373/EEG av den 13 juli 1987 om närmare villkor för utövandet av kommissionens genomförandebefogenheter(6).
(2) I sin resolution av den 8 juni 1993 om en gemensam politik för säkerhet till sjöss(7) godkände rådet i princip att det inrättas en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS) och uppmanade kommissionen att lägga fram ett förslag om att inrätta en sådan kommitté.
(3) COSS roll består av att centralisera uppgifterna för de kommittéer som inrättats enligt gemenskapslagstiftningen om sjösäkerhet, förhindrande av förorening från fartyg och skydd av boende- och arbetsförhållanden ombord på fartyg samt att bistå och ge kommissionen råd i alla frågor som rör sjösäkerhet och förebyggande eller minskning av miljöföroreningar från sjöfartsverksamhet.
(4) I enlighet med resolutionen av den 8 juni 1993 bör en kommitté för sjösäkerhet och förhindrande av förorening från fartyg inrättas och tilldelas de uppgifter som tidigare hört till de kommittéer som inrättats inom ramen för nämnda lagstiftning. All ny gemenskapslagstiftning som antas inom sjösäkerhetsområdet bör innehålla hänvisning till denna kommitté.
(5) Beslut 87/373/EEG har ersatts med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(8), vars bestämmelser bör tillämpas på COSS. Syftet med beslut 1999/468/EG är att fastställa tillämpliga kommittéförfaranden och att garantera mer uttömmande information till Europaparlamentet och allmänheten om kommittéernas arbete.
(6) De åtgärder som behövs för att genomföra nämnda lagstiftning bör antas i enlighet med beslut 1999/468/EG.
(7) Nämnda lagstiftning bör också ändras så att COSS ersätter den kommitté som inrättats genom direktiv 93/75/EEG eller, i förekommande fall, den ad hoc-kommitté som inrättas genom en viss rättsakt. Genom denna förordning bör framför allt relevanta bestämmelser i rådets förordningar (EEG) nr 613/91 av den 4 mars 1991 om överflyttning av fartyg från ett register till ett annat inom gemenskapen(9), (EG) nr 2978/94 av den 21 november 1994 om genomförande av IMO-resolution A.747(18) om tillämpningen av mätning av dräktighet av barlastutrymmen i oljetankfartyg med segregerade barlasttankar(10) och (EG) nr 3051/95 av den 8 december 1995 om säkerhetsorganisation för roll-on/roll-off-passagerarfartyg (ro-ro-fartyg)(11) samt Europaparlamentets och rådets förordning (EG) nr 417/2002 av den 18 februari 2002 om ett påskyndat införande av krav på dubbelskrov eller likvärdig konstruktion för oljetankfartyg med enkelskrov och om upphävande av rådets förordning (EG) nr 2978/94(12) ändras för infogande av en hänvisning till COSS och för tillämpning av det föreskrivande förfarande som anges i artikel 5 i beslut 1999/468/EG.
(8) Nämnda lagstiftning grundar sig på tillämpningen av regler som härrör från sådana internationella instrument som är i kraft vid tidpunkten för antagandet av den aktuella gemenskapsrättsakten eller vid en tidpunkt som anges i denna. Detta innebär att medlemsstaterna inte kan tillämpa senare ändringar av dessa internationella instrument, om inte gemenskapens direktiv eller förordningar ändras. Svårigheten att få tidpunkten för ikraftträdandet av ändringen på internationell nivå att sammanfalla med tidpunkten för ikraftträdandet av den förordning genom vilken ändringen infogas i gemenskapsrätten orsakar stora problem, och framför allt försenas tillämpningen av nyare och strängare internationella säkerhetsnormer inom gemenskapen.
(9) Skillnad måste emellertid göras mellan sådana bestämmelser i en gemenskapsrättsakt för vilkas tillämpning det hänvisas till ett internationellt instrument och sådana gemenskapsbestämmelser som ordagrant återger ett internationellt instrument helt eller delvis. I det sistnämnda fallet kan de senaste ändringarna av internationella instrument ändå inte tillämpas på gemenskapsnivå förrän de berörda gemenskapsbestämmelserna har ändrats.
(10) Medlemsstaterna bör därför tillåtas att tillämpa de senaste bestämmelserna i de internationella instrumenten, med undantag för bestämmelser som redan uttryckligen ingår i en gemenskapsrättsakt. Detta kan uppnås genom att man anger att den version av den internationella konvention som skall beaktas för det berörda direktivet eller den berörda förordningen skall vara "i gällande version", utan att ett datum anges.
(11) För insynens skull bör relevanta ändringar av de internationella instrument som är införlivade i gemenskapens sjöfartslagstiftning offentliggöras i gemenskapen genom Europeiska gemenskapernas officiella tidning.
(12) Ett särskilt förfarande för kontroll av överensstämmelse bör dock införas, så att kommissionen, efter samråd med COSS, kan vidta nödvändiga åtgärder för att undvika att ändringar av internationella instrument blir oförenliga med nämnda gällande lagstiftning eller gemenskapspolitik på områdena sjösäkerhet, förhindrande av förorening från fartyg samt skydd av boende- och arbetsförhållanden ombord på fartyg, eller med de mål som eftersträvas i denna lagstiftning. Ett sådant förfarande bör även göra det möjligt att förhindra att internationella ändringar försämrar den sjösäkerhet som uppnåtts inom gemenskapen.
(13) Förfarandet för kontroll av överensstämmelse kommer att få full verkan endast om de planerade åtgärderna antas så snart som möjligt, och under alla omständigheter innan den internationella ändringen träder i kraft. Följaktligen bör den tidsfrist som rådet enligt artikel 5.6 i beslut 1999/468/EG beviljas för att fatta beslut om förslag till åtgärder vara en månad.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte
Syftet med denna förordning är att förbättra genomförandet av den gemenskapslagstiftning som avses i artikel 2.2 om sjösäkerhet, förhindrande av förorening från fartyg samt boende- och arbetsförhållanden ombord på fartyg genom att
a) centralisera uppgifterna för de kommittéer som inrättats enligt gemenskapens sjöfartslagstiftning och som upphävs genom denna förordning, genom inrättande av en enda kommitté för sjösäkerhet och förhindrande av förorening från fartyg, kallad COSS,
b) påskynda uppdateringen och underlätta senare ändringar av gemenskapens sjöfartslagstiftning mot bakgrund av utvecklingen av de internationella instrument som avses i artikel 2.1.
Artikel 2
Definitioner
2. gemenskapens sjöfartslagstiftning: följande gällande gemenskapsrättsakter:
a) Rådets förordning (EEG) nr 613/91.
b) Rådets direktiv 93/75/EEG.
c) Rådets förordning (EG) nr 2978/94.
d) Rådets direktiv 94/57/EG av den 22 november 1994 om gemensamma regler och standarder för organisationer som utför inspektioner och utövar tillsyn av fartyg och för sjöfartsadministrationernas verksamhet i förbindelse därmed.(13)
e) Rådets direktiv 95/21/EG av den 19 juni 1995 om hamnstatskontroll.(14)
f) Rådets förordning (EG) nr 3051/95.
g) Rådets direktiv 96/98/EG av den 20 december 1996 om marin utrustning.(15)
h) Rådets direktiv 97/70/EG av den 11 december 1997 om att införa harmoniserade säkerhetsregler för fiskefartyg som har en längd av 24 meter och däröver.(16)
i) Rådets direktiv 98/18/EG av den 17 mars 1998 om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg.(17)
j) Rådets direktiv nr 98/41/EG av den 18 juni 1998 om registrering av personer som färdas ombord på passagerarfartyg som ankommer till eller avgår från hamnar i gemenskapens medlemsstater.(18)
k) Rådets direktiv 1999/35/EG av den 29 april 1999 om ett system med obligatoriska besiktningar för en säker drift av ro-ro-passagerarfartyg och höghastighetspassagerarfartyg i reguljär trafik.(19)
l) Europaparlamentets och rådets direktiv 2000/59/EG av den 27 november 2000 om mottagningsanordningar i hamn för fartygsgenererat avfall och lastrester.(20)
m) Europaparlamentets och rådets direktiv 2001/25/EG av den 4 april 2001 om minimikrav på utbildning för sjöfolk.(21)
n) Europaparlamentets och rådets direktiv 2001/96/EG av den 4 december 2001 om fastställande av harmoniserade krav och förfaranden för säker lastning och lossning av bulkfartyg.(22)
o) Europaparlamentets och rådets förordning (EG) nr 417/2002.
Artikel 3
Inrättande av en kommitté
1. Kommissionen skall biträdas av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg, nedan kallad COSS.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara en månad.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 4
Genomförande i gemenskapens lagstiftning av ändringar av internationella instrument
Gemenskapens sjöfartslagstiftning skall omfattas av de internationella instrument som har trätt i kraft, inbegripet de senaste ändringarna av dessa, med undantag för de ändringar som undantagits från tillämpningsområdet för gemenskapens sjöfartslagstiftning på grund av resultatet av det förfarande för kontroll av överensstämmelse som fastställs i artikel 5.
Artikel 5
Förfarande för kontroll av överensstämmelse
1. För att uppnå syftet med denna förordning och för att minska risken för en konflikt mellan gemenskapens sjöfartslagstiftning och internationella instrument skall medlemsstaterna och kommissionen samarbeta genom samordningsmöten och/eller på andra lämpliga sätt för att i förekommande fall fastställa en gemensam ståndpunkt eller strategi i behöriga internationella forum.
2. Ett förfarande för kontroll av överensstämmelse inrättas härmed i syfte att från tillämpningsområdet för gemenskapens sjöfartslagstiftning undanta en ändring av ett internationellt instrument endast om det, på grundval av en bedömning från kommissionens sida, finns en uppenbar risk att den internationella ändringen, inom ramen för tillämpningsområdet för de förordningar eller direktiv som avses i artikel 2.2, kommer att försämra den nivå på sjösäkerheten, förhindrandet av förorening från fartyg eller skydd av boende- och arbetsförhållandena ombord på fartyg som fastställs i gemenskapens sjöfartslagstiftning, eller vara oförenlig med denna lagstiftning.
Förfarandet för kontroll av överensstämmelse får användas enbart för att ändra gemenskapens sjöfartslagstiftning på de områden som uttryckligen omfattas av det föreskrivande förfarandet och strikt inom ramen för kommissionens genomförandebefogenheter.
3. Om det föreligger sådana omständigheter som avses i punkt 2 skall förfarandet för kontroll av överensstämmelse inledas av kommissionen, eventuellt på begäran av någon medlemsstat.
Kommissionen skall snarast efter antagandet av en ändring av ett internationellt instrument för COSS lägga fram ett förslag till åtgärder som syftar till att undanta den aktuella ändringen från den gemenskapstext som berörs.
Förfarandet för kontroll av överensstämmelse, i förekommande fall inbegripet förfarandena enligt artikel 5.6 i beslut 1999/468/EG, skall slutföras senast en månad innan den period löper ut som fastställts internationellt för underförstått godkännande av ändringen i fråga eller senast en månad före den planerade tidpunkten för ändringens ikraftträdande.
4. Om en sådan risk som avses i punkt 2 första stycket föreligger skall medlemsstaterna under förfarandet för kontroll av överensstämmelse avhålla sig från varje initiativ som syftar till att genomföra ändringen i den nationella lagstiftningen eller tillämpa denna ändring av det internationella instrumentet i fråga.
Artikel 6
Information
Alla relevanta ändringar av de internationella instrument som är införlivade i gemenskapens sjöfartslagstiftning i enlighet med artiklarna 4 och 5 skall i informationssyfte offentliggöras i Europeiska gemenskapernas officiella tidning.
Artikel 7
COSS befogenheter
COSS skall utöva de befogenheter som den tilldelas i enlighet med gällande gemenskapslagstiftning. Artikel 2.2 får ändras genom det förfarande som anges i artikel 3.2 i syfte att infoga en hänvisning till gemenskapsrättsakter som trätt i kraft efter antagandet av denna förordning och enligt vilka COSS tillerkänns genomförandebefogenheter.
Artikel 8
Ändring av förordning (EEG) nr 613/91
Förordning (EEG) nr 613/91 ändras på följande sätt:
1. Artikel 1 a skall ersättas med följande:
"a) Konventioner: 1974 års internationella konvention om säkerheten för människoliv till sjöss (Solas 1974), 1996 års internationella lastlinjekonvention (LL 66) och den internationella konventionen om förhindrande av förorening från fartyg (Marpol 73/78), i gällande version, och tillhörande bindande resolutioner, som har antagits av Internationella sjöfartsorganisationen (IMO)."
2. Artiklarna 6 och 7 skall ersättas med följande:
"Artikel 6
1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i Europaparlamentets och rådets förordning (EG) nr 2099/2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(23).
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(24) tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara två månader.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 7
Ändringarna av de internationella instrument som avses i artikel 1 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i förordning (EG) nr 2099/2002."
Artikel 9
Ändring av förordning (EG) nr 2978/94
Förordning (EG) nr 2978/94 ändras på följande sätt:
1. Artikel 3 g skall ersättas med följande:
"g) Marpol 73/78: 1973 års internationella konvention till förhindrande av förorening från fartyg, i dess lydelse enligt det därtill hörande protokollet av år 1978, i gällande version."
2. Följande stycke skall läggas till i artikel 6:"Ändringarna av de internationella instrument som avses i artikel 3 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i Europaparlamentets och rådets förordning (EG) nr 2099/2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(25)."
3. Artikel 7 skall ersättas med följande:
"Artikel 7
1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i förordning (EG) nr 2099/2002.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(26) tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning."
Artikel 10
Ändring av förordning (EG) nr 3051/95
Förordning (EG) nr 3051/95 ändras på följande sätt:
1. Följande stycke skall läggas till i artikel 9:"Ändringarna av de internationella instrument som avses i artikel 2 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i Europaparlamentets och rådets förordning (EG) nr.../2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(27)."
2. Artikel 10 skall ersättas med följande:
"Artikel 10
1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i förordning (EG) nr 2099/2002.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(28) tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara två månader.
3. Kommittén skall själv anta sin arbetsordning."
Artikel 11
Ändring av förordning (EG) nr 417/2002
Förordning (EG) nr 417/2002 ändras på följande sätt:
2. Artikel 10.1 skall ersättas med följande:
"1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i Europaparlamentets och rådets förordning (EG) nr 2099/2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(29)."
3. Följande stycke läggas till i artikel 11:"Ändringarna av de internationella instrument som avses i artikel 3.1 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i förordning (EG) nr 2099/2002."
Artikel 12
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2104/2002
av den 28 november 2002
om anpassning av rådets förordning (EG) nr 577/98 om anordnande av statistiska urvalsundersökningar av arbetskraften i gemenskapen och kommissionens förordning (EG) nr 1575/2000 om genomförande av rådets förordning (EG) nr 577/98 vad gäller förteckningen över variabler för utbildning samt deras kodning för användning vid överföring av data från och med 2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 577/98 av den 9 mars 1998 om anordnande av statistiska urvalsundersökningar av arbetskraften i gemenskapen(1), ändrad genom Europarlamentets och rådets förordning (EG) nr 1991/2002(2), särskilt artikel 4.3 i denna, och
av följande skäl:
(1) Utvecklingen av tekniker och begrepp, i synnerhet vad gäller skillnaden mellan formell utbildning och andra former av undervisningsaktiviteter och genomförandet av klassificeringen av inriktningen av utbildningen, framtvingar en anpassning av förteckningen över variabler för utbildning som anges i artikel 4.1 h i förordning (EG) nr 577/98.
(2) Härav följer att koderna för dessa variabler enligt vad som anges i bilagan till kommissionens förordning (EG) nr 1575/2000 av den 19 juli 2000(3) också skall anpassas. Den nya förteckningen och kodningen skall genomföras redan under 2003 så att full kompatibilitet med ad hoc-modulen för 2003 om livslångt lärande(4) kan garanteras.
(3) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från kommittén för det statistiska programmet, inrättad genom rådets beslut 89/382/EEG, Euratom(5).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 4.1 h i rådets förordning (EG) nr 577/98 skall ersättas med följande:
"h) Utbildning
deltagande i formell utbildning under de närmast föregående fyra veckorna
- nivå
- inriktning
deltagande i kurser och annan undervisningsaktivitet under de närmast föregående fyra veckorna
- total längd
- syfte för de senaste kurserna eller annan undervisningsaktivitet
- inriktning på den senaste undervisningsaktiviteten
- om den senaste undervisningsaktiviteten skett på arbetstid
utbildningsnivå
- högsta nivå för med framgång avslutad utbildning
- inriktning för denna högsta nivå av utbildning
- år då denna utbildning framgångsrikt avslutades"
Artikel 2
Koderna för de variabler för utbildning som skall användas för överföring av data under 2003 och framgent som anges i bilagan till denna förordning, ersätter motsvarande variabler i bilagan till kommissionens förordning (EG) nr 1575/2000.
Artikel 3
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens beslut
av den 23 december 2002
om tillämpning av rådets förordning (EEG) nr 1612/68 med avseende på förmedling av lediga platser och platsansökningar
(Text av betydelse för EES)
(2003/8/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1612/68 av den 15 oktober 1968 om arbetskraftens fria rörlighet inom gemenskapen(1), senast ändrad genom förordning (EEG) nr 2434/92(2), särskilt artikel 44 i denna, och
av följande skäl:
(1) Många framsteg har gjorts sedan nätverket för europeiska arbetsförmedlingar (EURES-nätverket) inrättades genom kommissionens beslut 93/569/EEG(3) om genomförandet av rådets förordning (EEG) nr 1612/68.
(2) Mot bakgrund av erfarenheterna sedan 1993 och för att beakta och befästa den nya utvecklingen av EURES-verksamheten, bör nätverket nu stärkas och fullt ut integreras i medlemsstaternas arbetsförmedlingsverksamhet. Den nuvarande ansvarsfördelningen och de nuvarande beslutsförfarandena bör få en ny utformning.
(3) Med hänsyn till den kommande utvidgningen av Europeiska unionen bör införandet av EURES-nätverket i kandidatländerna beaktas i full utsträckning samtidigt som man ser till att systemet fortfarande är effektivt och hanterbart.
(4) De möjligheter som ny informations- och kommunikationsteknik ger att ytterligare förbättra och rationalisera de tjänster som erbjuds bör också beaktas.
(5) EURES-nätverket bör därför befästas och stärkas som ett viktigt instrument för att övervaka den transnationella rörligheten, stödja arbetstagarnas fria rörlighet, integrera de europeiska arbetsmarknaderna och informera medborgarna om relevant gemenskapslagstiftning.
(6) Den yrkesmässiga och geografiska rörligheten behöver stimuleras i enlighet med den europeiska sysselsättningsstrategin med sikte på att genomföra handlingsplanen för kompetens och rörlighet(4) och rådets resolution av den 3 juni 2002 i samma fråga(5).
(7) För tydlighetens skull är det lämpligt att återupprätta EURES-nätverket och samtidigt tydligare fastställa dess sammansättning, uppbyggnad och funktioner. Detta innebär att beslut 93/569/EEG bör ersättas.
(8) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Tekniska kommittén för fri rörlighet för arbetstagare.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
EURES-nätverket
Kommissionen, medlemsstaternas arbetsförmedlingar och övriga nationella partner som de kan ha skall upprätta ett europeiskt nätverk för arbetsförmedlingar, som skall betecknas "EURES-nätverket" (EURopean Employment Services) och ansvara för utvecklingen av det informationsutbyte och samarbete som föreskrivs i del II i förordning (EEG) nr 1612/68.
Artikel 2
Mål
EURES-nätverket skall bidra till en samordnad tillämpning av bestämmelserna i del II i förordning (EEG) nr 1612/68. Nätverket skall stödja den europeiska sysselsättningsstrategin och bidra till att stärka EU:s gemensamma marknad.
EURES-nätverket skall särskilt till förmån för arbetssökande, arbetstagare och arbetsgivare sträva efter att främja
a) utveckling av europeiska arbetsmarknader som är öppna och tillgängliga för alla,
b) förmedling av lediga platser och platsansökningar mellan olika länder och regioner och i gränstrakter,
c) öppenhet och utbyte av information om europeiska arbetsmarknader, inklusive om levnadsvillkor och utbildningsmöjligheter,
d) utveckling av metoder och indikatorer för detta ändamål.
Artikel 3
Sammansättning
EURES-nätverket skall omfatta följande parter:
a) EURES-medlemmar, som skall vara särskilda förmedlingar som medlemsstaterna utser enligt artikel 13.2 i förordning (EEG) nr 1612/68, och Europeiska samordningsbyrån, enligt artiklarna 21, 22 och 23 i den förordningen, och
b) EURES samarbetspartner, enligt artikel 17.1 i förordning (EEG) nr 1612/68, dvs.
i) regionala arbetsförmedlingar i medlemsstaterna,
ii) arbetsförmedlingar som ansvarar för gränstrakter,
iii) särskilda arbetsförmedlingar som anmälts till kommissionen enligt artikel 17.2 i förordning (EEG) nr 1612/68.
Dessa parter skall inbegripa de fackliga organisationer och arbetsgivarorganisationer som EURES medlemmar utser.
Artikel 4
Europeiska samordningsbyråns roll
Kommissionens generaldirektorat för sysselsättning och socialpolitik skall ansvara för Europeiska samordningsbyrån.
Europeiska samordningsbyrån (nedan kallad "EURES samordningsbyrå") skall övervaka iakttagandet av bestämmelserna i del II i förordning (EEG) nr 1612/68 och hjälpa nätverket att genomföra sin verksamhet.
EURES samordningsbyrå skall särskilt
a) analysera den geografiska och yrkesmässiga rörligheten och utarbeta en generell metod för transnationell rörlighet i enlighet med den europeiska sysselsättningsstrategin,
b) utforma en samstämmig och övergripande metod samt lämpliga former för att främja samarbete och samordning mellan medlemsstaterna,
c) ansvara för den övergripande övervakningen och utvärderingen av EURES-verksamheten och vidta åtgärder för att kontrollera att den genomförs enligt bestämmelserna i förordning (EEG) nr 1612/68 och i det här beslutet.
Artikel 5
EURES-logotypen
Akronymen EURES får användas endast för verksamhet inom EURES-nätverket. Den skall illustreras med en logotyp som är definierad i ett grafiskt dokument.
Logotypen skall registreras som ett gemenskapsvarumärke vid Byrån för harmonisering inom den inre marknaden (varumärken och formgivning). Den får användas av EURES medlemmar och samarbetspartner.
Artikel 6
Högnivågrupp för strategiska frågor
En högnivågrupp för strategiska frågor inrättas härmed. Gruppen skall bestå av cheferna för EURES-medlemmarna och ha en företrädare för kommissionen som ordförande. Den skall bistå kommissionen med att främja och övervaka utvecklingen av EURES-nätverket.
Kommissionen skall samråda med högnivågruppen i frågor som rör strategisk planering, utveckling, genomförande, övervakning och utvärdering när det gäller de tjänster och verksamheter som avses i det här beslutet, inklusive
a) EURES-stadgan, enligt artikel 8.2,
b) EURES-nätverkets riktlinjer, enligt artikel 9.1,
c) kommissionens utkast till årsrapport som föreskrivs enligt artikel 19.1 i förordning (EEG) nr 1612/68,
d) den rapport som kommissionen vartannat år skall lämna till Europaparlamentet, rådet och Europeiska ekonomiska och sociala kommittén enligt artikel 19.3 i förordning (EEG) nr 1612/68.
Ledarna för arbetsmarknadsorganisationerna på EU-nivå skall inbjudas till att delta i gruppens möten.
Gruppen skall själv fastställa sina arbetsmetoder och anta sin arbetsordning. Gruppen skall sammankallas av ordföranden minst två gånger per år. Den skall anta sina yttranden med enkel majoritet.
EURES samordningsbyrå skall ställa sekreterartjänster till förfogande.
Artikel 7
Arbetsgrupp
För att bistå högnivågruppen med utvecklingen, genomförandet och övervakningen av EURES-verksamheten skall EURES samordningsbyrå inrätta en arbetsgrupp som består av EURES-ansvariga ("EURES-managers"), som var och en företräder en EURES-medlem. EURES samordningsbyrå skall bjuda in företrädare för arbetsmarknadens parter på EU-nivå och, i lämpliga fall, företrädare för andra samarbetspartner och experter inom EURES att delta i arbetsgruppens möten.
Artikel 8
EURES-stadga
1. EURES samordningsbyrå skall anta EURES-stadgan enligt de förfaranden som anges i artiklarna 14.2 och 15.2, artikel 22.1 a, b och c samt artikel 23 i förordning (EEG) nr 1612/68, efter samråd med den högnivågrupp för strategiska frågor som inrättas genom artikel 6 i det här beslutet.
2. Utifrån principen om att alla lediga platser och platsansökningar som offentliggörs av EURES medlemmar och samarbetspartner skall göras tillgängliga i hela Europeiska gemenskapen, skall EURES-stadgan särskilt innehålla följande information:
a) Beskrivningar av den verksamhet som EURES medlemmar och samarbetspartner skall bedriva, vilket inbegriper
i) arbetsförmedling, inklusive personlig vägledning och rådgivning till kunder, antingen de är arbetssökande, arbetstagare eller arbetsgivare,
ii) utveckling av samarbetet mellan olika länder och i gränstrakter, inklusive arbetsförmedling och social service, arbetsmarknadens parter och andra institutioner som berörs, med sikte på att arbetsmarknaderna skall fungera bättre och integreras samt på att öka rörligheten,
iii) främjande av en samordnad övervakning och bedömning av hinder för rörligheten, överskott och brist på kunskaper samt migrationsströmmar.
b) Verksamhetsmål för EURES-systemet, de kvalitetskrav som skall gälla samt EURES medlemmars och samarbetspartners skyldigheter, vilket inbegriper
i) integrering av medlemmarnas databaser för lediga platser i EURES-systemet för förmedling av lediga platser inom en tidsfrist som skall bestämmas,
ii) typ av information, t.ex. information om arbetsmarknaden, levnad- och arbetsvillkor, lediga platser och platsansökningar samt hinder för rörlighet, som de måste lämna till sina kunder och till nätverket,
iii) utbildning och kvalifikationer som krävs av EURES-personal samt villkor och förfaringssätt för att organisera besök och uppdrag för tjänstemän,
iv) utarbetande, inlämnande till EURES samordningsbyrå och genomförande av verksamhetsplaner, med särskilda regler för EURES-verksamhet som bedrivs över gränserna,
v) villkor för användning av EURES-logotypen för medlemmar och samarbetspartner,
vi) principer för övervakning och utvärdering av EURES-verksamheten.
c) Förfaranden för att upprätta ett enhetligt system och gemensamma former för utbyte av information om arbetsmarknaden och om transnationell rörlighet inom EURES-nätverket, i enlighet med artiklarna 14, 15 och 16 i förordning (EEG) nr 1612/68, inklusive information om lediga platser och utbildningsmöjligheter inom Europeiska unionen som skall integreras i en webbplats för information om rörlighet i arbetslivet.
Artikel 9
Riktlinjer och verksamhetsplaner
1. I enlighet med den EURES-stadga som föreskrivs i artikel 8 och efter samråd med den högnivågrupp för strategiska frågor som avses i artikel 6, skall EURES samordningsbyrå fastställa riktlinjer för EURES-verksamheten för en period på tre år.
I riktlinjerna skall villkoren för det ekonomiska stöd som Europeiska gemenskapen kan lämna i enlighet med punkt 4 anges.
2. Utifrån dessa riktlinjer skall EURES-medlemmarna lämna sina verksamhetsplaner för den period som riktlinjerna omfattar till EURES samordningsbyrå. Verksamhetsplanerna skall innehålla uppgifter om
a) den huvudsakliga verksamhet som EURES-medlemmen skall bedriva inom ramen för nätverket, inklusive sådan transnationell, gränsöverskridande och branschspecifik verksamhet som avses i artikel 17 i förordning (EEG) nr 1612/68,
b) den personal och de ekonomiska resurser som tilldelats för tillämpningen av del II i förordning (EEG) nr 1612/68,
c) formerna för övervakning och utvärdering av den planerade verksamheten, inklusive den information som skall lämnas till kommissionen varje år.
Verksamhetsplanerna skall även innehålla en utvärdering av verksamheten och de framsteg som gjorts under den föregående perioden.
3. EURES samordningsbyrå skall granska verksamhetsplanerna och den information som lämnats om deras genomförande för att bedöma om de följer riktlinjerna och bestämmelserna i del II i förordning (EEG) nr 1612/68. Resultaten av denna bedömning skall granskas tillsammans med EURES-medlemmarna varje år i enlighet med artikel 19.1 i den förordningen samt inbegripas i den rapport som kommissionen vartannat år skall lämna till Europaparlamentet, rådet och Ekonomiska och sociala kommittén i enlighet med artikel 19.3 i den förordningen.
4. Kommissionen får bevilja ekonomiskt stöd för genomförandet av verksamhetsplanerna i enlighet med bestämmelserna om de relevanta budgetmedlen.
Artikel 10
Upphävande
Beslut 93/569/EEG upphävs härmed. Det skall dock fortsätta att tillämpas på verksamhet för vilken en ansökan hade lämnats in innan det här beslutet trädde i kraft.
Artikel 11
Datum för tillämpning
Detta beslut skall tillämpas från och med den 1 mars 2003.
Artikel 12
Adressater
Detta beslut riktar sig till medlemsstaterna.
Europaparlamentets och rådets direktiv 2003/24/EG
av den 14 april 2003
om ändring av rådets direktiv 98/18/EG om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Genom rådets direktiv 98/18/EG av den 17 mars 1998 om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg(4) införs en enhetlig säkerhetsnivå för människoliv och egendom på nya och existerande passagerarfartyg och höghastighetspassagerarfartyg när dessa typer av fartyg används på inrikes resor, och fastställs förfaranden för förhandlingar på internationell nivå i syfte att harmonisera bestämmelserna för passagerarfartyg som används på internationella resor.
(2) Definitionen av fartområden är avgörande för hur direktiv 98/18/EG skall tillämpas på olika passagerarfartygsklasser. Direktivet innehåller ett förfarande för offentliggörandet av förteckningar av fartområden som visat sig vara svårt att genomföra. Det är därför nödvändigt att skapa ett praktiskt genomförbart och öppet förfarande som möjliggör en effektiv övervakning av direktivets genomförande.
(3) I syfte att harmonisera säkerhetsnivån för passagerarfartyg i hela gemenskapen bör det undantag som beviljats Grekland när det gäller tidtabellen för tillämpningen av säkerhetsbestämmelserna upphävas.
(4) Genom Europaparlamentets och rådets direktiv 2003/25/EG av den 14 april 2003 om särskilda stabilitetskrav för ro-ro-passagerarfartyg(5) införs skärpta stabilitetskrav för ro-ro-passagerarfartyg som går i internationell trafik till och från hamnar i gemenskapen; dessa krav bör även omfatta vissa kategorier av fartyg som går i inrikes trafik under motsvarande sjöförhållanden. Ro-ro-passagerarfartyg som inte uppfyller dessa stabilitetskrav bör tas ur trafik efter ett visst antal år i drift.
(5) Med tanke på de ombyggnader av existerande ro-ro-passagerarfartyg som kan vara nödvändiga för att de skall uppfylla de särskilda stabilitetskraven, bör dessa krav införas successivt under ett antal år, så att den del av branschen som berörs får tillräcklig tid att uppfylla kraven. En tidtabell för infasning av existerande fartyg bör därför fastställas. Denna tidtabell för infasning bör inte påverka tillämpningen av de särskilda stabilitetskraven i de fartområden som omfattas av bilagorna till Stockholmsöverenskommelsen av den 28 februari 1996.
(6) Ändringar i relevanta internationella texter, t.ex. Internationella sjöfartsorganisationens (IMO) konventioner, protokoll, koder och resolutioner, måste kunna beaktas på ett flexibelt och snabbt sätt.
(7) Enligt direktiv 98/18/EG är den internationella säkerhetskoden för höghastighetsfartyg - fastställd i IMO:s sjösäkerhetskommittés resolution MSC 36 (63) av den 20 maj 1994 - tillämplig på alla höghastighetspassagerarfartyg som går i inrikes trafik. IMO har antagit en ny kod för höghastighetsfartyg - Internationella säkerhetskoden för höghastighetsfartyg 2000 (HSC-koden 2000), fastställd i IMO:s sjösäkerhetskommittés resolution MSC 97 (73) av den 5 december 2000 - som är tillämplig på alla höghastighetsfartyg byggda den 1 juli 2002 eller senare. Det är viktigt att se till att direktiv 98/18/EG kan uppdateras på ett flexibelt sätt så att sådan utveckling på internationell nivå kan tillämpas, även på höghastighetspassagerarfartyg som går i inrikes trafik.
(8) Det är viktigt att vidta lämpliga åtgärder för att garantera att personer med nedsatt rörlighet under säkra former kan ta sig ombord på passagerarfartyg och höghastighetspassagerarfartyg i inrikes trafik i medlemsstaterna.
(9) Direktiv 98/18/EG bör därför ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 98/18/EG ändras enligt följande:
1. I artikel 2 skall följande punkter läggas till:
"ea) ro-ro-passagerarfartyg: ett fartyg som medför fler än tolv passagerare och som har ro-ro-lastutrymmen eller lastutrymmen av särskild kategori enligt definitionen i regel II-2/A/2 i bilaga I."
"ha) ålder: fartygets ålder uttryckt i antal år efter dess leveransdatum."
"w) personer med nedsatt rörlighet: alla personer som har särskilda problem med att använda allmänna transportmedel, inbegripet äldre, personer med funktionshinder, personer med sensoriska funktionshinder och rullstolsburna, gravida, och personer i sällskap med små barn."
2. I artikel 4 skall punkt 2 ersättas med följande:
"2. Varje medlemsstat skall
a) fastställa och vid behov uppdatera en förteckning över de fartområden som omfattas av deras jurisdiktion och fastställa zonerna för åretrunttrafik och, i förekommande fall, begränsad periodisk trafik för de olika fartygsklasserna enligt klassificeringskriterierna i punkt 1,
b) offentliggöra förteckningen i en offentlig databas som är tillgänglig på den behöriga sjöfartsmyndighetens webbplats på Internet, och
c) till kommissionen anmäla var denna information finns och när förteckningen senast ändrades.".
3. Följande artiklar skall införas:
"Artikel 6a
Stabilitetskrav för och utfasning av ro-ro-passagerarfartyg
1. Ro-ro-passagerarfartyg i klasserna A-C som kölsträcks eller är på motsvarande byggnadsstadium den 1 oktober 2004 eller senare skall uppfylla artiklarna 6, 8 och 9 i Europaparlamentets och rådets direktiv 2003/25/EG av den 14 april 2003 om särskilda stabilitetskrav för ro-ro-passagerarfartyg(6).
2. Ro-ro-passagerarfartyg i klasserna A och B som kölsträcks eller är på motsvarande byggnadsstadium före den 1 oktober 2004 skall uppfylla artiklarna 6, 8 och 9 i direktiv 2003/25/EG före den 1 oktober 2010 såvida de inte har tagits ur trafik den dagen eller vid en senare tidpunkt vid vilken de har uppnått en ålder av 30 år, dock senast den 1 oktober 2015.
Artikel 6b
Säkerhetskrav för personer med nedsatt rörlighet
1. Medlemsstaterna skall se till att lämpliga åtgärder vidtas, när så är praktiskt möjligt på grundval av riktlinjerna i bilaga III, för att passagerare med nedsatt rörlighet skall kunna ta sig ombord under säkra former på alla passagerarfartyg i klasserna A-D och alla höghastighetspassagerarfartyg som används för allmänna transporter och som kölsträcks eller befinner sig på motsvarande byggnadsstadium den 1 oktober 2004 eller senare.
2. Medlemsstaterna skall samarbeta och samråda med organisationer som företräder personer med nedsatt rörlighet när det gäller genomförandet av riktlinjerna i bilaga III.
3. När det gäller ombyggnaden av passagerarfartyg i klasserna A-D och höghastighetspassagerarfartyg som används för allmänna transporter och som kölsträcks eller befinner sig på motsvarande byggnadsstadium före den 1 oktober 2004, skall medlemsstaterna tillämpa riktlinjerna i bilaga III, i den mån det är rimligt och praktiskt möjligt i ekonomiskt hänseende.
Medlemsstaterna skall utarbeta nationella handlingsplaner för hur riktlinjerna skall tillämpas på sådana fartyg. Medlemsstaterna skall till kommissionen översända dessa handlingsplaner senast den 17 maj 2005.
4. Medlemsstaterna skall senast den 17 maj 2006 rapportera till kommissionen om genomförandet av denna artikel beträffande alla passagerarfartyg som avses i punkt 1, de passagerarfartyg som avses i punkt 3 och som är certifierade för fler än 400 passagerare samt alla höghastighetspassagerarfartyg."
4. Bilagan till detta direktiv skall läggas till som bilaga III.
Artikel 2
Artikel 6.3 g i direktiv 98/18/EG skall utgå med verkan från och med den 1 januari 2005.
Artikel 3
Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 17 november 2004. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 4
Kommissionens direktiv 2003/26/EG
av den 3 april 2003
om anpassning till den tekniska utvecklingen av Europaparlamentets och rådets direktiv 2000/30/EG i fråga om hastighetsbegränsande anordningar och avgasutsläpp från nyttofordon
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets direktiv 2000/30/EG av den 6 juni 2000 om vägkontroller av trafiksäkerheten hos nyttofordon i trafik i gemenskapen(1), särskilt artikel 8 i detta, och
av följande skäl:
(1) Direktiv 2000/30/EG rör den rättsliga ram för vägkontroller av nyttofordon, oavsett om de fraktar passagerare eller gods. Direktivet innehåller krav på att medlemsstaterna skall komplettera de årliga trafiksäkerhetsprovningarna med oanmälda vägkontroller av en representativ del av nyttofordonen varje år.
(2) Området trafiksäkerhet omfattas av rådets direktiv 96/96/EG av den 20 december 1996 om tillnärmning av medlemsstaternas lagstiftning om provning av motorfordons och tillhörande släpfordons trafiksäkerhet(2), senast ändrat genom kommissionens direktiv 2001/11/EG(3), som omfattar reguljära trafiksäkerhetsprovningar, samt av direktiv 2000/30/EG, som gäller vägkontroller av trafiksäkerheten hos tunga nyttofordon. I bägge direktiven förekommer samma kommitté och förfarande för tekniska anpassningar.
(3) Direktiv 96/96/EG har ändrats genom införande av skärpta utsläppsgränser för vissa kategorier av motorfordon och funktionsprovning av hastighetsbegränsande anordningar på tunga nyttofordon. Direktiv 2000/30/EG bör anpassas för att överensstämma med det direktivet genom att nya tekniska bestämmelser införs om att omborddiagnossystem och hastighetsbegränsande anordningar skall omfattas av vägkontrollerna. För att överensstämma med direktiv 96/96/EG, måste det införas nya tekniska bestämmelser i direktiv 2000/30/EG, vilket skall ske genom att omborddiagnossystem och hastighetsbegränsande anordningar skall omfattas av vägkontrollerna. Direktiv 2000/30/EG bör också uppdateras (tillsammans med direktiv 96/96/EG) så att det innehåller reviderade utsläppsgränsvärdena för vissa kategorier av motorfordon.
(4) De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från den kommitté för anpassning till den tekniska utvecklingen som inrättats genom artikel 8 i direktiv 96/96/EG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagorna I och II till direktiv 2000/30/EG ändras enligt bilagan till detta direktiv.
Artikel 2
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 2004. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 3
Europaparlamentets och rådets direktiv 2003/30/EG
av den 8 maj 2003
om främjande av användningen av biodrivmedel eller andra förnybara drivmedel
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175.1 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande(2),
med beaktande av Regionkommitténs yttrande(3),
i enlighet med förfarandet i artikel 251 i fördraget(4), och
av följande skäl:
(1) Europeiska rådet enades vid mötet i Göteborg den 15 och 16 juni 2001 om en gemenskapsstrategi för hållbar utveckling som omfattar ett antal åtgärder, däribland utvecklingen av biodrivmedel.
(2) Naturresurserna, som enligt artikel 174.1 i fördraget skall utnyttjas varsamt och rationellt, utgörs bland annat av olja, naturgas och fasta bränslen, vilka är viktiga energikällor, men de ger även upphov till de största koldioxidutsläppen.
(3) Det finns dock ett brett spektrum av biomassa som kan användas för att producera biodrivmedel och som härrör från jordbruks- och skogsbruksprodukter liksom från restprodukter och avfall från skogsbruk och skogs- och jordbrukslivsmedelsindustrin.
(4) Transportsektorn, som svarar för mer än 30 % av den slutliga energiförbrukningen i gemenskapen, expanderar och trenden kommer med all säkerhet att förstärkas och koldioxidutsläppen öka; denna expansion kommer att bli procentuellt högre i kandidatländerna efter deras anslutning till Europeiska unionen.
(5) Kommissionen anger i sin vitbok "Den gemensamma transportpolitiken fram till 2010: Vägval inför framtiden" att koldioxidutsläppen från transportsektorn förväntas öka med 50 % mellan 1990 och 2010 till omkring 1113 miljoner ton, varvid vägtransporterna, som svarar för 84 % av de transportrelaterade koldioxidutsläppen, bär det tyngsta ansvaret. I vitboken ställs det därför av miljöskäl upp krav på att oljeberoendet (för närvarande 98 %) inom transportsektorn skall minskas genom användning av alternativa drivmedel, såsom biodrivmedel.
(6) En ökad användning av biodrivmedel utgör en del av det åtgärdspaket som krävs för att följa Kyotoprotokollet, liksom av andra strategier för att uppfylla ytterligare åtaganden i detta hänseende.
(7) En ökad användning av biodrivmedel - utan att för den skulle utesluta användning av andra möjliga alternativa drivmedel, inbegripet motorgas (LPG) och komprimerad naturgas (CNG) för motorfordon - är ett av flera sätt för gemenskapen att minska sitt beroende av importerad energi och påverka drivmedelsmarknaden och således energiförsörjningstryggheten på medellång och lång sikt. Detta bör dock inte på något sätt minska vikten av att gemenskapslagstiftningen om bränslekvalitet, fordonsutsläpp och luftkvalitet efterlevs.
(8) Framsteg i tekniken har lett till att de flesta fordon som i dag är i bruk i Europeiska unionen utan problem kan använda en låg inblandning av biodrivmedel. De senaste tekniska framstegen gör det möjligt att använda högre halter av biodrivmedel i blandningen. I vissa länder används redan blandningar som innehåller halter av biodrivmedel på 10 % och däröver.
(9) Avgränsade fordonsflottor erbjuder möjligheten att använda biodrivmedel i högre koncentration. I vissa städer finns det redan avgränsade fordonsflottor som drivs med rent biodrivmedel, vilket i vissa fall har bidragit till att förbättra luftkvaliteten i städerna. Medlemsstaterna skulle därför ytterligare kunna främja användningen av biodrivmedel i offentliga transportmedel.
(10) Att främja användningen av biodrivmedel utgör ett steg mot en utökad användning av biomassa, vilket gör det möjligt att utveckla biodrivmedlen ytterligare i framtiden samtidigt som andra alternativ inte utesluts, särskilt inte vätgasalternativet.
(11) Medlemsstaternas forskningspolitik om ökad användning av biodrivmedel bör i avsevärd utsträckning omfatta vätgassektorn och främja detta alternativ, och därvid beakta gemenskapens alla relevanta ramprogram.
(12) Ren vegetabilisk olja från oljeväxter som framställs genom pressning, extraktion eller jämförbara metoder, rå eller raffinerad men kemiskt oförändrad, kan också användas som biodrivmedel i vissa fall där användningen är förenlig med motortyperna och motsvarande utsläppskrav.
(13) Nya typer av drivmedel bör uppfylla erkända tekniska standarder för att accepteras i större omfattning av konsumenter och fordonstillverkare, och därmed få spridning på marknaden. Tekniska standarder utgör också utgångspunkten för krav när det gäller utsläpp och övervakning av utsläpp. Nya drivmedelstyper kan ha svårt att uppfylla dagens tekniska standarder, som i stor utsträckning har utvecklats för konventionella fossila drivmedel. Kommissionen och standardiseringsorganen bör övervaka utvecklingen och aktivt anpassa och utveckla standarder, i synnerhet flyktighetsparametrar, så att nya typer av drivmedel kan införas med bibehållna krav på miljöprestanda.
(14) Bioetanol och biodiesel som i ren form eller i blandningar används i fordon bör uppfylla de kvalitetsstandarder som fastställts för att motorerna skall fungera optimalt. Det noteras att Europeiska standardiseringskommitténs standard prEN 14214 för fettsyrametylestrar (FAME) kan tillämpas i fråga om biodiesel för dieselmotorer, där tillverkningsalternativet är omförestring. Europeiska standardiseringskommittén bör sålunda fastställa lämpliga standarder för andra biodrivmedelsprodukter i Europeiska unionen.
(15) Att främja användningen av biodrivmedel i enlighet med hållbara jordbruks- och skogsbruksmetoder som föreskrivs i bestämmelserna inom den gemensamma jordbrukspolitiken kan skapa nya möjligheter till hållbar utveckling av landsbygden inom ramen för en mer marknadsinriktad gemensam jordbrukspolitik som är mer inriktad på den europeiska marknadens behov, en levande landsbygd och ett mångsidigare jordbruk och kan öppna en ny marknad för innovativa jordbruksprodukter i de nuvarande och framtida medlemsstaterna.
(16) I sin resolution av den 8 juni 1998(5) godkände rådet kommissionens strategi och handlingsplan för förnybara energikällor och efterlyste särskilda åtgärder när det gäller biodrivmedel.
(17) Kommissionens grönbok "Mot en europeisk strategi för trygg energiförsörjning" ställer upp målet att man senast år 2020 skall ha ersatt 20 % av konventionella drivmedel med alternativa drivmedel inom vägtransportsektorn.
(18) Om alternativa drivmedel skall lyckas komma in på marknaden, måste de vara lättillgängliga och konkurrenskraftiga.
(19) I sin resolution av den 18 juni 1998(6) krävde Europaparlamentet att marknadsandelen för biodrivmedel skulle öka till 2 % under de kommande fem åren genom ett åtgärdspaket som bland annat omfattar skattebefrielse, finansiellt stöd till förädlingsindustrin och fastställande av en obligatorisk andel biodrivmedel för oljeföretag.
(20) Den optimala metoden för att öka andelen biodrivmedel på de nationella marknaderna och gemenskapsmarknaderna är beroende av tillgången på resurser och råvaror, av den nationella politiken och gemenskapspolitiken för att främja biodrivmedel och av skattebestämmelser, samt av att alla intressenter/parter involveras på ett lämpligt sätt.
(21) Nationell politik för att främja användningen av biodrivmedel får inte hindra den fria rörligheten för drivmedel som uppfyller de harmoniserade miljöspecifikationerna i gemenskapslagstiftningen.
(22) Främjande av produktion och användning av biodrivmedel kan bidra till att beroendet av importerad energi och utsläppen av växthusgaser minskar. Dessutom kan biodrivmedel, i ren form eller i blandad form, i princip användas i befintliga motorfordon och användas i nuvarande bränslesystem för fordon. Blandning av biodrivmedel och fossila drivmedel kan underlätta en potentiell minskning av kostnaderna för distributionssystemet i gemenskapen.
(23) Eftersom målet för den föreslagna åtgärden, nämligen införandet av allmänna principer för att en minimiandel biodrivmedel skall kunna marknadsföras och distribueras, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna på grund av åtgärdens omfattning och det därför bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå detta mål.
(24) Forskning och teknisk utveckling när det gäller biodrivmedlens hållbarhet bör främjas.
(25) Ökad användning av biodrivmedel bör åtföljas av en noggrann analys av de miljömässiga, ekonomiska och sociala konsekvenserna för att man skall kunna avgöra huruvida det är lämpligt att öka andelen biodrivmedel i förhållande till konventionella drivmedel.
(26) Det bör föreskrivas ett förfarande för att snabbt anpassa förteckningen över biodrivmedel, andelen förnybart innehåll och tidsplanen för att införa biodrivmedel på transportmarknaden till den tekniska utvecklingen och till resultaten av en miljökonsekvensbedömning av den första introduktionsfasen.
(27) Åtgärder bör vidtas för att snabbt utveckla kvalitetsstandarderna för biodrivmedel som används inom fordonssektorn, både som rena biodrivmedel och som blandningskomponenter i konventionella drivmedel. Även om den biologiskt nedbrytbara delen av avfall är en potentiellt användbar källa för framställning av biodrivmedel, måste det i kvalitetsstandarderna tas hänsyn till att avfallet eventuellt kan vara kontaminerat, så att inte vissa komponenter skadar fordonet eller förvärrar utsläppen.
(28) Stödet för att främja användningen av biodrivmedel bör ske i överensstämmelse med försörjningstrygghet och miljömål, liksom de politiska målen och åtgärderna på området i varje medlemsstat. När så är fallet kan medlemsstaterna överväga vilka kostnadseffektiva sätt som finns för att informera om möjligheterna att använda biodrivmedel.
(29) De åtgärder som är nödvändiga för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(7).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syftet med detta direktiv är att främja användningen av biodrivmedel eller andra förnybara drivmedel som skall ersätta diesel eller bensin för transportändamål i varje medlemsstat, för att på så sätt bidra till mål som t.ex. att uppfylla åtaganden som rör klimatförändringar, bidra till försörjningstryggheten på ett miljövänligt sätt och främja förnybara energikällor.
Artikel 2
1. I detta direktiv avses med
a) biodrivmedel: flytande eller gasformigt bränsle för transport, som framställs av biomassa,
b) biomassa: den biologiskt nedbrytbara delen av produkter, avfall och restprodukter från jordbruk (inklusive material av vegetabiliskt och animaliskt ursprung), skogsbruk och därmed förknippad industri, liksom den biologiskt nedbrytbara delen av industriavfall och kommunalt avfall,
c) andra förnybara drivmedel: andra förnybara bränslen än biodrivmedel, som framställs från förnybara energikällor enligt definitionen i direktiv 2001/77/EG(8) och som används för transportändamål,
d) energiinnehåll: det nedre värmevärdet för ett drivmedel.
2. Åtminstone de produkter som förtecknas nedan skall anses vara biodrivmedel:
a) bioetanol: etanol som framställs av biomassa och/eller den biologiskt nedbrytbara delen av avfall och som skall användas som biodrivmedel.
b) biodiesel: metylester av dieselkvalitet från vegetabilisk eller animalisk olja, som skall användas som biodrivmedel.
c) biogas: en bränslegas som framställs av biomassa och/eller den biologiskt nedbrytbara delen av avfall som kan renas till naturgaskvalitet och som skall användas som biodrivmedel, eller vedgas.
d) biometanol: metanol som framställs av biomassa och skall användas som biodrivmedel.
e) biodimetyleter: dimetyleter som framställs av biomassa och skall användas som biodrivmedel.
f) bio-ETBE (etyltertiärbutyleter): ETBE som framställs av bioetanol. Volymandelen biodrivmedel i bio-ETBE beräknas till 47 %.
g) bio-MTBE (metyltertiärbutyleter): bränsle som framställs av biometanol. Volymandelen biodrivmedel i bio-MTBE beräknas till 36 %.
h) syntetiska biodrivmedel: syntetiska kolväten eller blandningar av syntetiska kolväten, som framställs av biomassa.
i) bioväte: vätgas som framställs av biomassa och/eller den biologiskt nedbrytbara delen av avfall, och som skall användas som biodrivmedel.
j) ren vegetabilisk olja: olja framställd från oljeväxter genom pressning, extraktion eller jämförbara metoder, rå eller raffinerad men kemiskt oförändrad, då den är förenlig med motortyperna och motsvarande utsläppskrav.
Artikel 3
1. a) Medlemsstaterna bör se till att en minsta andel biodrivmedel och andra förnybara bränslen släpps ut på deras marknader och skall fastställa nationella vägledande mål för detta.
b) i) Ett referensvärde för dessa mål skall vara 2 %, beräknat på energiinnehållet, av all bensin och diesel för transportändamål som släpps ut på deras marknader, senast den 31 december 2005.
ii) Ett referensvärde för dessa mål skall vara 5,75 %, beräknat på energiinnehållet, av all bensin och diesel för transportändamål som släpps ut på deras marknader, senast den 31 december 2010.
2. Biodrivmedel får tillhandahållas i följande form:
a) Rena biodrivmedel eller mineraloljederivat med hög halt av biodrivmedel i enlighet med särskilda kvalitetsnormer för transporttillämpningar.
b) Biodrivmedel som blandats i mineraloljederivat i enlighet med de tillämpliga europeiska standarder som beskriver de tekniska specifikationerna för drivmedel (EN 228 och EN 590).
c) Vätskor som framställs av biodrivmedel, t.ex. ETBE (etyltertiärbutyleter), som innehåller den procentandel biodrivmedel som anges i artikel 2.2.
3. Medlemsstaterna skall övervaka effekterna av en användning i icke-anpassade fordon av dieselblandningar som består av mer än 5 % biodrivmedel och skall, om så krävs, vidta åtgärder för att se till att den tillämpliga gemenskapslagstiftningen om utsläppsnormer följs.
4. Medlemsstaterna bör i sina åtgärder ta hänsyn till vilken inverkan på den totala klimat- och miljöbalansen som de olika biodrivmedlen och andra förnybara drivmedel har och får prioritera främjandet av sådana drivmedel som ger en mycket god kostnadseffektiv miljöbalans med beaktande av konkurrenskraft och försörjningstrygghet.
5. Medlemsstaterna skall se till att allmänheten upplyses om att biodrivmedel och andra förnybara drivmedel finns tillgängliga. Det skall föreskrivas att biodrivmedel som blandats i mineraloljederivat och som överstiger gränsvärdet på 5 % för fettsyrametylestrar (FAME) eller 5 % för bioetanol skall förses med en särskild märkning vid försäljningsställena.
Artikel 4
1. Medlemsstaterna skall före den 1 juli varje år rapportera till kommissionen om
- vilka åtgärder som vidtagits för att främja användningen av biodrivmedel eller andra förnybara drivmedel som skall ersätta diesel eller bensin för transportändamål,
- de nationella resurser som anslagits för produktion av biomassa för annan energianvändning än transport, och
- det föregående årets totala försäljning av drivmedel samt andelen biodrivmedel, rena eller blandade, och andra förnybara drivmedel som släppts ut på marknaden. I förekommande fall skall medlemsstaterna rapportera om exceptionella förhållanden när det gäller utbudet av råolja eller oljeprodukter som har påverkat försäljningen av biodrivmedel och andra förnybara drivmedel.
I sin första rapport efter ikraftträdandet av detta direktiv skall medlemsstaterna ange nivån på sina nationella vägledande mål för den första fasen. I rapporten för år 2006 skall medlemsstaterna ange sina nationella vägledande mål för den andra fasen.
I rapporterna skall avvikelser från de nationella målen i förhållande till referensvärdena i artikel 3.1 b motiveras och kan grundas på följande faktorer:
a) Objektiva faktorer, t.ex. den begränsade nationella potentialen för produktion av biodrivmedel från biomassa.
b) Storleken på de resurser som anslås till produktion av biomassa för annan energianvändning än transport samt de särskilda tekniska eller klimatmässiga förhållanden som kännetecknar den nationella marknaden för drivmedel.
c) Nationella strategier för att anslå jämförbara resurser till produktionen av andra drivmedel som baseras på förnybara energikällor och är förenliga med målen för detta direktiv.
2. Kommissionen skall senast den 31 december 2006 och vartannat år därefter utarbeta och till Europaparlamentet och rådet lämna en utvärderingsrapport om framstegen när det gäller användning av biodrivmedel och andra förnybara drivmedel i medlemsstaterna.
Denna rapport skall åtminstone omfatta följande:
a) Kostnadseffektiviteten för de åtgärder som medlemsstaterna har vidtagit för att främja användningen av biodrivmedel och andra förnybara drivmedel.
b) De ekonomiska aspekterna och miljökonsekvenserna av en ytterligare ökning av andelen biodrivmedel och andra förnybara drivmedel.
c) Biodrivmedel och andra förnybara drivmedel i ett livscykelperspektiv, för att ange möjliga åtgärder för det framtida främjandet av de av dem som är klimat- och miljövänliga och som kan bli konkurrenskraftiga och kostnadseffektiva.
d) Hållbarheten vid odling av grödor som används för att framställa biodrivmedel, särskilt markanvändning, grad av odlingsintensitet, växelbruk och användning av bekämpningsmedel.
e) Bedömning av användningen av biodrivmedel och andra förnybara drivmedel med avseende på deras olika konsekvenser för klimatförändringen och deras påverkan när det gäller att minska koldioxidutsläppen.
f) En genomgång av ytterligare mer långsiktiga alternativ när det gäller åtgärder för energieffektivitet på transportområdet.
Utifrån denna rapport skall kommissionen när det är lämpligt för Europaparlamentet och rådet lägga fram förslag om en anpassning av de mål som anges i artikel 3.1. Om rapportens slutsats blir att de vägledande målen sannolikt inte kommer att uppnås av skäl som är oberättigade och/eller inte hänför sig till nya vetenskapliga rön, skall dessa förslag ta upp nationella mål, inklusive eventuella bindande mål, i en lämplig form.
Artikel 5
Förteckningen i artikel 2.2 får anpassas till den tekniska utvecklingen i enlighet med förfarandet i artikel 6.2. Vid anpassning av förteckningen skall biodrivmedlens inverkan på miljön beaktas.
Artikel 6
1. Kommissionen skall biträdas av en kommitté.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 7
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 december 2004. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texten till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 8
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska unionens officiella tidning.
Artikel 9
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens direktiv 2003/60/EG
av den 18 juni 2003
om ändring av bilagorna till rådets direktiv 76/895/EEG, 86/362/EEG, 86/363/EEG och 90/642/EEG beträffande fastställande av gränsvärden för vissa bekämpningsmedelsrester i och på spannmål, livsmedel av animaliskt ursprung och vissa produkter av vegetabiliskt ursprung, inklusive frukt och grönsaker
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 76/895/EEG av den 23 november 1976 om fastställande av gränsvärden för bekämpningsmedelsrester i och på frukt och grönsaker(1), senast ändrat genom kommissionens direktiv 2002/79/EG(2), särskilt artikel 5 i detta,
med beaktande av rådets direktiv 86/362/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på spannmål(3), senast ändrat genom direktiv 2002/79/EG, särskilt artikel 10 i detta,
med beaktande av rådets direktiv 86/363/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på livsmedel av animaliskt ursprung(4), senast ändrat genom direktiv 2002/79/EG(5), särskilt artikel 10 i detta,
med beaktande av rådets direktiv 90/642/EEG av den 27 november 1990 om fastställande av gränsvärden för bekämpningsmedelsrester i och på produkter av vegetabiliskt ursprung inklusive frukt och grönsaker(6), senast ändrat genom kommissionens direktiv 2002/100/EG, särskilt artikel 7 i detta,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(7), senast ändrat genom kommissionens direktiv 2003/39/EG(8), särskilt artikel 4.1 f i detta, och
av följande skäl:
(1) De befintliga verksamma ämnena amitrol, dikvat, isoproturon och etofumesat infördes i bilaga I till rådets direktiv 91/414/EEG genom kommissionens direktiv 2001/21/EG(9), 2002/18/EG(10) respektive 2002/37/EG(11).
(2) De nya verksamma ämnena fenhexamid, acibenzolar-S-metyl, cyklanilid, pyraflufenetyl, iprovalikarb, prosulfuron, sulfosulfuron, cinidonetyl, cyhalofopbutyl, famoxadon, florasulam, metalaxyl-M, pikolinafen och flumioxazin infördes i bilaga I till direktiv 91/414/EEG genom kommissionens direktiv 2001/28/EG(12), 2001/87/EG(13), 2002/48/EG(14), 2002/64/EG(15) och 2002/81/EG(16).
(3) Införandet av de berörda verksamma ämnena i bilaga I till direktiv 91/414/EEG grundades på en utvärdering av de uppgifter som lämnats in om det föreslagna användningsområdet. Uppgifterna om användningen har lämnats in av vissa medlemsstater i enlighet med artikel 4.1 f i direktiv 91/414/EEG. Tillgängliga uppgifter har nu gåtts igenom, och de har befunnits vara tillräckliga för att vissa gränsvärden för bekämpningsmedelsrester skall kunna fastställas.
(4) Om det inte finns något permanent eller provisoriskt gränsvärde för bekämpningsmedelsrester på gemenskapsnivå måste medlemsstaterna fastställa ett provisoriskt nationellt gränsvärde i enlighet med artikel 4.1 f i direktiv 91/414/EEG innan växtskyddsmedel som innehåller dessa verksamma ämnen kan godkännas.
(5) För de verksamma ämnena klorfenapyr, fentinacetat och fentinhydroxid fattades beslut om att inte införa dem i bilaga I till direktiv 91/414/EEG genom kommissionens direktiv 2001/697/EG(17), 2002/478/EG(18) respektive 2002/479/EG(19). I besluten föreskrivs att användningen av växtskyddsmedel som innehåller dessa verksamma ämnen inte längre skall vara tillåten i gemenskapen. Det är därför nödvändigt att alla bekämpningsmedelsrester som uppstår genom användning av dessa växtskyddsmedel läggs till i bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG för att möjliggöra en ordentlig övervakning och kontroll av förbuden mot användning och för att skydda konsumenterna.
(6) För att berättigade förväntningar beträffande användning av befintliga lager av bekämpningsmedel skall kunna uppfyllas ges i kommissionens beslut om att inte godkänna de verksamma ämnena möjlighet till en utfasningsperiod, och därför bör beslut om gränsvärden för bekämpningsmedelsrester där ingen användning av det berörda ämnet är tillåten inom gemenskapen inte börja gälla förrän efter utgången av utfasningsperioden för det ämnet.
(7) Gemenskapens gränsvärden och de värden som rekommenderas i Codex alimentarius fastställs och utvärderas genom liknande förfaranden. I Codex alimentarius anges ett begränsat antal gränsvärden för dikvat och fentin (-acetat eller -hydroxid). Dessa har beaktats vid fastställandet av de gränsvärden som anges i detta direktiv. De gränsvärden i Codex alimentarius som inom en nära framtid kommer att rekommenderas att dras tillbaka har inte beaktats. De gränsvärden som grundas på gränsvärden i Codex alimentarius har utvärderats med avseende på riskerna för konsumenterna, och inga risker kunde påvisas med de toxikologiska endpoints som var baserade på studier som var tillgängliga för kommissionen.
(8) I samband med att de berörda verksamma ämnena infördes i eller uteslöts från bilaga I till direktiv 91/414/EEG avslutades de tekniska och vetenskapliga utvärderingarna genom kommissionens granskningsrapport. Utvärderingsrapporterna för de nämnda ämnena avslutades de datum som anges i de kommissions direktiv som anförs i skäl 1 och 2 samt i de kommissionsbeslut som anförs i skäl 5. I dessa rapporter fastställdes acceptabelt dagligt intag (ADI) och om nödvändigt akut referensdos (ARfD) för de berörda ämnena. Konsumenternas livstidsexponering genom livsmedel som behandlats med det berörda verksamma ämnet har uppskattats och utvärderats med hjälp av de metoder som används inom gemenskapen. Hänsyn har också tagits till de riktlinjer som offentliggjorts av Världshälsoorganisationen(20) samt yttrandet om de använda metoderna från den Vetenskapliga kommittén för växter(21). Slutsatsen har dragits att de föreslagna gränsvärdena inte leder till att acceptabla dagliga intag eller akuta referensdoser överskrids.
(9) För att konsumenterna skall få tillräckligt skydd mot exponering för bekämpningsmedelsrester till följd av otillåten användning av växtskyddsprodukter, bör de provisoriska gränsvärden som fastställs för de berörda kombinationerna av produkter/bekämpningsmedel motsvara den lägsta analytiska bestämningsgränsen.
(10) Att provisoriska gränsvärden fastställs på gemenskapsnivå hindrar inte medlemsstaterna från att fastställa provisoriska gränsvärden för de ämnen som anges i det här direktivet i enlighet med artikel 4.1 f i direktiv 91/414/EEG och bilaga VI till det direktivet. Fyra år anses vara en tillräckligt lång period för att godkänna ytterligare användningsområden för de berörda verksamma ämnena. De provisoriska gränsvärdena bör därefter bli permanenta.
(11) Det är därför nödvändigt att förteckna samtliga de bekämpningsmedelsrester som härrör från användningen av dessa växtskyddsprodukter i bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG för att möjliggöra en ändamålsenlig övervakning och kontroll av användningsförbudet och för att skydda konsumenterna. Bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG bör därför ändras.
(12) För att möjliggöra att det fastställs gränsvärden för resthalter av dikvat måste bestämmelserna i direktiv 76/895/EEG överföras till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG, och dessa bestämmelser måste strykas i direktiv 76/895/EEG. En del av dessa bestämmelser bör ändras som ett resultat av vetenskapliga och tekniska framsteg och på grund av förändrad användning och ändrade godkännanden på nationell nivå och gemenskapsnivå.
(13) Detta direktiv är förenligt med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilaga II till direktiv 76/895/EEG skall posterna beträffande dikvat utgå.
Artikel 2
De gränsvärden för bekämpningsmedelsrester som anges i bilaga I till detta direktiv skall läggas till i del A i bilaga II till direktiv 86/362/EEG.
Artikel 3
De gränsvärden för bekämpningsmedelsrester som anges i bilagorna II och III till detta direktiv skall läggas till i del A och B i bilaga II till direktiv 86/363/EEG.
Artikel 4
De gränsvärden för bekämpningsmedelsrester som anges i bilaga IV till detta direktiv skall läggas till i bilaga II till direktiv 90/642/EEG.
Artikel 5
Medlemsstaterna skall senast den 30 juni 2003 sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv, med undantag för bestämmelserna för fentinhydroxid, fentinacetat och klorfenapyr, som skall sättas i kraft senast den 30 juni 2004. De skall genast underrätta kommissionen om detta.
De skall tillämpa dessa bestämmelser från och med den 1 juli 2003, med undantag för bestämmelserna för fentinhydroxid, fentinacetat och klorfenapyr, som skall tillämpas från och med 1 juli 2004.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 6
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska unionens officiella tidning.
Artikel 7
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 568/2003
av den 28 mars 2003
om rättelse av de engelska och nederländska versionerna av förordning (EG) nr 2603/1999 om regler för övergången till den ordning för stöd till landsbygdens utveckling som föreskrivs i rådets förordning (EG) nr 1257/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1257/1999 av den 17 maj 1999 om stöd från Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) till utveckling av landsbygden och om ändring och upphävande av vissa förordningar(1), särskilt artikel 53.1 i denna, och
av följande skäl:
(1) Det är fel i de engelska och nederländska versionerna av kommissionens förordning (EG) nr 2603/1999(2), senast ändrad genom förordning (EG) nr 2055/2001(3). Dessa språkversioner bör därför rättas.
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för jordbrukets struktur och landsbygdens utveckling.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Rättelsen rör bara den nederländska versionen.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
Kommissionens förordning (EG) nr 1053/2003
av den 19 juni 2003
om ändring av Europaparlamentets och rådets förordning (EG) nr 999/2001 när det gäller snabbtest
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 999/2001 av den 22 maj 2001 om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati(1), senast ändrad genom kommissionens förordning (EG) nr 260/2003(2), särskilt första stycket i artikel 23 i denna, och
av följande skäl:
(1) I förordning (EG) nr 999/2001 fastställs för tillämpningen av den förordningen en förteckning över nationella referenslaboratorier för TSE. Grekland har bytt nationellt referenslaboratorium.
(2) I förordning (EG) nr 999/2001 fastställs även en förteckning över snabbtest som har godkänts för övervakning av TSE.
(3) Det företag som marknadsför ett av de snabbtest som har godkänts för TSE-övervakning har meddelat kommissionen att det har för avsikt att marknadsföra testet under ett nytt handelsnamn.
(4) Vetenskapliga styrkommittén rekommenderade i sitt yttrande av den 6 och 7 mars 2003 att två nya test skulle införas i förteckningen över de snabbtest som godkänts för övervakning av bovin spongiform encefalopati (BSE). Tillverkarna av båda testen har presenterat data som visar att deras test också får användas för övervakning av TSE hos får.
(5) För att garantera att godkända snabbtest håller samma prestandanivå efter godkännandet bör ett förfarande fastställas för eventuella ändringar av testet eller testprotokollet.
(6) Förordning (EG) nr 999/2001 bör därför ändras.
(7) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga X till förordning (EG) nr 999/2001 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Kommissionens förordning (EG) nr 1139/2003
av den 27 juni 2003
om ändring av Europaparlamentets och rådets förordning (EG) nr 999/2001 när det gäller övervakningsprogram och specificerat riskmaterial
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 999/2001 av den 22 maj 2001 om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati(1), senast ändrad genom kommissionens förordning (EG) nr 1053/2003(2), särskilt artikel 23 i denna, och
av följande skäl:
(1) Förordning (EG) nr 999/2001 innehåller bestämmelser om övervakning av transmissibel spongiform encefalopati (TSE) hos får och getter, inklusive övervakning av ett urval av djur som inte slaktas för att användas som livsmedel. Det är nödvändigt att klargöra definitionen av denna grupp av djur för att undvika olämplig riktning av proven.
(2) I förordning (EG) nr 999/2001 föreskrivs utrotningsåtgärder efter det att TSE har bekräftats hos får och getter. För att samla in epidemiologisk information bör riktade prov tas av djur som destruerats genom åtgärderna.
(3) Det finns en teoretisk möjlighet att bovin spongiform encefalopati (BSE) förekommer i får- och getpopulationen. Det är omöjligt att genom rutinmetoder skilja mellan BSE- och skrapiesmitta hos dessa djur. Infektiviteten i nedre delen av tunntarmen (ileum) är vid båda sjukdomarna signifikant redan i ett tidigt skede av infektionen. Som en förebyggande åtgärd bör ileum från får och getter i alla åldrar tillföras förteckningen över specificerat riskmaterial.
(4) I Vetenskapliga styrkommitténs yttrande av den 7 och 8 november 2002 om TSE-infektivitetens distribution i vävnader från idisslare rekommenderas att tonsiller från nötkreatur i alla åldrar bör anses medföra risk för BSE.
(5) Vetenskapliga styrkommittén har fastställt att kontaminering med vävnader från det centrala nervsystemet och tonsiller måste undvikas när tunga och kött från huvud tas ut från nötkreatur för att användas som livsmedel, för att undvika alla BSE-risker.
(6) Eftersom huvudets tillstånd huvudsakligen är beroende av att det hanteras varsamt och att skotthålet i pannan förseglas på ett säkert sätt liksom foramen magnum, måste det finnas kontrollsystem i slakterierna och i de styckningsanläggningar som särskilt godkänts.
(7) Bestämmelserna om sändning av slaktkroppar, halva slaktkroppar och kvartsparter av slaktkroppar som inte innehåller annat specificerat riskmaterial än ryggraden till övriga medlemsstater utan deras förhandsgodkännande bör utvidgas till att omfatta halva slaktkroppar som styckats i högst tre grossistdelar för att återspegla den faktiska handeln mellan medlemsstater.
(8) Europaparlamentets og rådets förordning (EG) nr 1774/2002(3), ändrad genom kommissionens förordning (EG) nr 808/2003(4), innehåller bestämmelser om djur- och folkhälsa vid insamling, transport, lagring, hantering, bearbetning och användning eller bortskaffande av alla animala biprodukter som inte skall användas som livsmedel, inklusive deras avyttring och, i vissa undantagsfall, export och transitering. Särskilda bestämmelser om avlägsnande och bortskaffande av sådana produkter i bilaga XI till förordning (EG) nr 999/2001 bör därför utgå.
(9) Förordning (EG) nr 999/2001 bör därför ändras.
(10) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagorna III och XI till förordning (EG) nr 999/2001 skall ändras i enlighet med bilagan till denna förordning.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Europaparlamentets och rådets förordning (EG) nr 1267/2003
av den 16 juni 2003
om ändring av rådets förordning (EG) nr 2223/96 med avseende på tidsfrister för sändningen av huvudaggregaten i nationalräkenskaperna, undantag när det gäller sändningen av huvudaggregaten i nationalräkenskaperna och sändning av uppgifter om sysselsättning angivna i arbetade timmar
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 285 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europeiska centralbankens yttrande(2),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Rådets förordning (EG) nr 2223/96 av den 25 juni 1996 om det europeiska national- och regionalräkenskapssystemet(4), innehåller en referensram bestående av gemensamma standarder, definitioner, klassifikationer och bokföringsregler för sammanställande av medlemsstaternas räkenskaper för gemenskapens statistikbehov, för att sinsemellan jämförbara resultat skall erhållas från medlemsstaterna.
(2) I den rapport om statistiska krav i den ekonomiska och monetära unionen (EMU), som framlagts av Monetära kommittén, och som godkändes av Ekofinrådet den 18 januari 1999, framhålls att effektiv övervakning och samordning av den ekonomiska politiken är av största vikt för den inre marknaden, och att detta kräver ett omfattande statistiksystem genom vilket beslutsfattarna förses med ett nödvändigt beslutsunderlag. I rapporten talas också om vikten av att sådana uppgifter finns tillgängliga för gemenskapen, i synnerhet för de medlemsstater som deltar i euroområdet.
(3) I rapporten betonades att man inom EMU kommer att behöva ägna större uppmärksamhet åt jämförelser mellan de olika ländernas arbetsmarknader.
(4) För att den kvartalsvisa statistiken skall kunna sammanställas för euroområdet, bör den beviljade tidsfristen för sändningen av huvudaggregaten i nationalräkenskaperna minskas till 70 dagar.
(5) Kvartalsvisa och årliga undantag som beviljats medlemsstaterna och som hindrar sammanställandet av huvudaggregaten i nationalräkenskaperna för euroområdet och gemenskapen bör avskaffas.
(6) I handlingsplanen avseende den statistik som krävs i samband med den ekonomiska och monetära unionen, godkänd av Ekofin-rådet den 29 september 2000, fastställs att leverans av sysselsättningsuppgifter i nationalräkenskaperna i enheten "arbetade timmar" prioriteras.
(7) Kommittén för det statistiska programmet och kommittén för valuta-, finans- och betalningsbalansstatistik har rådfrågats i enlighet med artikel 3 i rådets beslut 89/382/EEG, Euratom(5) och rådets beslut 91/115/EEG(6).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga B till förordning (EG) nr 2223/96 ändras enligt följande:
1. Texten som följer på rubriken "Leveransprogram för nationalräkenskapsdata" skall ändras på följande sätt:
a) Texten till "Tabellöversikt" skall ersättas med texten i bilaga I.
b) Texten till tabell 1, "Huvudaggregat - kvartalsvis och årlig redovisning" skall ersättas med texten i bilaga II.
2. Texten som följer på rubriken: "Avvikelser beträffande de tabeller som skall sändas i enlighet med frågeformuläret "ESA-95" per land" skall ersättas med texten i bilaga III.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Kommissionens förordning (EG) nr 1914/2003
av den 30 oktober 2003
om ändring av förordning (EG) nr 1488/2001 om tillämpningsföreskrifter för rådets förordning (EG) nr 3448/93 när det gäller att hänföra vissa kvantiteter av vissa basprodukter enligt bilaga I till Fördraget om upprättandet av Europeiska gemenskapen till förfarandet för aktiv förädling utan förhandskontroll av de ekonomiska kraven
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EG) nr 3448/93 av den 6 december 1993 om systemet för handeln med vissa varor som framställs genom bearbetning av jordbruksprodukter(1), senast ändrad genom förordning (EG) nr 2580/2000(2), särskilt artikel 11.1 tredje stycket i denna, och
av följande skäl:
(1) I artikel 11.1 i förordning (EG) nr 3448/93 föreskrivs att de ekonomiska villkor som anges i artikel 117 c i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3), senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 2700/2000(4), skall betraktas som uppfyllda för att tillåta att vissa kvantiteter av vissa basprodukter får hänföras till förfarandet för aktiv förädling för att användas vid framställning av varor. De detaljerade tillämpningsföreskrifter till denna bestämmelse som gör det möjligt att fastställa vilka basjordbruksprodukter som får hänföras till förfarandet för aktiv förädling samt att kontrollera och planera kvantiteterna därav, skall antas i enlighet med artikel 16 i förordning (EG) nr 3448/93.
(2) Kommissionens förordning (EG) nr 1488/2001(5), bör ändras för att klargöra att de förfaranden som avses i artikel 16 i förordning (EG) nr 3448/93 är tillämpliga för att fastställa vilka basjordbruksprodukter som skall hänföras till förfarandet för aktiv förädling samt för att kontrollera och planera kvantiteterna av dessa produkter.
(3) De åtgärder som föreskrivs i denna förordning står i överensstämmelse med yttrandet från Kommittén för övergripande frågor rörande handel med bearbetade jordbruksprodukter som inte omfattas av bilaga I till fördraget.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 1488/2001 ändras enligt följande:
1. I artikel 2 skall punkt 2 ersättas av följande:
"2. Om behoven av bidrag beräknas bli större än de tillgängliga ekonomiska medlen, skall kvantiteterna av de olika produkter som anges med sin åttasiffriga KN-kod, fastställas i enlighet med artikel 11.1 i förordning (EG) nr 3448/93 och med hjälp av prognosen."
2. I artikel 22 skall det andra stycket ersättas med följande:"Om de bidrag som skall betalas ut beräknas bli större än de tillgängliga ekonomiska medlen, skall den återstående kvantiteten för varje basprodukt fastställas i enlighet med artikel 11.1 i förordning (EG) nr 3448/93 med beaktande av redan licensierade kvantiteter och av de icke-utnyttjade kvantiteter som kommissionen informerats om i enlighet med artikel 25 i denna förordning. Denna kvantitet skall offentliggöras i Europeiska unionens officiella tidning en andra gång senast den 31 januari varje år och en tredje gång senast den 31 maj varje år."
3. Artikel 24 skall ersättas av följande:
"Artikel 24
Utfärdande av AF-licenser i nödfall
Kommissionens förordning (EG) nr 2151/2003
av den 16 december 2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 2195/2002 av den 5 november 2002 om en gemensam terminologi vid offentlig upphandling (CPV)(1), särskilt artikel 2 i denna, och
av följande skäl:
(1) Genom förordning (EG) nr 2195/2002 fastställdes ett enda klassificeringssystem för offentlig upphandling i syfte att standardisera de referenser som används av upphandlande myndigheter och enheter för att beskriva föremålet för upphandlingen.
(2) Uppbyggnaden av och koderna i CPV kan behöva anpassas, eller till och med ändras, i enlighet med marknadens utveckling och användarnas behov.
(3) Uppbyggnaden av och koderna i CPV bör uppdateras för att ta hänsyn till de särskilda behov som medlemsstaterna och användarna av CPV gett uttryck för samt för att rätta sakfel i de olika språkversionerna.
(4) De tekniska ändringar och förbättringar som kartlagts under lagstiftningsprocessen inför antagandet av förordning (EG) nr 2195/2002 men som inte kunde tas med i den förordningen, bör införas i samma förordnings bilagor.
(5) I sitt yttrande(2) om förslaget till en förordning om CPV poängterade Regionkommittén att klassificeringen av läkemedel måste förbättras och rekommenderade att Världshälsoorganisationens klassificeringssystem, ATC (Anatomic Therapeutic Chemical), används för att komplettera CPV-systemet och dess koder för läkemedel.
(6) Berörda parter och CPV-användare har bidragit med förslag till förbättring av CPV.
(7) Uppdateringen av CPV-koderna och CPV-strukturen bör även återspeglas i de vägledande konverteringstabellerna mellan CPV och FN:s centrala produktindelning (CPC Prov.), Europeiska gemenskapens statistiska näringsgrensindelning (NACE Rev. 1) och Kombinerade nomenklaturen (KN).
(8) För tydlighetens skull bör CPV och konverteringstabellen mellan CPV och CPC Prov. ersättas i sin helhet. Alla ändringar i CPV-koderna eller i deras beskrivningar bör anges i en separat ny bilaga till förordning (EG) nr 2195/2002.
(9) I och med att kommissionens förordning (EG) nr 204/2002 av den 19 december 2001 om ändring av rådets förordning (EEG) nr 3696/93 om den statistiska indelningen av produkter efter näringsgren (CPA) inom Europeiska ekonomiska gemenskapen(3) trädde i kraft, har konverteringstabellen mellan CPV och CPA 96 i bilaga II till förordning (EG) nr 2195/2002 blivit inaktuell.
(10) I gemensam ståndpunkt (EG) nr 33/2003 antagen av rådet den 20 mars 2003 inför antagandet av Europaparlamentets och rådets direktiv om samordning av förfarandena vid offentlig upphandling av byggentreprenader, varor och tjänster(4) och gemensam ståndpunkt (EG) nr 34/2003, antagen av rådet den 20 mars 2003 inför antagandet av Europaparlamentets och rådets direktiv om samordning av förfarandena vid upphandling på områdena vatten, energi, transporter och posttjänster(5), fastställs inte varuområden efter den statistiska indelningen av produkter efter näringsgren (CPA).
(11) Konverteringstabellen mellan CPV och CPA 96 i bilaga II till förordning (EG) nr 2195/2002 behöver därför inte uppdateras. Bilagan bör därför utgå.
(12) Förordning (EG) nr 2195/2002 bör därför ändras.
(13) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Rådgivande kommittén för offentlig upphandling.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 2195/2002 skall ändras enligt följande:
Bilaga I skall ersättas med texten i bilaga I till denna förordning.
Bilaga II skall ersättas med texten i bilaga II till denna förordning.
Bilaga III skall ersättas med texten i bilaga III till denna förordning.
Bilaga IV skall ändras i enlighet med bilaga IV till denna förordning.
Bilaga V skall ändras i enlighet med bilaga V till denna förordning.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Kommissionens förordning (EG) nr 317/2004
av den 23 februari 2004
om antagande av undantag för Österrike, Frankrike och Luxemburg från bestämmelserna i Europaparlamentets och rådets förordning (EG) nr 2150/2002 om avfallsstatistik
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 2150/2002 av den 25 november 2002 om avfallsstatistik(1), särskilt artikel 4.1 i denna,
med beaktande av Österrikes begäran av den 30 juni 2003,
med beaktande av Frankrikes begäran av den 12 juni 2003,
med beaktande av Luxemburgs begäran av den 25 juni 2003, och
av följande skäl,
(1) I enlighet med artikel 4.1 i förordning (EG) nr 2150/2002 får kommissionen under en övergångsperiod bevilja undantag från vissa bestämmelser i bilagorna till förordningen.
(2) Efter begäran bör sådana undantag beviljas Österrike, Frankrike och Luxemburg.
(3) Åtgärderna som fastställs i den här förordningen överensstämmer med yttrandet från Kommittén för det statistiska programmet som inrättades genom rådets beslut 89/382/EEG, Euratom(2).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Följande undantag från bestämmelserna i förordning (EG) nr 2150/2002 beviljas härmed:
a) Österrike beviljas undantag för redovisning av resultat avseende avsnitt 8.1.1, post 1 (jordbruk, jakt och skogsbruk) i bilaga I.
b) Frankrike beviljas undantag för redovisning av resultat avseende avsnitt 8.1.1, posterna 1 (jordbruk, jakt och skogsbruk), 2 (fiske) och 16 (tjänster) i bilaga I samt de som avser avsnitt 8.2 i bilaga II.
c) Luxemburg beviljas undantag för redovisning av resultat avseende avsnitt 8.1.1, posterna 1 (jordbruk, jakt och skogsbruk) och 2 (fiske) i bilaga I.
2. De undantag som beviljas i punkt 1 gäller endast uppgifter från det första referensåret, dvs. 2004.
Efter övergångsperiodens utgång skall Österrike, Frankrike och Luxemburg redovisa uppgifter från referensåret 2006.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den offentliggjorts i Europeiska unionens officiella tidning.
