med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 75.1 i detta,
Den gemensamma marknadens successiva uppbyggnad får inte försvåras av hinder inom transportsektorn. Det är nödvändigt att säkerställa en gradvis utbyggnad av de internationella godstransporterna på väg med tanke på utvecklingen av handeln och varuflödena inom gemenskapen.
1. Senast vid utgången av år 1962 skall varje medlemsstat, på det sätt som fastställts i punkterna 2 och 3 av denna artikel, liberalisera de typer av internationella yrkesmässiga vägtransporter som berör andra medlemsstater och som är förtecknade i bilagorna 1 och 2 till detta direktiv, om sådan transport utförs till eller från medlemsstaten eller passerar dess territorium i transit.
4. De båda bilagorna till detta direktiv skall utgöra en del av själva direktivet.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Exportlicenser för ris och brutet ris gäller till och med den femte månaden efter utfärdandemånaden men det finns för sådana produkter sällan en verkligt representativ terminsmarknad, annat än för den eller de närmaste terminerna. Det bör därför vara möjligt att fastställa ett korrektionsbelopp som är lägre än den ovannämnda skillnaden.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"När det exportbidrag för ris och brutet ris som anges i artikel 17.4 första stycket i förordning nr 359/67/EEG förutfastställs, skall exportbidraget vara det som gäller för export den dag då ansökan om exportlicens inlämnas - med avdrag för ett belopp som inte överstiger skillnaden mellan cif-priset för terminsköp och cif-priset, när det förstnämnda överstiger det sistnämnda med mer än 0,025 räkneenheter per 100 kg,
Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(1),
Förordningen av den 31 mars 1969 om "Sammansättningen hos avgaser som släpps ut från bensinmotorer i motorfordon" publicerades i Frankrike den 17 maj 1969 i Journal officiel. Förordningen gäller - från och med den 1 september 1971 för typgodkända fordon med en ny motortyp, dvs. en motortyp som inte tidigare monterats i ett typgodkänt fordon,
Vidare måste de tekniska kraven snabbt anpassas med hänsyn till tekniska framsteg. Därför bör det förfarande kunna tillämpas som fastslås i artikel 13 i rådets direktiv av den 6 februari 1970 om typgodkännande av motorfordon och släpvagnar till dessa fordon.
I detta direktiv avses med fordon varje fordon med förbränningsmotor med styrd tändning, avsett att användas på väg, med eller utan karosseri, som har minst fyra hjul, med en tillåten totalvikt på minst 400 kg och som är konstruerat för en högsta hastighet som uppgår till minst 50 km/tim. Jordbrukstraktorer, lantbruksmaskiner och arbetsfordon är undantagna.
- från och med den 1 oktober 1971, om fordonet även uppfyller kraven i punkt 3.2.1.1 och 3.2.2.1 i bilaga 1 och kraven i bilaga 3.
2. Bestämmelserna i 1 skall upphävas så snart rådets direktiv av den 6 februari 1970 om typgodkännande av motorfordon och släpvagnar till dessa fordon träder i kraft.
Artikel 5
1. Medlemsstaterna skall anta bestämmelser som innehåller de krav som är nödvändiga för att följa detta direktiv före den 30 juni 1970 och skall genast underrätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 103 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande, och
Förfaranden och instrument, lämpade att säkerställa ett snabbt genomförande av de åtgärder som är avsedda att dämpa försörjningssvårigheterna i fråga om råolja eller petroleumprodukter, bör fastställas i förväg.
I övrigt är det lämpligt att omedelbart bilda ett samrådsorgan som kan underlätta samordningen av konkreta åtgärder som medlemsstaterna kan ha vidtagit eller planerat på detta område.
Artikel 1
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättande av ett gemensamt råd och en gemensam kommission,
med beaktande av följande: Med hänsyn till en dom som nyligen avkunnats av domstolen samt till vissa tvingande sociala krav verkar det önskvärt att ändra en bestämmelse i rådets förordning (EEG, Euratom, EKSG) nr 260/681 av den 29 februari 1968 om villkoren för och förfarandet vid skatt till Europeiska gemenskaperna, senast ändrad genom förordning (Euratom, EKSG, EEG) nr 2531/722.
Rådets förordning (EEG, Euratom, EKSG) nr 260/68 av den 29 februari 1968 ändras på följande sätt:
RÅDETS DIREKTIV av den 17 december 1973 om tillnärmning av medlemsstaternas lagstiftning om inredningsdetaljer i motorfordon (passagerarutrymmets inre delar frånsett inre backspeglar, manöverorganens utformning, taket eller det öppningsbara taket, ryggstödet och sätenas baksida) (74/60/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: De tekniska krav som motorfordon måste uppfylla enligt nationell lagstiftning gäller bl.a. inredning avsedd att skydda föraren och passagerarna.
Harmoniserade krav bör minska risken för eller graden av skador i samband med olyckor som motorfordonsförare kan bli offer för och trygga trafiksäkerheten inom hela gemenskapen.
Artikel 1
Ingen medlemsstat får vägra att bevilja EEG-typgodkännande eller nationellt typgodkännande för ett fordon av skäl som hänför sig till sådana inredningsdetaljer som
- ryggstödet eller sätenas baksida,
Ingen medlemsstat får vägra eller förbjuda att ett fordon saluförs, registreras, tas i bruk eller används, av skäl som hänför sig till - passagerarutrymmets inre delar frånsett inre backspeglar,
- ryggstödet eller sätenas baksida,
Den medlemsstat som har beviljat EEG-typgodkännande måste vidta de åtgärder som krävs för att hålla sig informerad om varje ändring av en sådan del eller egenskap som avses i bilaga 1 punkt 2.2. De behöriga myndigheterna i staten skall avgöra om nya provningar behöver utföras på den ändrade fordonstypen och en ny rapport utformas. Om dessa provningar visar att kraven i detta direktiv inte uppfylls skall ändringen inte godkännas.
Artikel 6
Artikel 7
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag, och
Artikel 1
Denna förordning skall tillämpas från och med den 1 april 1974.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(1),
Dessa hinder för upprättandet av en väl fungerande gemensam marknad kan avlägsnas, om alla medlemsstater antar samma specifikationer, antingen utöver eller i stället för dem som fastlagts i deras nuvarande lagstiftning, och dessa specifikationer speciellt avser tillverkning och fyllning av aerosolbehållare och den volym de får anges ha.
Det är möjligt att vissa aerosolbehållare som finns på marknaden kan innebära en säkerhetsrisk, trots att de uppfyller kraven i detta direktiv och dess bilaga. Ett förfarande måste därför fastläggas för att motverka denna risk.
Detta direktiv skall gälla aerosolbehållare enligt definitionen i artikel 2 med undantag av sådana som har mindre volym än maximalt 50 ml och sådana som har större volym än vad som anges i punkt 3.1, 4.1.1, 4.2.1, 5.1 och 5.2 i bilagan till detta direktiv.
Artikel 3
Medlemsstaterna får inte, av skäl som sammanhänger med kraven i detta direktiv och dess bilaga, begränsa, hindra eller förbjuda att sådana aerosolbehållare släpps ut på marknaden som uppfyller kraven i detta direktiv och dess bilaga.
2. Kommittén skall själv fastställa sin arbetsordning.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom två månader. Yttranden skall antas med 41 rösters majoritet, varvid medlemsstaternas röster skall vägas enligt förslagets artikel 148.2. Ordföranden får inte rösta.
c) Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen anta förslaget till åtgärder.
b) Symbolen "3" (omvänt epsilon) som bevis för att produkten motsvarar kraven i detta direktiv.
e) Innehållets nettovikt och -volym.
Medlemsstaterna skall vidta nödvändiga åtgärder för att förhindra att märken eller påskrift som kan förväxlas med symbolen "3" (omvänt epsilon) används på aerosolbehållare.
2. Kommissionen skall inom sex veckor rådfråga berörda medlemsstater och därefter utan dröjsmål avge sitt yttrande och vidta lämpliga åtgärder.
1. Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv inom 18 månader efter dagen för anmälan och skall genast underrätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 43 och 100 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
Det är följaktligen lämpligt att harmonisera denna sektor som hittills har omfattats av nationell lagstiftning.
Det är lämpligt att tillåta att medlemsstaterna antar bestämmelser som underlättar plombering av små förpackningar med utsäde av stråsäd, utsädespotatis och utsäde av olje- och spånadsväxter.
Artikel 1
- Annat frö än monogermt frö eller tekniskt monogermfrö (precisionsfrö): högsta nettovikt 10 kg, exklusive, i förekommande fall, pesticider i pulverform, pelleteringsmedel eller andra fasta tillsatser."
3. Medlemsstaterna skall kräva att EEG-småförpackningar plomberas på sådant sätt att plomberingen skadas och inte kan anbringas på nytt när förpackningen öppnats. Förpackningar får inte omplomberas, varken en eller flera gånger, annat än under officiell övervakning.
"1. Medlemsstaterna skall kräva att förpackningar med basutsäde och certifikatutsäde, förutom då utsäde av den sistnämnda kategorin förpackas i EEG-småförpackningar..."
6. Följande artiklar skall läggas till efter artikel 11:
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(1), och
Syftet med den gemensamma jordbrukspolitiken är att uppnå de mål som fastställs i artikel 39 i fördraget. För att stabilisera marknaderna och tillförsäkra den berörda jordbruksbefolkningen en skälig levnadsstandard bör det inom fjäderfäköttsektorn införas bestämmelser om åtgärder för att underlätta anpassningen av utbudet till marknadens behov.
Det är nödvändigt att undvika störningar på gemenskapsmarknaden till följd av utbud på världsmarknaden till extremt låga priser. Därför bör slusspriser fastställas och om anbudspriserna fritt gränsen är lägre än slusspriserna bör importavgifterna höjas med en tilläggsavgift.
Beviljandet av vissa former av stöd kan äventyra förverkligandet av en enhetlig marknad. Följaktligen bör de bestämmelser i fördraget som gör det möjligt att värdera stödåtgärder som beviljats av medlemsstaterna och att förbjuda stödåtgärder som är oförenliga med den gemensamma marknaden göras tillämpliga på marknaden för fjäderfä.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
c) slaktade fjäderfä: döda höns, ankor, gäss, kalkoner och pärlhöns, hela och med eller utan slaktbiprodukter.
3. ätbara slaktbiprodukter enligt punkt 1 b,
6. produkter enligt punkt 1 f.
- Åtgärder för att förbättra kvaliteten.
Allmänna bestämmelser om dessa åtgärder skall antas i enlighet med det förfarande som föreskrivs i artikel 43.2 i fördraget.
Dessa normer får särskilt avse klassificering efter kvalitet och vikt, förpackning, lagring, transport, presentation och märkning.
De produkter som anges i artikel 1.1 skall vid import till gemenskapen beläggas med en importavgift som fastställs på förhand för varje kvartal i enlighet med det förfarande som föreskrivs i artikel 17.
Priserna på foderspannmål inom gemenskapen skall fastställas en gång om året för en tolvmånadersperiod som börjar den 1 augusti. Dessa priser skall baseras på tröskelpriserna på sådan spannmål och den månatliga höjningen av dessa priser.
2. Importavgiften för kycklingar skall beräknas på samma sätt som importavgiften för slaktat fjäderfä. Dock skall den kvantitet foderspannmål som skall användas vid beräkningen vara den kvantitet som åtgår till att inom gemenskapen producera en kyckling. Slusspriset skall vara det som gäller för kycklingar.
Artikel 5
3. Koefficienterna som uttrycker de förhållanden som avses i punkt 1 skall fastställas i enlighet med det förfarande som föreskrivs i artikel 17. De uppgifter som används vid fastställande av koefficienterna skall omprövas minst en gång om året.
Rådet skall på förslag av kommissionen och med kvalificerad majoritet anta allmänna tillämpningsföreskrifter för denna artikel.
2. Slusspriserna på slaktat fjäderfä skall utgöras av följande delar: a) Ett belopp som motsvarar världsmarknadspriset på den kvantitet foderspannmål, differentierad med hänsyn till art av fjäderfä, som åtgår till att i tredje land producera 1 kg slaktat fjäderfä.
Vid fastställande av det slusspris som skall gälla från den 1 november, den 1 februari och den 1 maj skall emellertid hänsyn tas till prisutvecklingen på världsmarknaden för foderspannmål endast om priset på kvantiteten foderspannmål uppvisar en minimiavvikelse från det pris som användes vid beräkning av slusspriset för föregående kvartal. De uppgifter som används för att fastställa det standardbelopp som avses i b skall omprövas minst en gång om året.
5. Rådet skall på förslag av kommissionen och med kvalificerad majoritet anta tillämpningsföreskrifter för denna artikel.
2. Importavgiften skall emellertid inte höjas med denna tilläggsavgift när det gäller tredje land som vill och är i stånd att garantera att importpriset till gemenskapen på produkter som har sitt ursprung i och kommer från deras territorium inte kommer att bli lägre än slusspriset för produkten i fråga och att varje snedvridning av handeln kommer att undvikas.
4. Närmare tillämpningsföreskrifter för denna artikel skall antas i enlighet med förfarandet i artikel 17.
1. I den mån det är nödvändigt för att göra det möjligt att exportera de produkter som avses i artikel 1.1 på grundval av världsmarknadspriserna på dessa produkter, får skillnaden mellan världsmarknadspriserna och priserna inom gemenskapen täckas av ett exportbidrag.
Vid fastställande av exportbidraget skall särskild hänsyn tas till behovet av att skapa en balans mellan användningen av gemenskapens basvaror vid framställningen av bearbetade varor för export till tredje land och användningen av produkter från tredje land som förts in enligt bestämmelserna för aktiv förädling.
3. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 17.
Artikel 11
- Införande av tullar eller avgifter med motsvarande verkan.
1. Om gemenskapsmarknaden för en eller flera av de produkter som anges i artikel 1.1, till följd av import eller export är utsatt för eller hotas av allvarliga störningar som kan äventyra de mål som fastställs i artikel 39 i fördraget, får lämpliga åtgärder avseende handeln med tredje land vidtas till dess att störningen eller hotet om störning har upphört.
3. En medlemsstat får hänskjuta kommissionens beslut om åtgärder till rådet inom tre arbetsdagar efter det att beslutet meddelades. Rådet skall sammanträda utan dröjsmål och får med kvalificerad majoritet ändra eller upphäva åtgärderna i fråga.
Artikel 14
Medlemsstaterna och kommissionen skall till varandra överlämna sådana uppgifter som är nödvändiga för att tillämpa denna förordning. Bestämmelser om överlämnande och spridning av sådana uppgifter skall fastställas i enlighet med det förfarande som föreskrivs i artikel 17.
2. Inom kommittén skall medlemsstaternas röster vägas enligt artikel 148.2 i fördraget. Ordföranden får inte rösta.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med en majoritet av 41 röster.
Artikel 18
Om inte annat följer av denna förordning, skall artikel 92 94 i fördraget gälla för produktionen av och handeln med de produkter som anges i artikel 1.1.
Artikel 21
1. Rådets förordning nr 123/67/EEG(5) av den 13 juni 1967 om den gemensamma organisationen av marknaden för fjäderfäkött, senast ändrad genom rådets beslut av den 1 januari 1973(6) om anpassning av dokumenten avseende de nya medlemsstaternas anslutning till Europeiska gemenskaperna, upphävs härmed.
Artikel 23
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
Tillnärmningen av den nationella lagstiftningen om motorfordon innefattar medlemsstaternas ömsesidiga erkännande av de kontroller som utförs av var och en av dem på grundval av gemensamma bestämmelser. För att ett sådant system skall bli framgångsrikt måste dessa bestämmelser tillämpas av alla medlemsstater från samma datum.
I detta direktiv avses med fordon varje motorfordon som är avsett att användas på väg, med eller utan karosseri, med minst fyra hjul och som är konstruerade för en högsta hastighet som överstiger 25 km/tim och släpvagnar till dessa fordon, dock med undantag av spårbundna fordon, traktorer och maskiner för jordbruk eller skogsbruk samt andra motorredskap.
Artikel 3
De ändringar som är nödvändiga för att anpassa kraven i bilagan till den tekniska utvecklingen skall antas enligt det förfarande som beskrivs i artikel 13 i direktiv 70/156/EEG.
Artikel 6
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 100 och 235 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
Inom detta område finns det vissa lagar och andra författningar i medlemsstaterna som direkt påverkar den gemensammamarknadens funktion. Fördraget ger dock inte alla de befogenheter som är nödvändiga för att vidta åtgärder.
Det bör föreskrivas att badvatten under vissa förhållanden skall anses uppfylla de relevanta parametervärdena, även om en viss procent av proven som tagits under badsäsongen inte överensstämmer med de gränsvärden som anges i bilagan.
Allmänhetens intresse för miljön och en förbättrad miljökvalitet ökar. Allmänheten bör därför få objektiv information om kvaliteten på badvatten.
- badning inte är förbjuden och traditionellt utövas av ett stort antal badare,
Artikel 2
1. Medlemsstaterna skall för alla badplatser eller för varje enskild badplats fastställa de värden som skall gälla för badvatten i fråga om de parametrar som anges i bilagan.
Artikel 5
- vattnet inte avviker från de relevanta parametervärdena med mer än 50 % utom för mikrobiologiska parametrar, pH och löst syre,
Artikel 8
Naturlig berikning avser den process genom vilken en viss vattenmassa, utan mänsklig påverkan, tillförs vissa ämnen ur marken.
Artikel 9
De skall antas i enlighet med det förfarande som fastställs i artikel 11.
3. a) Kommissionen skall själv anta förslaget om det är förenligt med kommitténs yttrande.
Artikel 12
Artikel 13
Artikel 14
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(1),
Harmonisering av lagar och andra författningar som avser dessa mätdon är också väsentlig som ett komplement till gällande bestämmelser om metoder att bestämma alkoholhalt utgående från mätresultat, så att alla risker avlägsnas för flertydighet i eller ifrågasättande av resultaten av sådana mätningar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 4
Artikel 5
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av kommissionens förslag,
med beaktande av följande: I artikel 5.1 b andra strecksatsen i förordning (EEG) nr 543/69 föreskrivs att förare av ett fordon som är avsett för transport av gods med en högsta tillåtna vikt över 7,5 metriska ton och som omfattas av förordningen, måste, om vederbörande inte har fyllt 21 år, inneha ett intyg om yrkeskompetens som är erkänt i en av medlemsstaterna. Intyget skall styrka att föraren har genomgått utbildning för förare av fordon som är avsedda för godstransporter på väg.
Artikel 1
3. Varje medlemsstat får kräva att förare som utför inrikestransporter på dess territorium och förare som utför internationella transporter med fordon registrerade i denna stat skall genomgå en mer omfattande utbildning än den som beskrivs i bilagan. Denna utbildning kan utgöras av utbildning som redan finns eller av utbildning som en medlemsstat beslutar införa i framtiden.
2. Rättigheter som förvärvats med stöd av de föreskrifter som avses i punkt 1 innan de nationella lagar och andra författningar som har antagits till följd av detta direktiv träder i kraft, skall förbli giltiga på samma sätt som utbildningsintyg, som utfärdats enligt detta direktiv.
2. Varje medlemsstat skall tillställa kommissionen prov på de utbildningsintyg eller likvärdiga dokument som staten inför för tillämpning av artikel 2.1. Kommissionen skall snarast vidarebefordra dessa underlag till de övriga medlemsstaterna.
RÅDETS FÖRORDNING (EEG) nr 2566/76 av den 20 juli 1976 om godkännande av avtalet i form av skriftväxling rörande ändringar i tabell I och II i bilaga till protokoll 2 till avtalet mellan Europeiska ekonomiska gemenskapen och Schweiz
med beaktande av kommissionens rekommendation, och
Härmed godkänns på gemenskapens vägnar avtalet i form av skriftväxling om ändringar i tabell I och II i bilaga till protokoll 2 till avtalet mellan Europeiska ekonomiska gemenskapen och Schweiz.
Rådets ordförande bemyndigas att utse den person som är behörig att med bindande verkan för gemenskapen underteckna avtalet.
RÅDETS ANDRA DIREKTIV av den 13 december 1976 om samordning av de skyddsåtgärder som krävs i medlemsstaterna av de i artikel 58 andra stycket i fördraget avsedda bolagen i bolagsmännens och tredje mans intressen när det gäller att bilda ett aktiebolag samt att bevara och ändra dettas kapital, i syfte att göra skyddsåtgärderna likvärdiga (77/91/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: Eftersom aktiebolagen spelar en framträdande roll i medlemsstaternas näringsliv och deras verksamhet ofta sträcker sig utöver de nationella gränserna, är det i fråga om dessa bolag särskilt viktigt att fortsätta den samordning som föreskrivs i artikel 54.3 g i fördraget och i Allmänna handlingsprogrammet för upphävande av begränsningar av etableringsfriheten och som inleddes med direktiv 68/151/EEG (3).
Sådana gemenskapsregler om att bevara det kapital som utgör borgenärernas säkerhet skall antas, som särskilt förbjuder en minskning av kapitalet genom utdelning till aktieägarna och begränsar bolagens möjligheter att förvärva egna aktier.
Artikel 1
- I Italien: la società per azioni.
- som inbjuder allmänheten att förvärva aktier i bolaget, och
Bolagsordningen eller stiftelseurkunden skall alltid innehålla minst följande uppgifter: a) bolagsform och firma;
- om bolaget har ett "auktoriserat" kapital, storleken av detta och det tecknade kapitalet vid bolagsbildningen eller då bolaget får tillstånd att börja sin verksamhet och vid varje ändring av det "auktoriserade" kapitalet, dock med förbehåll för vad som gäller enligt artikel 2.1 e i direktiv 68/151/EEG;
Artikel 3
c) antalet tecknade aktier utan nominellt belopp, om den nationella lagstiftningen tillåter att sådana aktier ges ut;
f) huruvida aktierna är ställda till viss man eller till innehavaren, om den nationella lagstiftningen tillåter båda formerna, och bestämmelser om hur aktierna omvandlas från den ena formen till den andra, om inte förfarandet är reglerat i lag eller annan författning;
i) identiteten hos de fysiska eller juridiska personer eller bolag av vilka eller i vilkas namn bolagsordningen eller stiftelseurkunden eller, om bolagsbildningen inte sker i ett sammanhang, utkasten till dessa handlingar har undertecknats;
Artikel 4
Artikel 5
3. När förordnandet om upplösning har meddelats, skall bolaget träda i likvidation.
Med en europeisk beräkningsenhet avses en sådan enhet som har bestämts genom kommissionens beslut nr 3289/75/EKSG (4). Som motvärde i nationell valuta gäller första gången motvärdet den dag då detta direktiv antas.
Det tecknade kapitalet får endast bestå av tillgångar som kan värderas ekonomiskt. I dessa tillgångar får dock inte inräknas åtaganden att utföra arbete eller att tillhandahålla tjänster.
2. Medlemsstaterna kan dock tillåta att de som yrkesmässigt åtar sig att placera aktier får betala mindre än fullt belopp för de aktier som de tecknar i ett sådant sammanhang.
2. Aktier som har getts ut mot apportegendom innan bolaget bildas eller får tillstånd att börja sin verksamhet skall vara fullt betalda inom fem år från bolagsbildningen eller tillståndet att börja verksamheten.
2. Sakkunnigutlåtandet skall minst beskriva apportegendomen samt ange vilka värderingsmetoder de sakkunniga har använt och huruvida de därvid beräknade värdena åtminstone motsvarar antal, nominellt värde eller, i avsaknad av sådant värde, bokfört parivärde och i förekommande fall överkurs i fråga om de aktier för vilka apportegendomen utgör vederlag.
b) avståendet har offentliggjorts enligt punkt 3;
e) det vid d angivna ansvaret har offentliggjorts enligt punkt 3;
1. Om ett bolag inom en tid som av den nationella lagstiftningen skall bestämmas till minst två år från det att bolagets bildades eller tilläts att börja sin verksamhet förvärvar tillgångar från en person eller ett bolag som avses i artikel 3 i mot ett vederlag som motsvarar minst en tiondel av det tecknade kapitalet, skall förvärvet granskas och offentliggöras enligt artikel 10 samt underställas bolagsstämman för godkännande.
Artikel 12
Om ett bolag av annat slag ombildas till aktiebolag skall medlemsstaterna, i avvaktan på en senare samordning av den nationella lagstiftningen, se till att minst de skyddsåtgärder som föreskrivs i artiklarna 2-12 iakttas.
Artikel 15
c) Det belopp som delas ut till aktieägarna får inte överstiga vinsten för det senast avslutade räkenskapsåret med tillägg för balanserad vinst och belopp från reserver som får användas för detta ändamål samt med avdrag för balanserad förlust och belopp som enligt lag eller bolagsordning har avsatts till reserver.
b) det belopp som skall delas ut får inte överstiga den vinst som har uppkommit efter det senaste räkenskapsår för vilket årsbokslut har upprättats, med tillägg för balanserad vinst och belopp från reserver som får användas för detta ändamål samt med avdrag för balanserad förlust och belopp som enligt lag eller bolagsordning skall föras över till reserver.
I denna punkt anses som förvaltningsbolag med fast kapital endast bolag: - som uteslutande har till föremål för sin verksamhet att placera sina medel i olika värdepapper, olika fastigheter eller andra tillgångar i det enda syftet att sprida investeringsriskerna och låta resultatet av kapitalförvaltningen komma aktieägarna till godo, och
b) får denna inte tillåta ett bolag som nu avses och vars nettotillgångar understiger det i punkt 1 a nämnda beloppet att dela ut medel till aktieägarna, om enligt årsredovisningen för det senaste räkenskapsåret summan av bolagets samtliga tillgångar på bokslutsdagen understiger eller till följd av utdelningen skulle komma att understiga en och en halv gånger beloppet av bolagets samtliga skulder enligt årsredovisningen;
En utdelning i strid med artikel 15 skall återbetalas av de aktieägare som har mottagit denna, om bolaget visar att aktieägarna kände till att utdelningen var olaglig eller att de med hänsyn till omständigheterna inte kunde vara okunniga om det.
2. Gränsen för betydande förlust enligt punkt 1 får i medlemsstaternas lagstiftning inte sättas högre än till hälften av det tecknade kapitalet.
2. Om aktierna i ett bolag har tecknats av någon i eget namn men för bolagets räkning, skall denne anses ha tecknat aktierna för egen räkning.
Artikel 19
c) Förvärvet får inte medföra att värdet av nettotillgångarna understiger det belopp som anges i artikel 15.1 a.
3. Medlemsstaterna behöver inte tillämpa punkt 1 a första meningen på aktier som förvärvas av bolaget, direkt eller av någon som handlar i eget namn men för bolagets räkning, för att fördelas bland de anställda i bolaget eller ett detta närstående bolag. Sådana aktier skall fördelas inom 12 månader från förvärvet.
b) aktier som förvärvas som ett led i en allmän förmögenhetsövergång;
e) aktier som förvärvas från en aktieägare på grund av bristande betalning av aktierna;
h) helt betalda aktier som har getts ut av ett förvaltningsbolag med fast kapital enligt artikel 15.4 andra stycket och som på placerarnas begäran förvärvas av detta bolag eller av ett detta närstående bolag. Artikel 15.4 a skall därvid tillämpas. Ett sådant förvärv får inte medföra att nettotillgångarna understiger det tecknade kapitalet ökat med de reserver som enligt lag inte får delas ut.
Artikel 21
1. Om lagstiftningen i en medlemsstat tillåter ett aktiebolag att förvärva egna aktier, direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall lagstiftningen för det fortsatta innehavet av aktierna alltid kräva att minst följande villkor iakttas:
b) antal och nominellt värde eller, i avsaknad av sådant värde, bokfört parivärde beträffande de aktier som har förvärvats och avyttrats under räkenskapsåret samt den andel av det tecknade kapitalet som dessa aktier utgör;
Artikel 23
3. Punkt 1 tillämpas inte på åtgärder som vidtas för att aktier skall förvärvas enligt artikel 20.1 h.
2. Medlemsstaterna behöver inte tillämpa punkt 1 på åtgärder i en banks eller något annat finansinstituts löpande verksamhet.
2. Bolagsordningen, stiftelseurkunden eller bolagsstämman, vilken senares beslut skall offentliggöras enligt punkt 1, får dock ge bemyndigande om att öka det tecknade kapitalet upp till ett högsta belopp som fastställs med hänsyn till eventuella lagregler om sådant högsta belopp. Inom ramen för det fastställda beloppet beslutar det bemyndigade bolagsorganet i förekommande fall om ökning av det tecknade kapitalet. Bemyndigandet gäller i högst fem år och kan förlängas av bolagsstämman en eller flera gånger med högst fem år varje gång.
Artikel 26
1. Om aktier ges ut mot apportegendom som ett led i ökningen av det tecknade kapitalet, skall aktierna vara helt betalda inom fem år från beslutet om ökning av det tecknade kapitalet.
Artikel 28
1. Vid varje ökning av det tecknade kapitalet, som skall betalas med pengar, skall aktierna med företrädesrätt erbjudas aktieägarna i förhållande till den andel av kapitalet som deras aktier representerar.
3. Erbjudandet om företrädesrätt och den tid inom vilken denna rätt får utnyttjas skall offentliggöras i den nationella tidning som har utsetts i överensstämmelse med direktiv 68/151/EEG. Lagstiftningen i en medlemsstat behöver dock inte föreskriva ett offentliggörande, om alla bolagets aktier är ställda till viss man. I sådant fall skall samtliga aktieägare underrättas skriftligen. Den tid inom vilken företrädesrätten skall utnyttjas får inte understiga 14 dagar från det att erbjudandet offentliggörs eller den skriftliga underrättelsen avsänds.
6. Punkterna 1-5 tillämpas vid emission av alla värdepapper som kan bytas ut mot aktier eller som är förenade med teckningsrätt till aktier, men inte vid själva utbytet av värdepapperen eller vid utnyttjandet av teckningsrätten.
Artikel 31
1. Om det tecknade kapitalet sätts ned har åtminstone de borgenärer, vilkas fordringar har uppkommit före offentliggörandet av beslutet om nedsättningen, rätt att minst få säkerhet för de fordringar som inte är förfallna till betalning vid offentliggörandet. Lagstiftningen i medlemsstaterna bestämmer under vilka förutsättningar denna rätt får utövas. Lagstiftningen får utesluta rätten endast om en borgenär har tillfredsställande säkerhet eller sådan inte behövs med hänsyn till bolagets ställning.
Artikel 33
Artikel 34
Om lagstiftningen i en medlemsstat tillåter att det tecknade kapitalet helt eller delvis löses in utan att kapitalet sätts ned, skall lagstiftningen minst kräva att följande villkor är uppfyllda: a) Om bolagsordningen eller stiftelseurkunden ger möjlighet till inlösen skall beslut om inlösen fattas av bolagstämman, som minst skall iaktta de allmänna villkoren för beslutförhet och majoritet. Om bolagsordningen eller stiftelseurkunden inte ger möjlighet till inlösen skall beslut om inlösen fattas av bolagstämman, som i så fall minst skall iaktta villkoren för beslutförhet och majoritet enligt artikel 40. Beslutet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
Artikel 36
c) Det bolagsorgan som beslutar om tvångsindragningen skall bestämma villkor och sätt för denna, om inte det har skett redan i bolagsordningen eller stiftelseurkunden.
2. Artikel 30 första stycket samt artiklarna 31, 33 och 40 tillämpas inte i de fall som avses i punkt 1.
2. Artikel 32 tillämpas utom i fråga om helt betalda aktier som har förvärvats utan vederlag eller med medel som får delas ut enligt artikel 15.1; i dessa fall skall ett belopp som motsvarar det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet för samtliga indragna aktier föras över till en reserv. Utom vid nedsättning av det tecknade kapitalet får denna reserv inte delas ut till aktieägarna; den får endast användas för att täcka en inträffad förlust eller för att öka det tecknade kapitalet genom överföring av reserver, i den mån medlemsstaterna tillåter en sådan åtgärd.
Om det finns flera slag av aktier skall i de fall som avses i artikel 35, artikel 36.1 b och artikel 37.1 bolagsstämmans beslut om inlösen av det tecknade kapitalet eller nedsättning av detta genom indragning av aktier bli föremål för en särskild omröstning minst för varje kategori av aktieägare vilkas rätt berörs av åtgärden.
b) aktierna skall vara helt betalda;
e) ett belopp som motsvarar det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet av alla återköpta aktier skall föras över till en reserv som inte får delas ut till aktieägarna i annat fall än då det tecknade kapitalet sätts ned; denna reserv får endast användas för att öka det tecknade kapitalet genom överföring av reserver;
h) återköpet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
2. Medlemsstaternas lagstiftning får dock föreskriva att enkel majoritet av rösterna enligt punkt 1 är tillräcklig, om minst hälften av det tecknade kapitalet är företrätt.
2. Medlemsstaterna får underlåta att tillämpa artikel 19.1 a första ledet samt artiklarna 30, 31 och 36-39 på bolag som bildas enligt särskild lagstiftning och som vid sidan av "kapitalaktier" ger ut "arbetsaktier" till förmån för de anställda som ett kollektiv, vilket på bolagsstämman företräds av fullmäktige med rösträtt.
Artikel 43
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
Om dessa skillnader skall kunna avlägsnas, vilket skulle leda till en ökning av jordbrukets produktivitet på området, måste handeln med alla renrasiga avelsdjur inom gemenskapen gradvis göras fri. En fullständig frihet i handeln förutsätter en ytterligare harmonisering, särskilt i fråga om godkännande för avel.
Det måste säkerställas att import av renrasiga avelsdjur av nötkreatur från icke-medlemsländer inte får ske på villkor som är mindre stränga än de som tillämpas inom gemenskapen.
I detta direktiv används följande beteckningar med de betydelser som här anges: a) renrasigt avelsdjur av nötkreatur: varje nötkreatur vars föräldrar samt far- och morföräldrar är införda eller registrerade i en stambok för samma ras och som självt är infört i eller är registrerat och berättigat till införande i en sådan stambok. b) stambok: varje bok, förteckning eller dataregister
Artikel 2
- Upprättande av stamböcker förutsatt att de uppfyller kraven enligt artikel 6.
Artikel 3
Artikel 4
Medlemsstaterna får kräva att renrasiga avelsdjur av nötkreatur samt sperma och embryon från sådana djur vid handel inom gemenskapen skall åtföljas av ett härstamningsintyg som har utformats enligt det förfarande som fastställs i artikel 8, särskilt då det gäller resultat från husdjurskontroll och avelsprövningar.
- Metoder för husdjurskontroll och avelsprövningar samt metoder för beräkning av djurens avelsvärde.
- Vilka uppgifter som skall anges i härstamningsintyget.
c) skall upprättandet av nya stamböcker även fortsättningsvis uppfylla de villkor som för närvarande gäller i varje medlemsstat.
Medlemsstaterna får inte tillåta import av renrasiga avelsdjur av nötkreatur från icke-medlemsländer om inte djuren åtföljs av ett härstamningsbevis som intygar att de är införda eller registrerade i en stambok i det exporterande icke-medlemslandet. Bevis måste framläggas på att djuren är införda i eller registrerade och berättigade till införande i en stambok i gemenskapen.
2. Inom kommittén skall medlemsstaternas röster vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas och tillämpa dem omedelbart såvida inte rådet med enkel majoritet har avvisat förslaget.
Artikel 10
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning nr 171/67/EEG av den 27 juni 1967 om exportbidrag och avgifter på olivolja(4), senast ändrad genom förordning (EEG) nr 2429/72(5), särskilt artikel 11 i denna, och
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för oljor och fetter.
Artikel 2 i förordning (EEG) nr 616/72 skall ändras på följande sätt:
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Villkoren för certifiering av majsutsäde bör anpassas till befintliga internationella program för sortcertifiering av utsäde.
Vissa standarder som skall uppfyllas av utsäde av ris bör anpassas till den utsädeskvalitet som normalt uppnås.
KOMMISSIONENS DIREKTIV av den 19 maj 1978 om anpassning till teknisk utveckling av rådets direktiv 76/114/EEG om tillnärmning av medlemsstaternas lagstiftning om föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt på motorfordon och släpvagnar till dessa fordon (78/507/EEG)
med beaktande av rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(1), i dess lydelse enligt anslutningsakten och särskilt artiklarna 11, 12 och 13 i denna,
Bestämmelserna i detta direktiv har tillstyrkts av Kommittén för anpassning till teknisk utveckling av direktiv om avskaffande av tekniska handelshinder inom motorfordonssektorn.
Bilagan till direktiv 76/114/EEG ändras enligt bilagan till detta direktiv.
- förbjuda att fordon tas i bruk
- Medlemsstaterna får vägra att bevilja nationellt typgodkännande för en typ av fordon för vilken föreskrivna skyltar och märkningar samt deras placering och fastsättning inte överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
Medlemsstaterna skall senast den 1 oktober 1978 sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv och skall genast underrätta kommissionen om detta.
RÅDETS FÖRORDNING (EEG) nr 1883/78 av den 2 augusti 1978 om allmänna bestämmelser för finansiering av interventioner genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ)
med beaktande av rådets förordning (EEG) nr 729/70 av den 21 april 1970 om finansiering av den gemensamma jordbrukspolitiken(1), senast ändrad genom förordning (EEG) nr 2788/72(2), särskilt artikel 3.2 i denna,
med beaktande av följande: I enlighet med artikel 3.2 i förordning (EEG) nr 729/70 bör allmänna bestämmelser för gemenskapsfinansiering av interventioner fastställas.
För de interventionsåtgärder för vilka ett belopp per enhet inte bestäms inom ramen för den gemensamma organisationen av marknaderna, bör grundläggande regler fastställas särskilt vad avser metoden för bestämning av de belopp som skall finansieras, finansieringen av utgifter som följer av att nödvändiga medel binds upp för interventionsköp av produkter, värderingen av lager som skall överföras från ett räkenskapsår till nästföljande och finansieringen av utgifter i samband med lagring och vid behov i samband med bearbetning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
När det inom ramen för den gemensamma organisationen av marknaden inte fastställs ett belopp per enhet för en interventionsåtgärd, skall denna finansieras av garantisektionen vid EUGFJ i enlighet med de bestämmelser som anges i artikel 4 8.
Artikel 5
Materiella åtgärder i samband med lagring och, i förekommande fall, bearbetning av interventionsprodukter, skall finansieras av garantisektionen vid EUGFJ med hjälp av schablonbelopp som är enhetliga inom hela gemenskapen och som skall fastställas enligt förfarandet i artikel 13 i förordning (EEG) nr 729/70, vid behov efter granskning av ärendet i den berörda förvaltningskommittén.
Artikel 8
Artikel 9
Förordning (EEG) nr 2824/72 upphör att gälla.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Med hänsyn till vunna erfarenheter och den tekniska utvecklingen är det nu möjligt att göra kraven strängare och att anpassa dem bättre till faktiska provningsförhållanden.
Artikel 1
Artikel 2
- förbjuda att fordon tas i bruk,
- inte längre utfärda det exemplar av det intyg som anges i sista strecksatsen i artikel 10.1 i direktiv 70/156/EEG med avseende på en fordonstyp vars bromsutrustning inte överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv,
4. Utan hinder av punkterna 1-3 skall medlemsstaterna tillämpa bestämmelserna i punkt 1.2.1 i bilaga 4 till direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv, endast från den 1 oktober 1983.
KOMMISSIONENS FÖRORDNING (EEG) nr 883/79 av den 3 maj 1979 om ändring av förordning (EEG) nr 2960/77 om närmare bestämmelser för försäljning av olivolja som innehas av interventionsorgan
med beaktande av av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(1), senast ändrad genom förordning (EEG) nr 590/79(2), särskilt artikel 12.4 i denna, och
För att underlätta avhämtningen av de sålda oljorna bör avhämtningstidens längd ändras genom att den anpassas efter det tilldelade partiets storlek.
Artikel 1
2. Artikel 6 andra stycket skall ersättas med följande:
4. Följande stycke skall läggas till i artikel 11.1:
2. Om det preliminära beloppet inte betalas inom den tid som anges i artikel 13.1, skall köpet automatiskt upphävas. I sådana fall skall den säkerhet som avses i artikel 8 förverkas.
Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av följande: Enligt artikel 227.2 tredje stycket i fördraget skall gemenskapens institutioner inom ramen för den ordning som anges i fördraget sörja för att den ekonomiska och sociala utvecklingen i de franska utomeuropeiska departementen möjliggörs.
Artikel 1
Artikel 2
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
När det gäller exportavgifterna kan det förekomma att avgiftsbeloppet är lägre än det belopp med vilket justeringen skall göras. För att undvika att företagen blir olika behandlade måste därför ett tillägg göras till den aktuella förordningen, enligt vilket skillnaden skall betraktas som ett exportbidrag som ges till den berörda parten i stället för utkrävandet av exportavgiften.
Artikel 1
"Om exportavgiften är lägre än det belopp med vilket den skall justeras, skall skillnaden mellan de två beloppen betraktas som ett exportbidrag som skall ges till den berörda parten. I sådana fall skall exportavgiften inte betalas."
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
Av detta skäl bör direktiv 77/541/EEG ändras.
"Artikel 9
"3.1 Fordonsutrustning
b) Avsnitt 3.1.1 skall ersättas med följande:
Med avseende på bilbältena skall vindrutan anses vara en del av referenszonen när den kan komma i statisk kontakt med provningsutrustningen enligt den metod som beskrivs i bilaga 2 till direktiv 74/60/EEG."
d) Lägg till ett nytt avsnitt 3.1.5 enligt följande:
Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv på samma dag som planerats för ikraftträdandet av bestämmelserna som krävs för att följa det direktiv som skall antas efter detta direktiv enligt artikel 10 i direktiv 77/541/EEG så att kraven i bilagorna till det sistnämnda direktivet kan anpassas till den tekniska utvecklingen. De skall genast underrätta kommissionen om detta.
RÅDETS DIREKTIV av den 19 oktober 1981 om ändring med anledning av Greklands anslutning av direktiv 79/869/EEG om mätmetoder samt provtagnings- och analysfrekvenser avseende ytvatten för dricksvattenframställning i medlemsstaterna (81/855/EEG)
med beaktande av kommissionens förslag,
I enlighet med artikel 198 första stycket i fördraget har rådet samrått med Ekonomiska och sociala kommittén om kommissionens förslag. Kommittén hade inte möjlighet att avge sitt yttrande inom den tidsgräns som rådet hade fastställt. Enligt artikel 198 andra stycket i fördraget skall avsaknaden av ett yttrande inte hindra rådet från att vidta åtgärder. Eftersom det är önskvärt att de nödvändiga ändringarna antas snabbt finner rådet det angeläget att utnyttja denna möjlighet.
I artikel 11.2 i direktiv 79/869/EEG skall "41" ersättas med "45".
Artikel 3
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(), och
Konventionens lydelse ändrades därför genom förordning (EEG) nr 653/80() men tillämpningen av ändringen var begränsad till och med den 31 december 1980 eftersom den var avsedd som en interimsåtgärd i enlighet med artikel 103 i fördraget.
Artikel 1
med beaktande av Europaparlamentets yttrande (),
Informationssystemets undersökningsområde måste bestå av alla jordbruksföretag av en viss ekonomisk storlek, oberoende av om jordbrukaren åtar sig annat arbete utanför företaget.
Det nationella samordningsorganet måste ha en nyckelroll i handhavandet av informationssystemet. I detta syfte bör det förses med nya uppgifter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2) Artikel 4 skall ersättas med följande:
2. För att bli behörigt som rapporterande företag skall ett jordbruksföretag
c) tillsammans med de övriga företagen och på områdesnivå vara representativt för undersökningsområdet.
3) Artikel 5 skall ersättas med följande:
2. Den nationella kommittén skall ha ansvaret för valet av rapporterande företag. För detta ändamål skall dess uppgifter framför allt omfatta godkännandet av
3. Ordföranden i den nationella kommittén skall utses av medlemsstaten bland medlemmarna i denna kommitté.
Den regionala kommittén skall särskilt ha som uppgift att arbeta med det samordningsorgan som anges i artikel 6 för att välja ut rapporterande företag.
"Artikel 6
b) att utarbeta och till den nationella kommittén överlämna för godkännande och därefter till kommissionen överlämna
c) att sammanställa
e) att överlämna de ifyllda företagsredovisningarna till kommissionen omedelbart efter kontrollen,
5) Artikel 9.2 andra stycket skall upphöra att gälla.
Denna begäran om uppgifter till den nationella kommittén, de regionala kommittéerna eller bokföringsbyråerna och svaren på dessa skall meddelas skriftligen genom samordningsorganet."
med beaktande av Europaparlamentets yttrande (), och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"Grekland
Denna förordning träder i kraft dagen efter dess offentliggörande i Europeiska gemenskapernas officiella tidning.
med beaktande av rådets direktiv 69/208/EEG av den 30 juni 1969 om saluföring av utsäde av olje- och spånadsväxter(), senast ändrat genom direktiv 81/126/EEG, särskilt artikel 20 a i detta, och
Det har i det nuvarande läget inte varit möjligt att, i fråga om solroshybrider, föreskriva om en harmonisering inom gemenskapen av de minimistandarder för sortrenhet som grödor och utsäde måste motsvara. Ett försök skall dock göras före den 1 juli 1983 att upprätta sådana standarder i syfte att uppnå en harmonisering.
Artikel 1
2. I andra och tredje meningen i punkt 4 skall orden "Raphanus sativus ssp. oleifera" utgå.
1. Punkt 1 i avsnitt I skall ersättas med följande:
Bilaga 1 till direktiv 69/208/EEG ändras på följande sätt:
- en per 10 m² vid produktion av certifikatutsäde."
Punkt 1 i avsnitt I skall ersättas med följande:
Lägsta sortrenhet skall främst undersökas vid fältbesiktningar som utförs enligt de villkor som fastställts i bilaga 1."
Artikel 6 I artikel 2.1 första strecksatsen i direktiv 78/388/EEG skall "den 1 januari 1982" ersättas med "vid ett datum som kommer att fastställas senare".
- bestämmelserna i artikel 5 och 6, med verkan från och med den 1 januari 1982,
2. Medlemsstaterna skall se till att utsäde inte underkastas några begränsningar av saluföringen till följd av olika datum för genomförandet av detta direktiv i enlighet med punkt 1, tredje strecksatsen.
med beaktande av protokollet om immunitet och privilegier för Europeiska gemenskaperna, särskilt artikel 13 i detta,
EUROPEISKA GEMENSKAPERNAS RÅD HAR FATTAT DETTA BESLUT
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
b) det område där motåtgärden skall tillämpas,
e) den tid under vilken motåtgärden skall tillämpas,
Det står medlemsstaterna fritt att ensidigt tillämpa nationella motåtgärder.
RÅDETS ÅTTONDE DIREKTIV av den 10 april 1984 grundat på artikel 54.3 g i fördraget, om godkännande av personer som har ansvar för lagstadgad revision av räkenskaper (84/253/EEG)
med beaktande av kommissionens förslag (1),
med beaktande av följande: Enligt direktiv 78/660/EEG (4) skall årsbokslutet i vissa företagsformer revideras av en eller flera personer som är behöriga att företa sådan revision. Endast företag som anges i artikel 11 i det direktivet får undantas från revisionen.
Genom en yrkesexamen måste en hög nivå garanteras när det gäller de teoretiska kunskaper och den förmåga att praktiskt tillämpa kunskaperna som behövs för en lagstadgad revision av räkenskaper.
Medlemsstaterna får godkänna såväl fysiska personer som revisionsbolag, vilka kan vara juridiska personer eller andra former av bolag eller sammanslutningar.
Om en medlemsstat då detta direktiv antas erkänner som revisorer vissa kategorier av fysiska personer vilka uppfyller i direktivet uppställda krav men vilkas yrkesexamen ligger på en lägre nivå än avslutad högskoleutbildning, bör denna medlemsstat i fortsättningen på vissa villkor och till dess ytterligare samordning sker få särskilt godkänna sådana personer att utföra lagstadgad revision i bolag och företagsgrupper av begränsad storlek. En förutsättning bör vara att medlemsstaten inte har utnyttjat de möjligheter till undantag från kravet på lagstadgad revision som lämnas i gemenskapsdirektiven om årsbokslut och sammanställt bokslut.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. De samordningsåtgärder som föreskrivs i detta direktiv skall vidtas i fråga om sådana lagar och andra författningar i medlemsstaterna som avser personer, vilka skall: a) utföra lagstadgad granskning av bolags och andra företags årsbokslut samt verifiera att innehållet i förvaltningsberättelserna är förenligt med årsboksluten, förutsatt att sådan granskning och verifiering föreskrivs i gemenskapsrätten,
AVSNITT II Regler om godkännande
b) Revisionsbolag som uppfyller minst följande villkor: i) De fysiska personer som på revisionsbolagets vägnar utför lagstadgad revision av de i artikel 1 angivna handlingarna skall uppfylla minst de i artikel 3-19 angivna villkoren; medlemsstaterna får föreskriva att sådana fysiska personer även skall vara godkända.
Med förbehåll för vad som gäller enligt artikel 14.2 skall godkännandet av ett revisionsbolag återkallas när något av kraven i b inte längre är uppfyllt. Medlemsstaterna får dock förordna om en frist på högst två år för att uppfylla kraven i b ii och iii.
Myndigheterna i en medlemsstat skall godkänna endast personer som har ett gott anseende och inte utövar någon form av verksamhet som enligt medlemsstatens lagar är oförenlig med lagstadgad revision av de i artikel 1.1 angivna handlingarna.
Artikel 5
- extern redovisning,
- intern revision och kontroll,
b) i den utsträckning det har betydelse för revisionen: - associationsrätt,
- civil- och handelsrätt,
- företagsekonomi, nationalekonomi och finansiering,
Artikel 7
Artikel 8
Artikel 9
Artikel 10
Artikel 11
2. Artikel 3 skall tillämpas.
2. Inträder en fysisk person i en av staten erkänd yrkesförening får detta anses som ett godkännande genom förvaltningsbeslut av behörig myndighet enligt punkt 1, om inträdet enligt lagstiftningen i den staten ger föreningsmedlemmen rätt att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna.
Artikel 14
3. Fysiska personer som till dess de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas utför lagstadgad revision av de i artikel 1.1 angivna handlingarna för ett revisionsbolags räkning, får därefter meddelas tillstånd att fortsätta att utföra sådan revision även om de inte uppfyller alla villkor i detta direktiv.
Artikel 16
2. Artikel 3 skall tillämpas.
Artikel 20
Om bolaget ingår i en grupp av företag vars räkenskaper skall sammanställas och som överskrider gränserna för två av de tre kriterierna i artikel 27 i direktiv 78/660/EEG, får dock inte sådana personer utföra lagstadgad revision i bolaget av de handlingar som anges i artikel 1.1 a i detta direktiv.
Artikel 22
Artikel 23
Medlemsstaterna skall föreskriva att dessa personer inte får utföra en lagstadgad revision, om de inte är oberoende enligt lagstiftningen i den medlemsstat som kräver revisionen.
Artikel 26
Medlemsstaterna skall säkerställa att i varje fall de aktieägare och andra delägare i godkända revisionsbolag samt de ledamöter i dessa bolags förvaltnings-, lednings- och övervakningsorgan, som i en medlemsstat inte personligen uppfyller villkoren enligt artikel 3-19, inte ingriper i revisionsarbetet på något sätt som äventyrar oberoendet hos de fysiska personer som på revisonsbolagens vägnar reviderar de i artikel 1.1 angivna handlingarna.
1. Medlemsstaterna skall säkerställa att namn och adress för alla fysiska personer och revisionsbolag som av dem har godkänts att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna är offentligt tillgängliga.
c) Namn och adress för ledamöter i revisionsbolagets företagsledning.
Artikel 29
Artikel 30
3. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av följande: Genom artikel 5 i förordning nr 136/66/EEG införs en form av produktionsstöd för olivolja. Detta stöd för områden som är planterade med olivträd på ett visst datum beviljas odlare som är medlemmar av de producentorganisationer som anges i artikel 20c.1 i förordning nr 136/66/EGG och vars genomsnittliga produktion är minst 100 kg olja per regleringsår och till andra odlare på grundval av antalet olivträd samt produktionspotentialen och avkastningen från dessa träd, fastställd enligt en standardmetod, och under förutsättning att de odlade oliverna verkligen har skördats.
För att säkerställa att stödsystemet fungerar på rätt sätt bör rättigheterna och skyldigheterna för alla berörda parter, nämligen odlare, producentorganisationer och sammanslutningar av producentorganisationer samt de berörda medlemsstaterna, fastställas.
För att förvaltningen skall fungera på rätt sätt skall producentorganisationer och sammanslutningar av dessa hos de behöriga nationella myndigheterna ansöka om godkännande i god tid före regleringsårets början. Den behöriga medlemsstaten bör besluta om dessa ansökningar inom en skälig tid.
För att säkerställa att systemet med produktionsstöd till odlare som tillhör producentorganisationer fungerar på rätt sätt, bör bestämmelser införas om att stöd endast bör utbetalas för de kvantiteter som erhålls från godkända fabriker. För att bli godkända bör fabrikerna i fråga uppfylla flera villkor.
Erfarenheten har visat, att trots de många särskilda kontroller som införts är en noggrann och effektiv kontroll och verifiering svår att genomföra, på grund av det stora antalet odlare som skall kontrolleras. Dessa svårigheter måste lösas genom att ett dataregister upprättas i varje medlemsstat som innehåller all nödvändig information för att underlätta kontrollen och snabbt upptäcka oegentligheter.
Från och med regleringsåret 1984/1985 skall de allmänna bestämmelser som fastställs i denna förordning tillämpas vid beviljande av produktionsstöd för olivolja enligt artikel 5 i förordning nr 136/66/EEG.
För andra olivodlare skall stödet beviljas enligt artikel 5.2 andra strecksatsen i förordning nr 136/66/EEG, och stödet skall motsvara det stöd som erhålls om avkastningen från oliver och olivolja, fastställd enligt den standardmetod enligt artikel 18, tillämpas för antalet olivträd i produktion.
Artikel 3
- en kopia av den deklaration som lämnats för sammanställning av registret över olivodling. Denna deklaration får, när det gäller Grekland och till dess att registret över olivodling är sammanställt i den medlemsstaten, ersättas av den deklaration som anges i artikel 1.1 i förordning (EEG) nr 1590/83.
4. De olivodlare som avses i punkt 3 skall lämna skördedeklarationen och ansökan om stöd via sin organisation.
- en deklaration om att de har skördat sina oliver för regleringsåret i fråga, och
Artikel 4
b) i övriga fall, består av minst 1 200 olivodlare. Skulle en eller flera organisationer som producerar och ökar marknadsvärdet av oliver och olivolja vara medlemmar i organisationen i fråga, skall de berörda odlarna beaktas individuellt vid beräkning av det minsta antalet odlare som fordras, eller
För att uppnå detta skall olivodlare överlämna de upplysningar som behövs till de producentorganisationer som de tillhör för att fastställa att de brukar en olivodling samt uppgifter om alla förändringar som skett sedan de ansökte om medlemsskap.
Artikel 5
Tillståndet skall träda i kraft från början av det regleringsår som följer efter ansökningsåret.
Om villkoren inte längre uppfylls eller om organisationens struktur inte gör det möjligt att kontrollera medlemmarnas produktion, skall den behöriga myndigheten snarast och senast före det följande regleringsårets början återkalla godkännandet och anmäla sitt beslut om detta till kommissionen.
- lämna in skördedeklarationer från alla sina medlemmar enligt artikel 3.1,
Alla ansökningar som gäller produktionen från ett enda regleringsår skall, med risk för uteslutning, inlämnas före en fastställd dag.
Den kvantitet av olja för vilken stöd erhålls får inte vara större än den kvantitet som fastställs genom standardmetoden enligt artikel 18, dvs. att den fastställda skörden av oliver och olja tillämpas för antalet olivträd i produktionen, om en olivodlare som är medlem i en producentorganisation
- har blivit medlem i organisationen under regleringsåret.
- att den produktion av oliver, av varje odlare deklarerad som pressad i en godkänd fabrik, stämmer överens med de uppgifter som lämnats i hans skördedeklaration, på grundval av kännetecken som skall fastställas,
- Om de upplysningar som anges i punkt 1 första strecksatsen inte förefaller att stämma överens, efter det att organisationen har erhållit alla stöddokument och alla upplysningar som kan användas för att fastställa den kvantitet som verkligen producerats.
Artikel 9
2. Bestämmelserna om godkännande och återkallande av godkännande enligt vad som anges i artikel 5 skall även tillämpas för sammanslutningar. Artikel 10
- skall överlämna de skördedeklarationer och ansökningar om stöd som inlämnats till dem av de organisationer som de består av till de behöriga myndigheterna,
1. Det belopp som innehållits enligt artikel 20d.1 i förordning nr 136/66/EEG skall användas på följande sätt:
- antalet individuella ansökningar om stöd som inges till varje organisation av dess medlemmar,
3. Om beloppen inte används, helt eller delvis, såsom anges i punkt 2 skall de återbetalas till den behöriga medlemsstaten och avräknas från de utgifter som finansieras av EUGFJ.
Artikel 12
- det belopp som erhålls genom tillämpning av skörden av oliver och olja, fastställd enligt artikel 18, för antalet olivträd i produktion enligt skördedeklarationen eller det belopp som erhålls för den uppgivna kvantiteten i ansökan, om den kvantiteten är mindre än den som anges ovan, eller
1. Medlemsstaterna skall endast godkänna fabriker vars ägare
c) under det föregående regleringsåret inte blivit föremål för åtgärder beroende på oriktigheter som upptäckts vid kontroller enligt artikel 14 och denna artikel, beträffande godkännande för regleringsåret 1984/1985,
d) samtycka till att föra en standardiserad lagerredovisning enligt kriterier som skall fastställas.
Detta tillfälliga godkännande skall bli definitivt så snart den berörda medlemsstaten har förvissat sig om att de villkor för godkännande som fastställs i punkt 1 är uppfyllda.
5. I de fall godkännandet återkallas i enlighet med punkt 3 eller 4 får ingen ny ansökan om godkännande under den tid då godkännandet är återkallat beviljas.
Artikel 14
3. Under varje regleringsår och framför allt under den tid då oljan pressas, skall de producerande medlemsstaterna på plats kontrollera verksamheten och bokföringen hos en viss procent av de godkända fabrikerna, vilken skall fastställas.
- att skördedeklarationerna är riktiga,
5. Medlemsstaterna skall bl. a. använda de dataregister som föreskrivs i artikel 16 för dessa kontroller och verifieringar.
1. Medlemsstaterna skall besluta vilken kvantitet av olja är berättigad till stöd på grundval av de ansökningar som överlämnas enligt artiklarna 3 och 6, med hänsyn tagen till alla dithörande fakta och särskilt till alla kontroller och godkännanden som föreskrivs i denna förordning.
4. Som underlag för bestämmandet av den kvantitet som är berättigad till stöd, i de fall som omfattas av punkt 2 och 3, skall medlemsstaten framför allt använda skörden av oliver och olja, fastställd enligt den standardmetod som anges i artikel 18.
2. Dessa register skall innehålla minst följande information:
- de kvantiteter av producerad olja, för vilka en ansökan om produktionsstöd har inlämnats samt den kvantiteten för vilken stöd har utbetalats,
c) För fabriker som framställer olivolja och för varje regleringsår: de uppgifter som finns i lagerbokföringen, information om den tekniska utrustningen och pressningskapaciteten samt resultaten av de kontroller som utförts enligt denna förordning.
1. De register som anges i artikel 16 skall vara konfidentiella.
- Kommissionens tjänstemän i samarbete med de behöriga tjänstemännen i medlemsstaterna och enligt förordning (EEG) nr 729/70(), senast ändrad genom förordning (EEG) nr 3509/80(), särskilt med tanke på de fastställda förfarandena.
Artikel 18
Tillämpningsföreskrifter för denna förordning skall antas enligt förfarandet i artikel 38 i förordning nr 136/66/EEG.
- De belopp som anges i artikel 11.1 a.
Artikel 21
Medlemsstaterna skall anmäla de åtgärder som genomförs enligt denna förordning till kommissionen.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
Bestämmelserna i direktiv 64/433/EEG omfattar endast färskt kött som kan komma att föras i handel inom gemenskapen. Medlemsstaternas myndigheter har dock infört nationella kontroller av färskt kött som enbart är avsett för den nationella marknaden.
För att undanröja sådana skillnader bör harmoniserade regler fastställas för finansieringen av dessa hygienundersökningar och kontroller.
Artikel 1
P för att dels säkerställa lika behandling enligt artikel 15 i direktiv 71/118/EEG och dels täcka de omkostnader som avses i direktiv 72/462/EEG tar ut en avgift för det kött som avses i dessa direktiv och som importeras från tredje land,
2. Medlemsstaterna kan debitera en summa som överstiger den eller de belopp som avses i punkt 1, under förutsättning att den sammanlagda avgift som uttas i varje medlemsstat är lägre än eller lika med de faktiska kostnaderna för undersökningarna.
Artikel 4
Artikel 5
med beaktande av Europaparlamentets yttrande(),
Det förefaller ändå önskvärt att vissa bestämmelser införs för att underlätta det faktiska utövandet av etableringsrätten.
Inom ramen för ländernas hälso- och sjukvårdspolitik, som bl.a. går ut på att garantera en tillfredsställande utlämning av läkemedel överallt inom respektive lands territorium, begränsar vissa medlemsstater antalet nya apotek som får inrättas medan det i andra länder inte finns några bestämmelser av detta slag; under dessa omständigheter är det för tidigt att bestämma att följderna av ett erkännande av utbildnings-, examens- och andra behörighetsbevis i farmaci även skall omfatta utövandet av apotekarverksamhet som innehavare av ett apotek som varit öppet för allmänheten mindre än tre år; detta problem skall inom en viss bestämd tidsfrist utredas på nytt av kommissionen och rådet.
Detta direktiv påverkar inte medlemsstaternas lagar eller författningar med bestämmelser som förbjuder bolag att utöva vissa former av verksamhet eller ålägger dem vissa villkor för detta.
När det gäller verksamhet som anställd fastslås inte några särskilda bestämmelser i rådets förordning (EEG) nr 1612/68 av den 15 oktober 1968 om arbetskraftens fria rörlighet inom gemenskapen som hänför sig till god vandel eller gott anseende, yrkesansvar eller användningen av yrkestitlar(); beroende på den enskilda medlemsstaten tillämpas eller får dessa regler tillämpas på såväl anställda som självständigt verksamma yrkesutövare; sådan verksamhet för vilken det i alla medlemsstater krävs innehav av utbildnings-, examens- eller andra behörighetsbevis i farmaci utövas av såväl anställda som självständigt verksamma yrkesutövare eller av samma personer omväxlande som anställd eller som självständigt verksam yrkesutövare under deras yrkeskarriär; för att i möjligaste mån uppmuntra dessa yrkesutövares fria rörlighet inom gemenskapen förefaller det nödvändigt att utvidga detta direktiv till att även omfatta anställda.
Artikel 2
Fem år efter utgången av den tidsfrist som fastställts i artikel 19.1 skall kommissionen lägga fram en rapport för rådet om det sätt på vilket medlemsstaterna har tillämpat föregående stycke och om möjligheten att utvidga verkningarna av ett ömsesidigt erkännande av de utbildnings-, examens- och andra behörighetsbevis som avses i punkt 1. Den skall föreslå lämpliga åtgärder.
Så länge som Grekland använder denna undantagsbestämmelse och utan att det påverkar tillämpningen av artikel 45 i 1979 års anslutningsakt skall de övriga medlemsstaterna endast åläggas att tillämpa bestämmelserna i artikel 2 om de examensbevis som avses i artikel 4 d, såvida det gäller utövande av de former av verksamhet som avses i artikel 1 som anställd i enlighet med förordning (EEG) nr 1612/68.
De utbildnings-, examens- och andra behörighetsbevis som avses i artikel 2 är följande:
b) I Danmark:
1) Zeugnis über die staatliche Pharmazeutische Prüfung (statligt examensbevis för farmaceuter) som utfärdas av de behöriga myndigheterna,
Ðéáôïðïéçôéêü ôùí áñìïäßùí áñ÷þí, éêáíüôçôáò Üóêçóçò ôçò öáñìáêåõôéêÞò, ÷ïñçãïýìåíï ìåôÜ êñáôéêÞ åîÝôáóç (det intyg som visar att innehavaren av detta är behörig att utöva verksamhet som farmaceut) som utfärdas av de behöriga myndigheterna efter statsexamen;
f) I Irland:
Examensbevis eller intyg som innebär rätt att utöva verksamhet som farmaceut och som förvärvas efter statsexamen.
i) I Nederländerna:
Intyg som Registered Pharmaceutical Chemist.
Detta godkännande skall emellertid inte tillämpas på den tvååriga yrkeserfarenhet som krävs i Luxemburg för att tilldelas ett statligt tillstånd att driva ett apotek som är öppet för allmänheten.
och i båda fallen,
Artikel 7
Artikel 8
4. Medlemsstaterna skall garantera de lämnade upplysningarnas konfidentiella natur.
2. Om värdlandet har ingående kunskap om ett allvarligt sakförhållande som har uppstått utanför dess territorium, innan personen i fråga etablerade sig i det landet, och som sannolikt kommer att påverka rätten att inom dess territorium utöva verksamheten i fråga, får det landet underrätta ursprungslandet eller det senaste hemvistlandet om detta.
Om värdlandet kräver intyg om den fysiska och psykiska hälsan av de egna medborgare som vill påbörja eller utöva sådan verksamhet som avses i artikel 1, skall det landet som tillräckligt bevis godta den handling som krävs i ursprungslandet eller det senaste hemvistlandet.
Handlingar som utfärdats i enlighet med artikel 8, 9 och 10 får när de företes inte vara äldre än tre månader.
2. I de fall som avses i artikel 8.3 och 9.2 skall en begäran om utredning medföra att den tidsfrist som fastställts i punkt 1 förlängs.
Artikel 13
Om användningen av yrkestiteln för sådan verksamhet som avses i artikel 1 är reglerad i ett värdland, skall medborgare från andra medlemsstater som uppfyller villkoren i artikel 2, 5 och 6 använda den titel i värdlandet, som i det landet motsvarar denna utbildningsnivå, även i titelns förkortade form.
För detta ändamål får medlemsstaterna upprätta informationskontor där dessa personer kan få de upplysningar som behövs. Vid etablering får värdlandet kräva att personerna i fråga kontaktar dessa kontor.
Artikel 16
Inom den tidsfrist som fastställts i artikel 19.1 skall medlemsstaterna utse de myndigheter och organ som är behöriga att utfärda eller motta utbildnings-, examens- och andra behörighetsbevis samt de handlingar och upplysningar som avses i detta direktiv. De skall genast underrätta övriga medlemsstater och kommissionen om detta.
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta direktiv före den 1 oktober 1987. De skall genast underrätta kommissionen om detta.
Om det vid tillämpningen av detta direktiv skulle uppstå allvarligare svårigheter för en medlemsstat inom vissa områden, skall kommissionen i samverkan med det landet undersöka dessa svårigheter och begära yttrande från den farmaceutiska nämnd som upprättats enligt beslut 75/320/EEG().
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Europaparlamentets yttrande (2),
Med hänsyn till dessa målsättningar bör gemensamma grundregler införas om auktorisation, tillsyn, organisation och verksamheter för medlemsstaternas företag för kollektiva investeringar hemmahörande i medlemsstaterna och för den information de skall offentliggöra.
Den fria marknadsföringen av andelar som utgivits av fondföretag som fått tillstånd att placera upp till 100% av sina tillgångar i överlåtbara värdepapper från samma emittent (stat, lokal myndighet, etc.) får varken direkt eller indirekt åstadkomma störningar i kapitalmarknadens funktion eller medlemsstaternas finansiering eller skapa ekonomiska situationer av det slag som artikel 68.3 i fördraget avser att förhindra.
AVSNITT I Allmänna bestämmelser och räckvidd
4. Detta direktiv skall emellertid inte tillämpas på investeringsbolag vars tillgångar via dotterbolag är placerade huvudsakligen i annat än överlåtbara värdepapper.
7. Bestämmelserna i punkt 6 hindrar inte en medlemsstat att på fondföretag hemmahörande i den egna staten ställa krav som är strängare eller som går utöver vad som föreskrivs i artikel 4 och följande artiklar, förutsatt att kraven är generellt tillämpbara och inte står i strid med bestämmelserna i detta direktiv.
- Kategorier av fondföretag enligt vad som föreskrivs av medlemsstater där företagen hör hemma och för vilka bestämmelserna i avsnitt V och artikel 36 inte är ändamålsenliga med hänsyn till den placerings- och upplåningsinriktning som företagen har.
Vid tillämpningen av detta direktiv skall ett fondföretag anses hemmahörande i den medlemsstat där investeringsbolaget eller förvaltningsbolaget har sitt stadgeenliga säte; medlemsstaterna skall föreskriva att företagets huvudkontor skall vara beläget i samma medlemsstat som dess stadgeenliga säte.
1. Inget fondföretag får bedriva verksamhet utan auktorisation av behöriga myndigheter i den medlemsstat där företaget hör hemma (i fortsättningen kallade "behöriga myndigheter").
3. De behöriga myndigheterna får inte auktorisera ett fondföretag, om de som ingår i den verkställande ledningen för förvaltningsbolaget, investeringsbolaget eller förvaringsinstitutet inte har erforderlig vandel eller om de saknar tillräcklig erfarenhet för att kunna utföra sina uppgifter. För detta ändamål skall de behöriga myndigheterna utan dröjsmål underrättas om namnen på personer i sådan ledande ställning samt namnen på var och en som efterträder dem.
AVSNITT III Bestämmelser om värdepappersfonders organisation
Artikel 6
1. Tillgångarna i en värdepappersfond skall förvaras hos ett förvaringsinstitut.
e) tillse att en värdepappersfonds intäkter används i enlighet med lag eller annan författning och med fondbestämmelserna.
2. Ett förvaringsinstitut skall stå under offentlig tillsyn. Det skall också kunna ställa erforderliga ekonomiska garantier samt besitta tillfredsställande sakkunskap och kompetens för att kunna effektivt bedriva verksamhet som förvaringsinstitut och uppfylla därmed förenade åtaganden.
Ett förvaringsinstitut skall i enlighet med den nationella lagstiftningen i den stat där förvaltningsbolaget har sitt stadgeenliga säte vara ansvarigt mot förvaltningsbolaget och andelsägarna för förluster som drabbar dem som följd av att institutet allvarligt försummat sina förpliktelser eller fullgjort dem på ett oriktigt sätt. Detta ansvar kan av andelsägarna åberopas antingen direkt eller indirekt genom förvaltningsbolaget, beroende på hur rättsförhållandet mellan förvaringsinstitutet, förvaltningsbolaget och andelsägarna är utformat.
2. Förvaltningsbolaget och förvaringsinstitutet skall utföra sina respektive uppgifter självständigt och uteslutande i andelsägarnas intresse.
AVSNITT IV Bestämmelser om investeringsbolags organisation och och om deras förvaringsinstitut
Artikel 13
1. Ett investeringsbolags tillgångar skall förvaras hos ett förvaringsinstitut.
a) tillse att försäljning, utgivning, återköp, inlösen och makulering av andelar, som sker av eller på uppdrag av ett investeringsbolag, genomförs i enlighet med lag eller annan författning och med bolagsordningen,
Artiklarna 34, 37 och 38 skall inte gälla sådana bolag som nu sagts. Bestämmelserna om värdering av sådana bolags tillgångar måste emellertid vara angivna i lag eller annan författning eller i bolagsordningen.
b) agera (intervenera) på marknaden för att hindra att marknadsvärdet för andelarna avviker mer än 5% från nettovärdet,
6. Medlemsstaterna skall underrätta kommissionen om de investeringsbolag för vilka säregler, medgivna enligt punkterna 4 och 5, tillämpas.
1. Ett förvaringsinstitut skall antingen ha sitt stadgeenliga säte i samma medlemsstat som investeringsbolaget eller vara etablerat där om det har sitt stadgeenliga säte i en annan medlemsstat.
Artikel 16
1. Ett företag får inte samtidigt vara investeringsbolag och förvaringsinstitut.
Villkoren för utbyte av förvaringsinstitut skall, liksom regler till skydd för andelsägarna vid sådana utbyten, föreskrivas i lag eller annan författning eller anges i investeringsbolagets bolagsordning.
b) överlåtbara värdepapper som är föremål för handel på någon annan reglerad marknad i en medlemsstat och vilken marknadsplats fungerar fortlöpande och är erkänd och öppen för allmänheten, och/eller
b) en medlemsstat får föreskriva att ett fondföretag får placera högst 10% av sina tillgångar i fordringsbevis som med hänsyn till sin natur kan jämställas med överlåtbara värdepapper och för vilka bland annat gäller att de är överlåtbara och likvida och vars värde kan nöjaktigt bestämmas när som helst eller i vart fall så ofta som sägs i artikel 34,
3. Summan av placeringar som nämns i punkt 2 a och b får aldrig motsvara mer än 10% av ett fondföretags tillgångar.
b) närmare upplysningar om alla ändringar de avser att göra i förteckningar enligt a eller om andra instrument som de avser att jämställa med överlåtbara värdepapper, med angivande av skälen.
Artikel 22
3. Medlemsstaterna får höja den gräns som anges i punkt 1 till högst 35% om de överlåtbara värdepapperen är utgivna eller garanterade av en medlemsstat, av dess lokala myndigheter, av en icke-medlemsstat eller av offentliga internationella organ i vilka en eller flera medlemsstater är medlemmar.
De behöriga myndigheterna får medge sådana undantag endast om de finner att andelsägarna i fondföretaget har ett skydd likvärdigt med det som tillkommer andelsägarna i fondföretag som iakttar de gränsvärden som anges i artikel 22.
3. De fondföretag som avses i punkt 1 skall vidare i sina prospekt och reklambroschyrer på framträdande plats omnämna tillståndet och ange de stater, lokala myndigheter och/eller offentliga internationella organ i vars värdepapper de har för avsikt att placera eller har placerat mer än 35% av fondtillgångarna.
2. Ett fondföretag får placera högst 5% av sina tillgångar i andelar i sådana företag för kollektiva investeringar.
4. Punkt 3 skall även gälla i fall där ett investeringsbolag förvärvar fondandelar i ett annat investeringsbolag till vilket det är anknutet på det sätt som anges i punkt 3.
- 10% av de skuldebrev som en enskild emittent givit ut,
d) Ett fondföretags innehav av aktier i ett bolag beläget i en icke-medlemsstat och vars tillgångar placeras huvudsakligen i värdepapper utgivna av emittenter med sitt stadgeenliga säte i den staten, då den statens lagstiftning inte gör det möjligt för fondföretaget att på något annat sätt placera sina fondtillgångar i värdepapper med utgivare i staten. Detta undantag gäller dock endast om bolaget från icke-medlemsstaten vid sina placeringar följer de gränsvärden som anges i artiklarna 22, 24 och 25.1 och 25.2. Om gränsvärdena i artikel 22 och 24 har överskridits skall artikel 26 gälla i tillämpliga delar.
1. Fondföretag behöver inte iaktta de gränsvärden som anges i detta avsnitt när de utnyttjar teckningsrätter för överlåtbara värdepapper som ingår i fondtillgångarna.
Bestämmelser om information till andelsägarna A. Offentliggörande av prospekt och periodiska rapporter
- Två månader för halvårsrapporter.
2. Årsrapporten skall innehålla en balansräkning eller en redovisning av tillgångar och skulder, en specificerad resultaträkning för räkenskapsåret, en verksamhetsberättelse för räkenskapsåret samt den information som anges i lista B i bilagan till detta direktiv, liksom all annan väsentlig information som möjliggör för investerare att göra en välgrundad bedömning av utvecklingen av fondföretagets verksamhet och av dess resultat.
1. Fondbestämmelserna eller investeringsbolagets bolagsordning skall utgöra en del av prospektet och skall bifogas till detta.
All väsentlig information i ett prospekt måste hållas aktuell.
Artikel 32
1. Den som avser att teckna sig för förvärv av fondandelar skall innan avtalet ingås erbjudas att kostnadsfritt få prospektet, den senaste halvårsrapporten samt, i förekommande fall, den därpå följande halvårsrapporten.
B. Offentliggörande av annan information
Artikel 35
Artikel 36
- av fondens värde, i fråga om en värdepappersfond, förutsatt att upplåningen är av tillfällig art,
1. Ett fondföretag skall återköpa eller inlösa andelar när andelsägare begär det.
Artikel 38
Utdelningen eller återinvestering av en värdepappersfonds eller ett investeringsbolags intäkter skall ske i enlighet med lag eller annan författning och fondbestämmelserna eller investeringsbolagets bolagsordning.
Artikel 41
2. Bestämmelserna i punkt 1 skall inte hindra sådana företag från att förvärva överlåtbara värdepapper som inte är till fullo betalda.
I lag eller annan författning eller i fondbestämmelserna skall det anges vilken ersättning och vilka kostnader ett förvaltningsbolag har rätt att debitera en värdepappersfond och vilken metod som skall tillämpas för beräkning av sådana vederlag.
Artikel 44
3. Bestämmelserna i punkterna 1 och 2 får inte tillämpas på ett diskriminerande sätt.
Artikel 46
- där det anses lämpligt, sin senaste årsrapport och eventuell senare halvårsrapport, samt - upplysningar om de åtgärder som vidtagits för försäljning av dess andelar i den andra medlemsstaten.
Ett fondföretag skall i sin verksamhet ha rätt att använda samma företagsbeteckning (t.ex. investeringsbolag eller värdepappersfond) inom hela gemenskapen som det använder i den medlemsstat där det är hemmahörande. Om det finns risk för förväxling kan värdmedlemsstaten i förtydligande syfte begära att namnet skall åtföljas av något förklarande tillägg.
1. Medlemsstaterna skall utse de myndigheter som skall fullgöra de uppgifter som föreskrivs i detta direktiv. Medlemsstaterna skall underrätta kommissionen om detta och i förekommande fall ange hur uppgifterna fördelats mellan myndigheterna.
4. De berörda myndigheterna skall ges alla de befogenheter som de behöver för att utföra sina uppgifter.
2. Medlemsstaterna skall föreskriva att alla som är eller har varit anställda hos de myndigheter som avses i artikel 49 skall vara bundna av tystnadsplikt. Detta innebär att ingen konfidentiell information som erhållits i tjänsten får röjas för någon person eller myndighet annat än med stöd av bestämmelser i lag eller annan författning.
Artikel 51
Artikel 52
3. Myndigheterna i den medlemsstat där ett fondföretag är beläget skall utan dröjsmål underrätta myndigheterna i de medlemsstater där företaget utbjuder sina andelar om beslut som avser återkallelse av auktorisation, andra allvarliga åtgärder som riktar sig mot företaget samt uppskov med återköp eller inlösen.
1. En kontaktkommitté, i fortsättningen kallad kommittén, skall inrättas vid sidan av kommissionen. Dess funktion skall vara
c) att, om så erfordras, föreslå kommissionen tillägg till eller ändringar i detta direktiv.
4. Kommittén skall sammankallas av dess ordförande antingen på dennes eget initiativ eller på begäran av en medlemsstats delegation. Kommittén skall självständigt fastställa sin arbetsordning.
Uteslutande med avseende på danska fondföretag skall "pantebreve" utställda i Danmark jämställas med de överlåtbara värdepapper som avses i artikel 19.1 b.
Artikel 56
Artikel 57
3. Grekland och Portugal tillåts att uppskjuta genomförandet av detta direktiv till senast den 1 april 1992.
Artikel 58
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Europaparlamentets yttrande (2),
Ett sådant samarbete kan möta svårigheter av rättslig, skattemässig eller psykologisk natur. Ett ändamålsenligt rättsligt instrument på gemenskapsnivå i form av en europeisk ekonomisk intressegruppering skulle bidra till att ovannämnda mål uppnås och behövs därför.
En gruppering skiljer sig från ett bolag främst i fråga om ändamålet, vilket endast är att underlätta eller utveckla medlemmarnas ekonomiska verksamhet för att göra det möjligt för dessa att förbättra sina egna resultat. På grund av denna stödjande karaktär måste grupperingens verksamhet ha samband med medlemmarnas ekonomiska verksamhet och får inte ersätta denna i sådan utsträckning att grupperingen t.ex. i förhållande till tredje man utövar en självständig yrkesmässig verksamhet, varvid begreppet ekonomisk verksamhet skall ges en vidsträckt tolkning.
Förordningens bestämmelser om möjlighet att av hänsyn till allmänna intressen förbjuda eller begränsa rätten att delta i en gruppering inverkar inte på de rättsregler i medlemsstaterna som behandlar utövande av verksamhet och som kan föreskriva ytterligare förbud eller begränsningar eller annan kontroll eller tillsyn i fråga om rätten för fysiska personer, bolag eller andra rättsliga enheter eller kategorier därav att delta i en gruppering.
Frågor om fysiska personers rättsliga handlingsförmåga och rättskapacitet samt om juridiska personers rättskapacitet regleras av nationell lagstiftning.
Denna förordning föreskriver att det endast är grupperingens medlemmar som skall beskattas för resultatet av grupperingens verksamhet. Därutöver tillämpas nationella skatteregler, bl.a. när det gäller fördelningen av vinst, taxeringsförfarandet och alla förpliktelser som medlemsstaternas skattelagstiftning innehåller.
- konkurrensrätt,
Det står medlemsstaterna fritt att tillämpa eller anta lagar eller förordningar eller vidta administrativa åtgärder som inte strider mot tillämpningsområdet för eller syftet med denna förordning.
De som avser att bilda en gruppering skall ingå ett avtal och låta registrera grupperingen enligt artikel 6.
a) direkt eller indirekt utöva någon form av styrning eller kontroll över medlemmarnas egen verksamhet eller över något annat företags verksamhet, särskilt inte i personal-, finansierings- eller investeringsfrågor,
d) utnyttjas av ett bolag för att lämna lån till ledningen i ett bolag eller till någon ledningen närstående person, om rätten att bevilja sådana lån är begränsad eller underkastad kontroll enligt medlemsstaternas bolagsrätt; en gruppering får inte heller utnyttjas för att föra över egendom mellan ett bolag och dess ledning eller någon ledningen närstående person utöver vad som är tillåtet enligt medlemsstaternas bolagsrätt; i denna bestämmelse avses med att lämna lån även att medverka i transaktioner med motsvarande verkan, och med egendom avses lös och fast egendom,
1. Endast följande kan vara medlemmar i en gruppering:
2. En gruppering skall omfatta minst
c) ett bolag eller någon annan rättslig enhet som avses i punkt 1 och en fysisk person, av vilka den förstnämnda har sitt huvudkontor i en medlemsstat och den senare utövar sin huvudsakliga verksamhet i någon annan medlemsstat.
Artikel 5
b) Grupperingens säte.
e) Tiden för grupperingens bestånd, om inte denna tid är obestämd.
Artikel 7
b) Uppgift om inrättande eller nedläggning av ett huvudkontor eller avdelningskontor för grupperingen.
e) Uppgift om när en medlem enligt artikel 22.1 har överlåtit sin andel eller en del av denna.
h) Uppgift om att likvidationen av en gruppering har avslutats enligt artikel 35.2.
Artikel 8
b) Registreringsnummer, datum och ort för registreringen samt uppgift om att denna har upphört.
Artikel 9
Artikel 10
Efter offentliggörandet i den i artikel 39.1 avsedda tidningen skall i Europeiska gemenskapernas officiella tidning föras in uppgifter om bildandet av en gruppering och om avslutandet av en grupperings likvidation med uppgift om grupperingens registreringsnummer, datum och plats för registreringen, datum och plats för offentliggörandet samt den förstnämnda tidningens namn.
Sätet skall vara beläget
Artikel 13
Artikel 14
2. En gruppering får avföras ur det tidigare registret först sedan det visats att grupperingen har tagits in i det nya registret.
Artikel 15
3. Ett avgörande varigenom ogiltigheten av en gruppering fastställs eller tillkännages kan göras gällande mot tredje man enligt artikel 9.1.
1. Medlemmarna gemensamt och en eller flera företagsledare utgör grupperingens organ.
Artikel 17
a) ändra föremålet för grupperingens verksamhet,
d) förlänga grupperingens varaktighet utöver den tid som har bestämts i avtalet om att bilda grupperingen,
g) vidta andra ändringar i avtalet om att bilda grupperingen än som anges i denna punkt, om inte annat är bestämt i avtalet.
Artikel 19
- enligt den lagstiftning som gäller för honom, eller
inte får tillhöra styrelsen eller direktionen i ett bolag, inte får leda ett företag eller inte får vara företagsledare i en europeisk ekonomisk intressegruppering.
Förbuden enligt punkt 1 gäller också för representanterna.
1. Endast företagsledaren eller, om de är flera, var och en av dem företräder grupperingen mot tredje man.
2. I avtalet om att bilda grupperingen kan bestämmas att endast två eller flera företagsledare i förening får företräda denna. En sådan bestämmelse kan göras gällande mot tredje man enligt artikel 9.1 endast om den har offentliggjorts enligt artikel 8.
2. Grupperingens medlemmar skall bidra till att betala belopp varmed utgifterna överstiger inkomsterna enligt vad som är bestämt i avtalet om att bilda grupperingen eller, om sådana bestämmelser saknas, med lika delar.
2. En medlem kan endast med de övriga medlemmarnas enhälliga medgivande använda sin andel i grupperingen som säkerhet, om inte något annat är bestämt i avtalet om att bilda grupperingen. Innehavaren av en sådan säkerhet kan inte bli medlem på grund av säkerheten.
1. Medlemmarna svarar obegränsat solidariskt för alla grupperingens förbindelser. Följderna av detta ansvar bestäms av den nationella lagstiftningen.
På brev, beställningssedlar och liknande handlingar skall följande tydligt anges:
c) Adressen för grupperingens säte.
Varje enligt artikel 10 registrerat kontor skall på de nu nämnda handlingarna som härrör från kontoret lämna de angivna uppgifterna och motsvarande uppgifter som gäller kontorets egen registrering.
2. Varje ny medlem svarar enligt artikel 24 för grupperingens förbindelser, inräknat sådana som har uppkommit i verksamheten före medlemmens inträde.
2. En medlem kan uteslutas på de grunder som anges i avtalet om att bilda grupperingen och under alla förhållanden, om medlemmen väsentligt åsidosätter sina skyldigheter eller vållar eller hotar att vålla allvarliga störningar i grupperingens verksamhet.
1. Ett medlemskap upphör när medlemmen dör eller inte längre uppfyller de i artikel 4.1 angivna villkoren.
Artikel 29
Utom då avtalet att bilda grupperingen föreskriver något annat och med förbehåll för den rätt som någon kan ha förvärvat enligt artiklarna 22.1 och 28.2, skall grupperingen efter det att ett medlemskap har upphört fortsätta att bestå med de kvarvarande medlemmarna och på de villkor som är bestämda i avtalet om att bilda grupperingen eller som de sistnämnda medlemmarna enhälligt beslutar.
a) tiden för grupperingens bestånd enligt avtalet om att bilda denna har löpt ut eller någon annan i avtalet angiven grund för upplösning föreligger, eller
3. En gruppering skall även upplösas genom ett beslut av medlemmarna eller den kvarvarande medlemmen om de i artikel 4.2 angivna villkoren inte längre är uppfyllda.
1. På ansökan av den som saken angår eller en behörig myndighet skall rätten förordna att en gruppering skall upplösas om bestämmelserna i artikel 3, 12 eller 31.3 har åsidosatts, såvida inte rättelse vidtas innan rätten har avgjort ärendet.
Artikel 33
Artikel 34
1. Avvecklingen av en gruppering skall ske genom likvidation.
4. Likvidatorerna skall vidta de åtgärder som avses i artiklarna 7 och 8.
Artikel 37
Artikel 38
Medlemsstaterna skall vidare se till att var och en har möjlighet att vid det register som avses i artikel 6 respektive 10 ta del av de i artikel 7 angivna handlingarna och att, även med post, få fullständiga eller partiella kopior av dessa handlingar.
3. Medlemsstaterna skall bestämma lämpliga påföljder för underlåtenhet att iaktta föreskrifterna om offentliggörande i artiklarna 7, 8 och 10 och föreskrifterna i artikel 25.
Artikel 41
Artikel 42
b) vid behov ge kommissionen råd om tillägg till eller ändringar i förordningen.
med beaktande av rådets förordning (EEG) nr 1035/72/EEG(1) av den 18 maj 1972 om den gemensamma organisationen av marknaden för frukt och grönsaker, senast ändrad genom förordning (EEG) nr 1332/84(2),
De blanketter som avses i rådets förordning (EEG) nr 850/80(5) bör därför anpassas till de nya bestämmelserna.
Enda artikel
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: I artikel 2 i förordning (EEG) nr 3117/85 fastställs vissa villkor för beviljande av ekonomisk kompensation för produkterna, att den kvantitativa begränsningen skall vara 2 000 ton, vilka mottagarna av stödet skall vara samt metoden för beräkning av detta.
De former av beredning som är tillåtna bör preciseras i syfte att klart ange omfattningen av den aktuella ordningen.
Enligt artikel 2.3 i anslutningsfördraget får gemenskapens institutioner före anslutningen vidta de åtgärder som anges i artiklarna 171 och 358 i akten.
- fångats av medlemmarna,
a) frysning,
Artikel 3
Om någon av de beredningsprocesser som anges i artikel 2.2 utförs i en annan medlemsstat än den som erkänt den producentorganisation som säljer produkten, skall bevis om att sådan beredning ägt rum företes i form av kontrollformulär T nr 5 i enlighet med bestämmelserna i kommissionens förordning (EEG) nr 223/77() och i denna förordning.
- I fält 104 en av följande angivelser med versaler:
2. Beredaren skall skriftligt åta sig att bereda de produkter som ingår i avtalet i enlighet med bestämmelserna i artikel 2. Han måste därför i sin lagerförteckning kunna identifiera de kvantiteter som inköpts i samband därmed. Beredaren skall förplikta sig att upplåta sina lokaler för varje form av inspektion av de behöriga myndigheterna.
1. De berörda medlemsstaterna skall införa ett kontrollsystem för att säkerställa att de produkter för vilka ansökan om bidrag lämnats in berättigar till sådant och att bestämmelserna i denna förordning följts.
- Mottagaren av bidraget skall lämna in de handlingar på vilka han grundar sina anspråk på rätt till bidraget.
Artikel 7
3. På grundval av den information som framkommit vid kontrollen enligt artikel 6 skall i förekommande fall bidragets storlek korrigeras.
Artikel 9
med beaktande av följande: I kommissionens förordning (EEG) nr 3143/85 av den 11 november 1985 om försäljning till sänkt pris av interventionssmör för användning till direkt konsumtion i form av koncentrerat smör(3), senast ändrad genom förordning (EEG) nr 3338/85(4), föreskrivs att förpackningar med koncentrerat smör skall vara försedda med vissa påskrifter som är skrivna med klart synliga och läsliga tryckbokstäver. På grund av ett fel motsvarar påskriften på italienska språket inte den påskrift som antagits i den text som förelagts Förvaltningskommittén för mjölk och mjölkprodukter för röstning. Följaktligen bör nämnda förordning rättas.
I artikel 5.4 första stycket skall den näst sista strecksatsen ersättas med följande:
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Europaparlamentets yttrande (),
Rådets resolution av den 10 april 1984 om gemenskapspolitik på turistområdet () understryker behovet av samråd mellan medlemsstaterna och kommissionen i fråga om turism.
I avsikt att ha samråd inom turistområdet bör informationsutbyte säkerställas mellan medlemsstaterna och kommissionen.
Artikel 1
Kommitténs uppgift skall vara att underlätta informationsutbyte, samråd och, när så är lämpligt, samarbete om turism och då i synnerhet tjänster för turister.
Kommissionen skall underrätta de andra medlemsstaterna om detta.
4. Den information och det samråd som föreskrivs i detta beslut skall omfattas av tystnadsplikt.
Kommissionen skall tillhandahålla sekreterartjänster åt kommittén.
I enlighet med artikel 2.3 i Fördraget om Spaniens och Portugals anslutning får gemenskapens institutioner besluta om de åtgärder som åsyftas i artikel 396 i anslutningsakten, vilka åtgärder skall träda i kraft om och när fördraget träder i kraft.
Med verkan från den 1 januari 1986 skall artikel 11 k i direktiv 85/384/EEG kompletteras med följande:
Syftet med sådana minimikrav på kvalitet är att förhindra framställning av produkter som inte efterfrågas eller produkter som skulle leda till en snedvridning av marknaden. Kraven måste baseras på traditionella och sunda framställningsmetoder.
Förvaltningskommittén för bearbetade produkter av frukt och grönsaker har inte lämnat något yttrande inom den tidsfrist som dess ordförande har bestämt.
Denna förordning fastställer de minimikvalitetskrav som produkter som framställs av tomater enligt definitionen i artikel 1.2 i förordning (EEG) nr 1599/84 skall uppfylla för att få del av det produktionsstöd som avses i artikel 2.1 i förordning (EEG) nr 426/86.
I denna avdelning betyder "skalade tomater"
1. Skalade tomater får endast tillsättas
P tomatkoncentrat,
Som tillsatsämnen vid framställning av skalade tomater får endast citronsyra (E 330) och kalciumklorid (509) användas.
Artikel 5
3. Mögeltalet för skalade tomater (tomaterna och den omgivande vätskan) skall inte överstiga 50 % positiva fält och pH-värdet får inte överstiga 4,5.
P skador: 35 cm2 sammantagen yta,
P tomater i bitar: 1 250 cm2 sammantagen yta.
a) skador: områden där skador på ytan har trängt igenom och som därigenom skiljer sig starkt i färg eller konsistens från den normala tomatvävnaden och som normalt borde ha avlägsnats under bearbetningen,
1. Vad avser skalade konserverade tomater skall tomaterna och den omgivande vätskan uppta minst 90 % av behållarens volym.
Artikel 8
1. Tomatsaft och tomatkoncentrat får endast tillsättas följande:
2. Som tillsatsämne vid framställning av tomatsaft och tomatkoncentrat får citronsyra (E 330) användas. Vidare, vid framställning av
3. Kvantiteten tillsatt vanligt salt får inte överstiga
Vid bestämning av kvantiteten tillsatt vanligt salt skall det naturliga innehållet av klorider anses vara lika med 2 % av torrsubstansinnehållet.
a) en karakteristisk röd färg, och
a) fria från synligt främmande beståndsdelar av vegetabiliskt ursprung, däribland skal, frön och andra hårda delar av tomater,
a) eventuella främmande beståndsdelar av vegetabiliskt ursprung endast kan urskiljas genom en noggrann undersökning med blotta ögat, och
a) en jämnt fördelad konsistens och beskaffenhet som visar att en korrekt bearbetningsmetod har använts,
d) en flyktig surhet, uttryckt som ättiksyra på högst 0,4 viktprocent av torrsubstansen, minskat med eventuell tillsats av vanligt salt,
Artikel 11
1. Tomatflingor skall
c) vara fria från främmande smaker och lukter.
4. Som tillsatsämne vid framställning av tomatflingor får endast kiseldioxid (551) användas. Kiseldioxidinnehållet får dock inte överstiga 1 viktprocent.
2. Bestämmelserna i punkt 1 skall även gälla andra tomatbaserade produkter om sådana produkter vid bearbetningstillfället förpackas i behållare i vilka de skall lämna bearbetningsanläggningen. Om de förvaras i tankar eller liknande behållare ämnade för senare förpackning eller vidare bearbetning, skall datumet eller datumen för framställningen anges på behållarna. När sådana produkter förpackas i de slutliga behållarna skall det på dessa finnas en referens som gör det möjligt att fastställa datumet eller datumen för framställningen samt bearbetningsföretaget.
Bearbetningsföretaget skall dagligen och med jämna mellanrum under bearbetningen kontrollera att produkterna uppfyller kraven för beviljande av stöd. Resultatet av kontrollen skall registreras. Artikel 15
b) naturliga lösliga substanser,
e) den totala surheten,
h) pH-värde,
Artikel 16
med beaktande av följande: Artikel 30 och följande i fördraget, om avskaffande av kvantitativa restriktioner och alla åtgärder med motsvarande verkan, gäller utan åtskillnad för de varor som har sitt ursprung i gemenskapen och sådana som har övergått till fri omsättning i någon av medlemsstaterna oberoende av ursprung.
En fullständig tillämpning av dessa principer förutsätter emellertid en fungerande gemensam handelspolitik.
För detta ändamål har kommissionen befogenhet att til låta medlemsstater att, utan hinder av principen om fri rörlighet inom gemenskapen, besluta om övervakningsåtgärder eller skyddsåtgärder inom gemenskapen gentemot varor som har sitt ursprung i tredje land och som övergått till fri omsättning i någon av medlemsstaterna. I artikel 115 föreskrivs emellertid att sådana åtgärder enbart kan tillåtas om de är nödvändiga och att kommissionen skall ge företräde åt åtgärder som vållar de minsta störningarna när det gäller den gemensamma marknadens funktion. Följden är att på det nuvarande stadiet av genomförandet av den gemensamma marknaden åtgärder enligt artikel 115 i fördraget bör tillåtas endast i fall där en störning i handeln leder till ekonomiska svårigheter eller äventyrar effektiviteten av handelspolitiska åtgärder som medlemsstater har vidtagit i överensstämmelse med gemenskapens internationella åtaganden.
I de fall då en övervakningsåtgärd tillåts måste en importhandling utfärdas automatiskt och utan avgift, inom en given frist och för varje begärd mängd. Om övervakningsåtgärder begärs på grund av att import kan leda till ekonomiska svårigheter för en medlemsstat, bör en sådan risk bedömas mot bakgrund av de störningar i handeln som dittills iakttagits och av storleken av de importmöjligheter gemenskapen har beviljat tredje land i fråga.
Om så är nödvändigt bör kommissionen få företa en undersökning för att kontrollera giltigheten av de uppgifter som den har fått till sitt förfogande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Detta beslut gäller för import till en medlemsstat av varor med ursprung i tredje land, som har övergått till fri omsättning inom gemenskapen och inte är underkastade enhetliga importvillkor i medlemsstaterna.
1. När det kan befaras att import till en medlemsstat av en sådan vara som avses i artikel 1 kan leda till ekonomiska svårigheter, får som villkor för import med tidsbegränsat tillstånd från kommissionen, krävas att en importhandling utfärdas.
b) importmöjligheter som gemenskapen har öppnat för varan gentemot det tredje land som är ursprungsland inte överstiger 1 % av de sammanlagda importmöjligheterna som gemenskapen har öppnat gentemot alla tredje länder för vilka liknande regler gäller.
a) En beskrivning av varan med närmare uppgifter om dess handelsbeteckning, dess nummer i Gemensamma tulltaxan, dess NIMEXE-nummer och dess ursprungsland.
- i tredje landet i fråga, med fördelning på direkt import och varor i fri omsättning,
d) Risken för ekonomiska svårigheter som åberopas och huruvida de framgår av sådana faktorer som förbrukningen av varan och de marknadsandelar som gäller för inhemsk produktion, för tredje landet i fråga och för alla tredje länder.
a) Uppgifter som identifierar importören samt avsändaren i den exporterande medlemsstaten.
- dess handelsbeteckning,
e) Planerad dag eller planerade dagar för leverans.
Skyddsåtgärder
3. För att få tillstånd skall medlemsstaten i sin ansökan till kommissionen lämna följande uppgifter utöver de uppgifter som avses i artikel 2.4 a och 2.4 b:
c) Den faktiska eller tillåtna importvolymen eller importmängden för varan i fråga
- med ursprung i alla tredje länder,
e) De åberopade ekonomiska svårigheterna, vilka framgår av sådana faktorer som produktion, kapacitetsutnyttjande, förbrukning, försäljning, marknadsandelarna för det tredje landet i fråga, för alla tredje länder och för inhemsk produktion, samt priser (dvs. pressade priser eller uteblivna normala prisstegringar), vinster eller förluster, sysselsättning.
5. I de fall då medlemsstaten finner att den volym eller den sammanlagda mängd som omfattas av ansökningar under prövning avseende import av varan i fråga med ursprung i tredje landet överstiger antingen 5 % av eventuell direkt import från det tredje landet eller 1 % av den sammanlagda importen från länder utanför EEG under den senaste tolvmånadsperiod för vilken statistiska uppgifter finns tillgängliga, skall dock följande gälla:
6. Medlemsstaten skall sända in sin ansökan om tillstånd till skyddsåtgärder med telex eller telefax. En kopia skall samtidigt och på samma sätt sändas till de behöriga myndigheter som för detta syfte har utsetts av de andra medlemsstaterna. Medlemsstaten skall vidare underrätta dem som har ansökt om importhandlingar om att en ansökan om skyddsåtgärder har lämnats in.
Ursprungsbevis
Slutbestämmelser De förfaranden som fastställs genom detta beslut skall gälla när verkan av de handelspolitiska åtgärder som en medlemsstat tillämpar i överensstämmelse med gemenskapens internationella åtaganden äventyras av en störning i handeln med undantag för vad som avses i artiklarna 2.4 d och 3.3 e.
2. Kommissionens beslut 80/47/EEG skall upphöra att gälla från och med samma dag. Hänvisningar till det upphävda beslutet skall betraktas som hänvisningar till detta beslut.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(2), och
För att förfarandet för typgodkännande skall kunna tillämpas fullständigt är det nödvändigt att det omfattar såväl komponenter som särskilda tekniska enheter och att varje begrepp definieras noggrant.
Ett förtydligande behövs för de administrativa förfaranden som styr förhållandet mellan medlemsstaterna, i det fall en medlemsstat påvisar att ett antal fordon inte överensstämmer med den godkända typen för den medlemsstat som har utfärdat typgodkännandet och att det därför finns skäl att anta att produktionens överensstämmelse inte har kontrollerats i tillräcklig grad.
Artikel 1
- fordon: dels varje motordrivet fordon avsett att användas på väg, med eller utan karosseri, som har minst fyra hjul och som är konstruerad för en högsta hastighet som överstiger 25 km/tim, dels släpvagnar till dessa fordon, spårbundna fordon, jordbrukstraktorer och lantbruksmaskiner är undantagna,
Artikel 2
-"agrément par type"/"typegoedkeuring" i belgisk lagstiftning,
- "Ýãêñéóç ôýðïõ" i grekisk lagstiftning,
- "type approval" i irländsk lagstiftning,
- "typegoedkeuring" i nederländsk lagstiftning,
b) EEG-typgodkännande avser det förfarande genom vilket en medlemsstat fastställer att en fordonstyp, en särskild teknisk enhet eller komponent, uppfyller de tekniska kraven i särdirektiven och de kontroller som anges i EEG-typgodkännandeintyget. En förebild för detta visas i bilaga 2 och skall, i tillämpliga fall, kompletteras enligt bilagan till typgodkännandeintyget i det berörda direktivet."
1. Varje medlemsstat skall godkänna alla fordonstyper som uppfyller följande villkor:
2. En medlemsstat som har beviljat ett typgodkännande skall vidta nödvändiga åtgärder för att, i nödvändig utsträckning och vid behov i samarbete med behöriga myndigheter i andra medlemsstater, kontrollera att tillräckliga åtgärder har gjorts som säkerställer att serietillverkade fordon överensstämmer med den godkända typen.
Artikel 5
3. Tillverkaren eller dennes representant i registreringslandet skall för varje fordon som tillverkas i enlighet med den godkända typen utfärda ett intyg om överensstämmelse, för vilket en förebild visas i bilaga 3.
Ett fordon anses inte överensstämma med den godkända typen om det avviker från uppgifterna i typgodkännandeintyget och/eller det tekniska underlaget förutsatt att dessa avvikelser inte har godkänts under artikel 6.2 eller 6.3 av den medlemsstat som har beviljat typgodkännandet. Ett fordon skall inte anses avvika från den godkända typen om toleranser som anges i särdirektiv inte överskrids."
1. Om en medlemsstat som har utfärdat EEG-typgodkännandet finner att ett antal fordon med intyg om överensstämmelse inte överensstämmer med den godkända typen, skall den vidta nödvändiga åtgärder för att säkerställa att serietillverkade exemplar överensstämmer med den godkända typen. De behöriga myndigheterna i denna stat skall upplysa motsvarande myndigheter i de andra medlemsstaterna om vidtagna åtgärder vilket, om så är påkallat, kan leda till att EEG-typgodkännandet återkallas. 2. Om en medlemsstat påvisar att ett antal fordon med intyg om överensstämmelse inte överensstämmer med den godkända typen kan denna stat begära att medlemsstaten som har utfärdat EEG-typgodkännandet visar att serietillverkade fordon överensstämmer med den godkända typen. Medlemsstaten som utfärdade EEG-typgodkännandet skall, inom sex månader räknat från dagen för en begäran, kontrollera att produktionen är i överensstämmelse med den godkända typen. Kontrollen kan, om så bedöms nödvändigt, utföras i samarbete med den medlemsstat som begärde att en sådan kontroll skulle utföras.
4. Om medlemsstaten som beviljade EEG-typgodkännandet ifrågasätter den påpekade avvikelsen, skall de berörda medlemsstaterna bemöda sig att bilägga tvisten.
"Artikel 9a
3. Emellertid skall innehavaren av EEG-typgodkännande för en särskild teknisk enhet eller en komponent, vilka beviljats i enlighet med denna artikel, utfärda intyget som beskrivs i artikel 5.3 och märka varje enhet eller komponent som tillverkats i enlighet med den godkända typen med handelsbeteckning eller varumärke, typen och, om så anges i särdirektivet, typgodkännandets nummer. I det senare fallet medför detta ingen skyldighet att utfärda intyget som föreskrivs i artikel 5.3.
"- vid ansökan från en tillverkare eller dennes representant och inlämnandet av de upplysningar som krävs enligt särdirektivet, skall den berörda medlemsstaten färdigställa intyget om typgodkännande i enlighet med det tillgängliga särdirektivet. En kopia av intyget skall sändas till sökanden. Andra medlemsstater skall, för fordon av samma typ, acceptera denna kopia som bevis på att nödvändiga provningar har utförts."
Artikel 3
Artikel 4
med beaktande av följande: Vetenskapliga och tekniska framsteg medför att vissa ändringar måste göras i bilagan till direktiv 79/117/EEG.
De åtgärder som föreskrivs genom detta direktiv är förenliga med yttrandet från Ständiga kommittén för växtskydd.
2. I del B, "Svårnedbrytbara organiska klorföreningar", under 1, "Aldrin", skall texten till b i andra kolumnen ändras genom att orden "Irland och" utgår.
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(1), senast ändrad genom förordning nr (EEG) 1454/86(2), särskilt artikel 5.4 i denna,
Innan medlemsstaterna har möjlighet att definitivt godkänna en fabrik skall de utföra vissa kontroller. För att göra det möjligt för fabrikerna att börja sin verksamhet bör bestämmelser införas för beviljande av ett tillfälligt tillstånd under en begränsad tid, så snart som ansökan har lämnats in.
Första stycket i artikel 13.3 i förordning (EEG) nr 2261/84 skall ersättas med följande:
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 113 i detta,
med beaktande av följande: Enligt beslut 83/539/EEG(3) har gemenskapen provisoriskt tillämpat Internationella kaffeavtalet 1983 sedan denna provisoriskt trädde i kraft den 1 oktober 1983.
För att säkerställa en effektiv förvaltning av systemet och för att klargöra frågan under vilken tid denna förordning faktiskt kommer att gälla, och för att uppfylla regel 11 i bilagan till denna förordning och till regel 47 i bilagan till förordning (EEG) nr 3761/83, bör åtgärder vidtas för kommissionen, enligt de beslut som fattats av de behöriga organen i Internationella kaffeorganisationen och vid den tid då kvoterna är tillfälligt upphävda eller återinförs, för att ange den dag då åtgärderna i fråga skall bli tillämpliga eller upphöra att vara tillämpliga.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
I artikel 6.3 i kommissionens förordning (EEG) nr 3440/84() fastställs att det är tillåtet att sätta fast en förstärkande nätkasse på trålar, danska snurrevadar och liknande nätredskap under förutsättning att dess maskstorlek är minst 80 millimeter.
Definitionerna på nätkategorierna i artiklarna 5 och 6 i förordning (EEG) nr 3440/84 behöver därför ändras.
Artikel 1
"5. Det är förbjudet att använda ett övre slitskydd tillsammans med förstärkande nätkassar, med undantag för trålar med en maskstorlek på 60 mm eller mindre."
"2. Det är bara tillåtet att använda en förstärkande nätkasse åt gången, med undantag för trålar med en maskstorlek på högst 60 mm, för vilka två förstärkande nätkassar får användas."
- Punkt 6 skall ersättas med följande:
"7. Trots punkt 1 får en förstärkande nätkasse som är mindre än lyftet sättas fast på redskap med en maskstorlek på högst 60 mm."
KOMMISSIONENS FÖRORDNING (EEG) nr 4155/87 av den 22 december 1987 om ändring av vissa förordningar om tillämpningen av den gemensamma organisationen av marknaden för ägg till följd av införandet av Kombinerade nomenklaturen
Artikel 1 i kommissionens förordning nr 54/65/EEG () av den 7 april 1965 om icke-fastställande av en tilläggsavgift för polska ägg skall ersättas med följande: "Artikel 1 I enlighet med artikel 8.2 i förordning (EEG) nr 2771/75 skall de importavgifter som skall betalas vid import av fjäderfäägg med skal (undernummer 0407 00 i Kombinerade nomenklaturen) som har sitt ursprung i och kommer från Polen, inte höjas med en tilläggsavgift."
Artikel 3
Artikel 1 i kommissionens förordning nr 765/67/EEG av den 26 oktober 1967 om icke-fastställande av en tilläggsavgift för australiska ägg () skall ersättas med följande: "Artikel 1 Importavgifter som fastställts i enlighet med artikel 3 i förordning (EEG) nr 2771/75 skall inte höjas med en tilläggsavgift när det gäller import av färska, konserverade, kokta eller på annat sätt värmebehandlade fjäderfäägg med skal, undantaget kläckägg som omfattas av undernummer 0407 00 30 i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Australien."
2. Artikel 2 skall ersättas med följande: "Artikel 2 Importförändringar som fastställts i enlighet med artikel 2 i förordning (EEG) nr 2783/75 avseende produkter som omfattas av följande undernummer i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Österrike, skall inte höjas med en tilläggsavgift: () EGT nr L 186, 1.7.1974, s. 14. () EGT nr 260, 27.10.1967, s. 24. () EGT nr L 130, 31.5.1969, s. 4. >Plats för tabell>
Artikel 7
Denna förordning träder i kraft den 1 januari 1988.
med beaktande av rådets förordning (EEG) nr 1898/87 av den 2 juli 1987 om skydd för beteckningar som används vid saluförande av mjölk och mjölkprodukter(1), senast ändrad genom förordning (EEG) nr 222/88(2), särskilt artikel 4.2 b i denna, och
Artikel 2 Detta beslut riktar sig till medlemsstaterna.
För fordon i kategori N2 med en massa över 7,5 ton och andra fordon än dragfordon för påhängsvagn i kategori N3 har nuvarande krav visat sig otillräckliga vad avser det yttre siktfältet längs fordonets sida och bakåt. För att råda bot på denna brist är det nödvändigt att möjliggöra montering av en extra backspegel av s.k. vidvinkeltyp.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
- eller förbjuda att fordon tas i bruk,
- Medlemsstaterna får inte längre utfärda dokumentet enligt artikel 10.1 tredje strecksatsen i direktiv 70/156/EEG för en typ av fordon, vars backspeglar inte överensstämmer med bestämmelserna i det här direktivet.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Europaparlamentets yttrande(),
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 11.2 skall ersättas med följande:
"Artikel 22
"Kapitel IIa
Sändningar som innehåller varuprov av referenssubstanser som godkänts av Världshälsoorganisationen för kvalitetskontroll av material som används vid tillverkning av läkemedel och som är adresserade till mottagare som är bemyndigade av medlemsstaternas behöriga myndigheter att ta emot sådana försändelser utan att erlägga skatt skall vara skattebefriade vid införsel."
6. Artiklarna 62 och 63 skall ersättas med följande:
a) varor som är till salu eller uthyrning av en person som är etablerad utanför införselmedlemsstaten, eller
Artikel 63
b) Varje försändelse får innehålla högst ett dokument eller ett enda exemplar av varje dokument om det består av flera dokument. Försändelser innefattande flera exemplar av samma dokument får emellertid beviljas befrielse, om deras sammanlagda bruttovikt inte överstiger ett kilogram.
7. Följande tillfogas till artikel 79:
"Bränslen och smörjmedel som finns i motorfordon och specialcontainrar"
b) bränsle som finns i reservdunkar som fraktas av privata motorfordon och motorcyklar, dock högst 10 liter per fordon, med förbehåll för nationella bestämmelser om innehav och transport av bränsle.
- varor,
- tankar som av tillverkaren är fast monterade i alla containrar av samma typ som containern i fråga och vars fasta installation gör det möjligt att använda bränslet direkt för att under transporten driva kylsystem och övriga system som specialcontainrar är utrustade med.
- I inledningen införs orden "och specialcontainrar" efter orden "kommersiella motorfordon".
12. Följande tillfogas till artikel 91:
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta direktiv senast den 1 januari 1989. De skall genast underrätta kommissionen om detta.
med beaktande av rådets förordning (EEG) nr 3878/87 av den 18 december 1987 om produktionsstöd för vissa rissorter(1), senast ändrad genom förordning (EEG) nr 1424/88(2), särskilt artikel 2.3 i denna, och med beaktande av följande:
De analysmetoder som skall användas när dessa morfologiska och kvalitativa kännetecknen fastställs, bör närmare anges.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- En klibbighet på högst 2,50 gcm.
1. De medlemsstater som vill få en rissort som berättigar till stöd införd i bilaga B till förordning (EEG) nr 3878/87, skall senast den 31 juli varje år till kommissionen överlämna en ansökan där sortens namn anges samt dess inskrivningsreferenser i den nationella sortlistan över jordbruksgrödor.
2. Varje prov som sänds in till laboratorierna för analys skall bestå av minst 100 g råris och minst 750 g helt slipat ris. Proven skall endast bestå av hela riskorn, dock skall hela men kritaktiga korn avlägsnas från prov av helt slipat ris.
2. Om en och samma sort är föremål för två eller flera ansökningar, skall dess kännetecken bestämmas som medelvärdet av provresultaten enligt punkt 1.
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Förordning (EEG) nr 2658/87 fastställer de allmänna bestämmelserna för tolkningen av Kombinerade nomenklaturen och dessa bestämmelser gäller också varje annan nomenklatur som helt eller delvis grundar sig på denna eller som lägger ytterligare underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser med tanke på tillämpningen av tulltaxebestämmelser eller andra bestämmelser som rör varuhandeln.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
med beaktande av kommissionens förslag(1),
Med hänsyn till den viktiga roll som dessa organ kan spela för att säkerställa att avtalen om produktionsstöd tillämpas på ett korrekt och enhetligt sätt, bör en metod föreskrivas för finansiering av deras faktiska utgifter som gör det möjligt för dem att ha en smidig och effektiv verksamhet inom ramen för en självständig administration som föreskrivs i dessa bestämmelser. Det syftet kan uppnås genom en metod som förenar gemenskapsfinansiering med finansiering av medlemsstaten.
Artikel 1
- För Italien 100 % för de första tre åren upp till högst 14 miljoner ecu och 50 % för det fjärde och femte året,
För Spanien och Portugal skall 100 % av organets faktiska utgifter under tiden från den 1 mars 1986 till den 31 oktober 1990 täckas av de europeiska gemenskapernas allmänna budget upp till högst 9 300 000 ecu för Spanien och 4 700 000 ecu för Portugal. Under tiden från den 1:a november 1990 till den 31 oktober 1992 skall 50 % av de ifrågavarande utgifterna täckas av denna budget.
Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
i samarbete med Europaparlamentet(2),
Direktiv enligt artikel 118a i fördraget får inte medföra sådana administrativa, ekonomiska och rättsliga hinder, som skulle kunna hämma bildandet och utvecklingen av små och medelstora företag.
Europaparlamentet antog i februari 1988 fyra resolutioner i anslutning till debatten om den inre marknaden och arbetarskydd; i dessa resolutioner anmodas kommissionen uttryckligen att utarbeta ett ramdirektiv, som skall ligga till grund för särdirektiv, vilka skall omfatta alla risker förknippade med säkerhet och hälsa på arbetsplatsen.
Antalet arbetsolycksfall och arbetssjukdomar är alltjämt för högt; förebyggande åtgärder måste införas eller förbättras utan dröjsmål för att trygga arbetstagarnas säkerhet och hälsa och säkra en högre skyddsnivå.
Förbättring av arbetarskyddet för arbetstagarna är ett mål som inte skall underordnas rent ekonomiska hänsyn.
En kommitté bestående av ledamöter nominerade av medlemsstaterna behöver tillsättas för att bistå kommissionen med de tekniska bearbetningarna för de särdirektiv, som föreskrivs i detta direktiv.
3. Detta direktiv skall inte hindra tillämpningen av sådana gällande eller framtida bestämmelser i medlemsstaterna och i gemenskapen som är gynnsammare vad gäller skyddet för arbetstagarnas säkerhet och hälsa.
1. Detta direktiv skall tillämpas på all verksamhet, såväl privat som offentlig ( industri, jordbruk, handel, förvaltning, tjänster, undervisning, kultur- och fritidsverksamhet etc.).
Artikel 3
a) arbetstagare, varje person anställd av en arbetsgivare, inklusive praktikanter och lärlingar men inte arbetstagare i arbetsgivarens hushåll,
d) förebyggande, alla mått och steg som vidtas eller planeras i något skede av verksamheten för att förebygga eller minska risker i arbetet.
2. Medlemsstaterna skall i synnerhet se till att en ändamålsenlig kontroll och tillsyn säkerställs.
Allmänna bestämmelser
3. Arbetstagarnas skyldigheter på arbetarskyddsområdet skall inte inverka på arbetsgivarens ansvar.
1. Inom ramen för sina skyldigheter skall arbetsgivaren vidta tillräckliga åtgärder till skydd för arbetstagarnas säkerhet och hälsa, inbegripet förebyggande av risker i arbetet och tillhandahållande av information och utbildning samt iordningställande av erforderlig organisation och nödvändiga resurser.
3. Utan att det inskränker de övriga bestämmelserna i detta direktiv skall arbetsgivaren göra följande med beaktande av verksamhetens art:
- garantera en förbättring av skyddsnivån för arbetstagarna med avseende på säkerhet och hälsa,
c) Arbetsgivaren skall se till att planläggning och införande av ny teknik blir föremål för överläggningar med arbetstagarna och/eller deras representanter i fråga om följdverkningarna för arbetstagarnas säkerhet och hälsa i samband med val av utrustning och förändringar i arbetsbetingelser och arbetsmiljön.
5. Åtgärder som rör säkerhet, hygien och hälsa i arbetet får under inga förhållanden medföra några kostnader för arbetstagarna.
1. Utan att det inskränker skyldigheterna enligt artiklarna 5 och 6 skall arbetsgivaren ge en eller flera arbetstagare i uppgift att verka för skydd mot och förebyggande av risker i arbetet inom företaget och/eller verksamheten.
4. I de fall då arbetsgivaren anlitar sakkunnig hjälp utifrån skall han informera de personer som anlitas om de faktorer som påverkar eller misstänks påverka arbetstagarnas säkerhet och hälsa och personerna skall ha tillgång till sådan information som avses i artikel 10.2.
- utifrån anlitade företag eller personer ha tillräckliga kunskaper och tillräckliga personella och professionella resurser, och
7. Med hänsyn tagen till verksamheternas art och företagens storlek skall medlemsstaterna ange de verksamhetsgrenar, där arbetsgivaren, under förutsättning att han har kompetens, själv kan ta ansvaret för de åtgärder som avses i punkt 1.
Artikel 8
- upprätta alla behövliga kontakter med utomstående serviceorgan, framför allt i fråga om första hjälpen, akutvård, räddningsarbete och brandbekämpning.
3. Arbetsgivaren skall
c) utom i sådana undantagsfall då det finns väl underbyggda skäl för det, avhålla sig från att anmoda arbetstagarna att återgå till arbetet i ett läge, där en allvarlig och överhängande fara fortfarande föreligger.
Arbetstagarnas åtgärder får inte leda till att de på något sätt missgynnas, såvida de inte handlat vårdslöst eller visat grov försumlighet.
1. Arbetsgivaren skall
c) föra ett register över arbetsolycksfall, som resulterat i att arbetstagaren varit arbetsoförmögen under mer än tre dagar,
Artikel 10
a) arbetsmiljörisker och skydds- och förebyggande åtgärder och verksamhet med avseende såväl på företaget och/eller verksamheten i stort som varje enskild arbetsplats och/eller varje enskilt arbete,
3. Arbetsgivaren skall vidta lämpliga åtgärder, så att arbetstagare med särskilda uppgifter i skyddsfrågor eller arbetstagarrepresentanter med särskilt ansvar för skyddsfrågor, för de skall kunna utföra sina uppgifter och i enlighet med nationell lagstiftning och praxis, får tillgång till
c) den kunskap som skydds- och förebyggande åtgärder, tillsynsmyndigheter och arbetsmiljöansvariga organ avkastar.
1. Arbetsgivarna skall inhämta synpunkter från arbetstagarna och/eller deras representanter och låta dem delta i diskussioner om alla frågor som gäller säkerhet och hälsa på arbetsplatsen.
- rätt för arbetstagarna och/eller deras representanter att lägga fram förslag,
a) varje åtgärd som på ett väsentligt sätt kan påverka arbetsmiljön,
d) i förekommande fall, anlitande av tjänster eller personer utifrån enligt artikel 7.3,
4. De arbetstagare, som avses i punkt 2, och de arbetstagarrepresentanter, som avses i punkterna 2 och 3, får inte missgynnas på något sätt på grund av sin verksamhet enligt punkterna 2 och 3.
Artikel 12
- anställning,
- införande av ny teknik.
- vid behov upprepas regelbundet.
4. Den utbildning som avses i punkterna 1 och 3 får inte bekostas av arbetstagarna eller arbetstagarrepresentanterna.
AVSNITT III ARBETSTAGARNAS SKYLDIGHETER
Artikel 14
2. De åtgärder som avses i punkt 1 skall vara av sådan karaktär att varje arbetstagare, som så önskar, kan genomgå regelbundna hälsokontroller.
Riskgrupper
1. Efter förslag från kommissionen med stöd av artikel 118a i fördraget skall rådet anta särdirektiv, bland annat på de områden som uppräknas i bilagan.
Artikel 17
- antagandet av direktiv om teknisk harmonisering och standardisering, och/eller
2. Kommissionens företrädare skall till kommittén lämna ett förslag till åtgärder som skall vidtas.
Vid omröstningen i kommittén skall de röster som avges av representanterna för medlemsstaterna vägas enligt artikeln i fördraget. Ordföranden får inte delta i omröstningen.
Om rådet inte fattar beslut inom tre månader från det att förslaget har mottagits, skall kommissionen besluta att de föreslagna åtgärderna skall vidtas.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de redan har antagit eller som de antar på det område som omfattas av detta direktiv.
4. Kommissionen skall regelbundet överlämna en rapport till Europaparlamentet, rådet och Ekonomiska och sociala kommittén om tillämpningen av detta direktiv med beaktande av punkterna 1, 2 och 3.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(),
I avvaktan på att skattegränserna upphävs såsom behövs för att uppnå en verklig inre marknad, är det nödvändigt att harmonisera och lätta på vissa formaliteter som krävs för beviljandet av den införselbefrielse som föreskrivs i direktiv 83/183/EEG, särskilt vad beträffar upprättandet av en förteckning över egendomen och bevisning om den normala hemvisten. Det är nödvändigt att lätta på gällande regler om användningstiden för importerad egendom och de kvantitativa begränsningarna för vissa artiklar.
Direktiv 83/183/EEG ändras på följande sätt:
För de varor som avses i punkt a andra meningen får medlemsstaterna kräva att den flyttande skall ha haft dem i bruk före flyttningen minst
4. I artikel 7 görs följande ändringar:
5. I artikel 8.2 görs följande ändringar:
6. I artikel 9 görs följande ändringar:
b) Punkt 2 skall ersättas med följande:
a) I punkt 1 skall orden "Fram till ikraftträdandet av de gemenskapsskatteregler som införs i överensstämmelse med artikel 14.2 i direktiv 77/388/EEG skall medlemsstaterna" utgå och punkten inleds därefter med "Medlemsstaterna skall".
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
På det veterinära området utnyttjas för närvarande gränserna för att utföra kontroller som syftar till att värna om hälsan hos människor och djur.
Denna lösning förutsätter ett ökat förtroende för de veterinära kontroller som utförs av den avsändande staten. Den senare måste säkerställa att dessa veterinära kontroller utförs på ett lämpligt sätt.
Ett förfarande bör fastställas för att bilägga eventuella tvister i fråga om sändningar från någon anläggning, något produktionsställe eller något företag.
Dock föreligger alltjämt med avseende på vissa epizootiska sjukdomar olika hälsosituationer inom medlemsstaterna och i avvaktan på ett ställningstagande från gemenskapens sida vad gäller sätten att bekämpa dessa sjukdomar bör frågan om kontroll av handeln med husdjur inom gemenskapen tills vidare lämnas utanför och en kontroll av handlingar bör vara tillåten under transporten. Med hänsyn till det rådandet läget vad gäller frågan om harmonisering och i avvaktan på gemenskapsregler bör varor som inte är underkastade harmoniserade regler uppfylla de krav som gäller inom destinationslandet, förutsatt att de senare står i överensstämmelse med artikel 36 i fördraget.
Kommissionen bör bemyndigas att vidta åtgärder för tillämpningen av detta direktiv. I detta syfte bör det utarbetas rutiner för att upprätta ett nära och effektivt samarbete mellan kommissionen och medlemsstaterna inom Ständiga veterinärkommittén.
Medlemsstaterna skall se till att de veterinära kontroller som skall utföras på produkter av animaliskt ursprung, som omfattas av de direktiv som räknas upp i bilaga A eller i artikel 14 och som är avsedda för handel, inte längre sker vid gränserna utan verkställs i enlighet med detta direktiv, utan att det påverkar tillämpningen av artikel 6.
1. veterinär kontroll: varje fysisk undersökning eller administrativt förfarande som gäller de varor som avses i artikel 1 och som syftar till att direkt eller på annat sätt värna om människors eller djurs hälsa,
4. behörig myndighet: den centrala myndighet i en medlemsstat som det åligger att utföra veterinära kontroller eller varje myndighet till vilken denna uppgift har överförts,
1. Medlemsstaterna skall se till att inga andra produkter görs till föremål för handel än sådana som avses i artikel 1 och som har anskaffats, kontrollerats, stämplats och märkts i enlighet med gemenskapens regler för den angivna destinationen och som fram till den slutlige mottagare som uppgivits åtföljs av ett hälsointyg, djurhälsocertifikat eller något annat dokument som fastställts genom gemenskapens veterinära bestämmelser.
När det finns anledning att misstänka att kraven inte uppfylls skall den behöriga myndigheten utföra nödvändiga kontroller och, i de fall misstanken bekräftas, vidta lämpliga åtgärder, vilket kan innefatta indragning av godkännandet.
3. Medlemsstater som valt att föra in produkter från vissa länder utanför gemenskapen skall meddela kommissionen och övriga medlemsstater om förekomsten av sådan import.
Artikel 4
- de produkter som omfattas av bilaga B inte förs ut till någon annan medlemsstats territorium, om de inte kan försäljas inom medlemsstatens eget territorium av skäl som har stöd i artikel 36 i fördraget.
a) Den behöriga myndigheten får på destinationsorten för varorna genom icke-diskriminerande veterinära stickprov kontrollera att de krav som uppställs i artikel 3 har uppfyllts. Provtagning får ske samtidigt.
- för en anläggning som står under tillsyn av en officiell veterinär, skall denne se till att endast sådana produkter släpps in i denna anläggning som uppfyller kraven i artikel 3.1 med avseende på märkning och medföljande dokument eller, vad gäller de produkter som avses i bilaga B, åtföljs av de dokument som fastställs i destinationslandets bestämmelser,
De garantier som skall företes av de mottagare som avses i andra och tredje strecksatserna skall specificeras i ett avtal med den behöriga myndigheten att undertecknas vid tiden för den registrering som föreskrivits i punkt 3. Den behöriga myndigheten skall utföra stickprovskontroller för att förvissa sig om att dessa garantier uppfylls.
a) de dessförinnan skall bli föremål för registrering, om den behöriga myndigheten kräver detta,
d) de skall under den tid som fastställts av den behöriga myndigheten, dock under minst sex månader, arkivera de hälsointyg och dokument som avses i artikel 3 för att vid anfordran företes för den behöriga myndigheten.
Artikel 6
b) Vid införsel av produkter från länder utanför gemenskapen, skall de sändas under tullövervakning till inspektionsställen där veterinär besiktning kan utföras.
- antingen underkastas veterinär besiktning som visar att de uppfyller de bestämmelser som utfärdats i den medlemsstat till vilken de destinerats, eller
2. Dock skall från den 1 januari 1993 och utan hinder av punkt 1 alla produkter som transporteras genom reguljära och direkta transportmedel som förbinder två geografiska punkter inom gemenskapen vara underkastade de bestämmelser om inspektion som fastställs i artikel 5.
a) förekomst av smittämnen som orsakar någon av de sjukdomar som nämns i direktiv 82/894/EEG(4), senast ändrat genom kommissionens beslut 89/162/EEG(5), någon zoonos eller sjukdom eller något annat som kan tänkas orsaka allvarlig fara för djur och människor eller om produkterna kommer från ett område som är smittat med en epizootisk sjukdom, skall de utom vad gäller djurhälsoaspekter, i fråga om produkter som är föremål för någon av de behandlingar som avses i artikel 4 i direktiv 80/215/EEG(6), senast ändrat genom direktiv 88/660/EEG(7), beordra att transportförpackningen i fråga förstörs eller används på något annat sätt som fastställts genom gemenskapsregler.
De skyddsåtgärder som anges i artikel 9 får tillämpas.
- förstöra varorna eller
2. I enlighet med det förfarande som fastställs i artikel 18 skall kommissionen upprätta en förteckning över de smittämnen och sjukdomar som avses i punkt 1 och fastställa detaljerade regler för hur denna artikel skall tillämpas.
Om myndigheten i den första medlemsstaten befarar att dessa åtgärder är otillräckliga, skall de behöriga myndigheterna i de två medlemsstaterna gemensamt söka finna en lösning. Om det är lämpligt kan detta innefatta inspektion på platsen.
- sända en inspektionsgrupp till den berörda anläggningen, eller
Den skall underrätta medlemsstaterna om vad som framkommit.
Den mottagande medlemsstaten får å sin sida utöka kontrollerna av produkter som kommer från samma anläggning.
2. Rätten enligt medlemsstatens gällande lagstiftning att begära prövning av beslut som fattats av de behöriga myndigheterna skall inte påverkas av detta direktiv.
Om tvist skulle uppkomma, och utan att det påverkar tillämpningen av den nyssnämnda rätten till prövning, får dock de två berörda parterna, om överenskommelse träffas om detta inom en period av högst två månader, hänskjuta tvisten för avgörande till någon expert vars namn finns med på en av kommissionen upprättad förteckning över gemenskapens experter. Kostnaden för att anlita denna expert skall betalas av gemenskapen.
Artikel 9
I avvaktan på att åtgärder vidtas i enlighet med punkt 4 får den mottagande medlemsstaten, när särskilt allvarliga folk- eller djurhälsoskäl föreligger, vidta tillfälliga skyddsåtgärder gentemot de berörda anläggningarna eller, i fråga om en epizootisk sjukdom, vad gäller det skyddsområde som fastställs i gemenskapens regler.
3. Om kommissionen inte har informerats om vilka åtgärder som vidtagits, eller om den anser de vidtagna åtgärderna otillräckliga, får den, i samarbete med den berörda medlemsstaten och i avvaktan på att den Ständiga veterinärkommittén sammanträder, vidta tillfälliga skyddsåtgärder gentemot produkter från den region som berörs av den epizootiska sjukdomen eller produkter från en viss anläggning. Dessa åtgärder skall underställas Ständiga veterinärkommittén snarast möjligt för att fastställas, ändras eller upphävas i enlighet med förfarandet i artikel 17.
Artikel 10
Medlemsstaterna skall se till att tjänstemännen inom deras veterinärmyndigheter, om så är lämpligt i samarbete med tjänstemännen inom andra myndigheter som anförtrotts denna uppgift särskilt ges fullmakt och möjlighet att
- ta prover på produkter som finns i lager för att förvaras, släppas ut på marknaden eller transporteras,
Artikel 12
3. I direktiv 74/461/EEG(11), senast ändrat genom direktiv 87/489/EEG(12),
4. Artikel 7.3 och artiklarna 12 och 16 i direktiv 77/99/EEG(13), senast ändrat genom direktiv 89/227/EEG(14), utgår.
ii) i artikel 7a skall hänvisningarna till artikel 7 ersättas med en hänvisning till artikel 9 i direktiv 89/662/EEG.
8. Artiklarna 8 och 9 i direktiv 89/437/EEG(17) utgår.
1. Följande artikel skall läggas till direktiven 64/433/EEG och 71/118/EEG:
"Artikel 15
4. Följande artikel skall läggas till direktiven 85/397/EEG och 88/657/EEG:
"Artikel 17
Medlemsstaterna skall före det datum som fastställs i artikel 19 meddela vilka villkor och förfaranden som för närvarande tillämpas vid handeln med de produkter som avses i första stycket.
I artikel 9 i direktiv 64/432/EEG(19)skall följande punkt införas:
1. Medlemsstaterna skall senast tre månader före det datum som fastställs i artikel 19.1 tillställa kommissionen ett program som redovisar de nationella åtgärder som kommer att vidtas för att förverkliga de angivna målen med detta direktiv, särskilt hur ofta kontrollerna kommer att utföras.
Artikel 17
Rådet skall fatta sitt beslut med kvalificerad majoritet.
1. När det förfarande som fastställs i denna artikel skall tillämpas, skall ordföranden utan dröjsmål hänskjuta ärendet till den ständiga veterinärmedicinska kommittén (i det följande kallad "kommittén") som inrättats genom beslut 68/361/EEG.
4. Om förslaget inte är förenligt med yttrandet från kommittén eller om inget yttrande avgives, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas.
1. Före den 31 december 1990 skall rådet fatta sitt beslut med kvalificerad majoritet om kommissionens förslag rörande veterinärkontroller vid handel mellan medlemsstaterna med levande djur.
Artikel 20
- verkställa kontroller av handlingar under transporten av produkter som importerats från tredje land och som är avsedda för medlemsstaterna.
Artikel 22
Artikel 23
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
i samarbete med Europaparlamentet (2),
Gällande bestämmelser för tillämpning av direktiven på såväl nationell som gemenskapsnivå är inte alltid tillräckliga för att garantera efterlevnad av i sammanhanget relevanta gemenskapsregler, i synnerhet inte i ett skede, då överträdelser kan korrigeras.
Det är nödvändigt att se till att lämpliga förfaranden finns inom alla medlemsstater, så att beslut i strid mot dess bestämmelser kan upphävas och ersättning kan ges till dem som skadats av överträdelserna.
Tillämpningen av detta direktiv bör utvärderas inom en period av fyra år från genomförandet på grundval av information från medlemsstaterna om prövningsförfarandets funktion i respektive länder.
1. Medlemsstaterna skall vidta nödvändiga åtgärder för att garantera, att en upphandlande myndighets beslut prövas effektivt, vad beträffar upphandling inom ramen för direktiv 71/305/EEG och 77/62/EEG. I synnerhet skall prövningar göras skyndsamt enligt reglerna i följande artiklar, där särskilt uppmärksammas artikel 2.7 för de fall upphandlingsbeslut innefattar överträdelse av gemenskapsrätten för offentlig upphandling eller nationella bestämmelser om införande av sådan lag.
Artikel 2
b) antingen åsidosätta eller garantera åsidosättande av olagliga beslut, vilket innefattar undanröjandet av diskriminerande tekniska, ekonomiska eller finansiella specifikationer i anbuds- eller kontraktshandlingarna eller i varje annat dokument som har samband med upphandlingen,
3. Prövningsförfarandet i sig behöver inte automatiskt bidra till att upphandlingen skjuts upp.
Medlemsstaterna får dessutom bestämma att, utom i fall där ett beslut måste undanröjas innan ersättning ges ut, prövningsorganets behörighet sedan ett upphandlingsavtal genomförts skall begränsas till att lämna ersättning till den som lidit skada av överträdelsen.
Medlemmarna i ett sådant oberoende organ skall tillsättas och frånträda på samma villkor som gäller för rättsliga instanser, tillämpade av den myndighet som utnämner och avsätter dem, samt bestämmer ämbetsperiodens längd. Åtminstone ordföranden i prövningsorganet skall ha domarkompetens. Det oberoende organet skall fatta sina beslut i ett förfarande, där båda parter hörs, och besluten skall vara lagligen bindande enligt regler bestämda av medlemsstaten.
2. Kommissionen skall underrätta den berörda medlemsstaten och den upphandlande myndigheten om de skäl, som föranlett bedömningen att en klar och konkret överträdelse föreligger och kräva rättelse.
b) förklaring till varför rättelse ej skett, eller
5. Då uppgift har lämnats om att en upphandling har avbrutits enligt punkt 3 c, skall medlemsstaten underrätta kommissionen om när upphandlingsförfarandet återupptas, eller när någon annan upphandlingsprocedur med hel eller delvis anknytning till upphandlingen påbörjats. Underrättelsen skall bekräfta, att den påstådda överträdelsen har rättats eller om så inte är fallet, skälen till varför rättelse inte har skett.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
Förordning (EEG) nr 2658/87 fastställer de allmänna bestämmelserna för tolkningen av Kombinerade nomenklaturen och dessa bestämmelser gäller också varje annan nomenklatur som helt eller delvis grundar sig på denna eller som lägger ytterligare underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser med tanke på tillämpningen av tulltaxebestämmelser eller andra bestämmelser som rör varuhandeln.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
med beaktande av följande: För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen som är en bilaga till förordning (EEG) nr 2658/87 vad avser tulltaxeklassificering av anoraker, skidjackor, vindjackor och liknande artiklar som omfattas av bl.a. KN-nummer 6101, 6102, 6201 och 6202, är det nödvändigt att ange vissa kännetecknande egenskaper för dessa klädesplagg.
Nomenklaturkommittén har inte avgivit något yttrande inom den tid som dess ordförande bestämt.
Endast klädesplagg med långa ärmar skall klassificeras som anoraker, skidjackor, vindjackor och liknande artiklar enligt KN-nummer 6101, 6102, 6201 och 6202.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(2),
För somliga rubriker hade dock inga gränsvärden fastställts i avvaktan på beslut av rådet efter ytterligare utredning, främst av vetenskapliga experter.
Vissa andra uppgifter i denna bilaga bör också anpassas till de senaste vetenskapliga rönen inom detta område.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Tillämpningsföreskrifter till denna förordning, en lista över mindre viktiga livsmedel tillsammans med de gränsvärden som skall tillämpas på dessa, samt gränsvärden för djurfoder, skall antas enligt artikel 30 i förordning (EEG) 804/68, som skall tillämpas på motsvarande sätt. För detta ändamål skall en kommitté tillsättas."
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
I brev av den 26 september 1989 har myndigheterna i Spanien till kommissionen framfört en begäran om undantag från punkt 45 c i bilaga 1 till direktiv 64/433/EEG i fråga om styckning av färskt nötkött, fårkött och griskött. I begäran föreslås hygienkrav. Det är nödvändigt att de alternativa hygienkrav som fastställs i det begärda undantaget i fråga om styckning av färskt kött lägst motsvarar kraven i punkt 45 c i bilaga 1 till direktiv 64/433/EEG.
med beaktande av rådets direktiv 64/433/EEG av den 26 juni 1964 om hygienproblem som påverkar handeln med färskt kött inom gemenskapen(1), senast ändrat genom direktiv 88/657/EEG(2), särskilt artikel 13 i detta, och
De hygienkrav som föreslås a
med beaktande av rådets förordning (EEG) nr 2658/87(1) om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan, senast ändrad genom förordning (EEG) nr 3945/89(2), särskilt artikel 9 i denna, och med beaktande av följande:
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt de tillämpliga KN-nummer som anges i kolumn 2, av de skäl som anges i kolumn 3.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Enligt bestämmelserna i direktiv 77/93/EEG får växter av vissa släkten, med undantag för frukter och fröer, med ursprung i andra länder eller regioner än dem som har erkänts vara fria från Erwinia amylovora (Burr.) Winsl. et al. inte föras in till vissa medlemsstater från och med den 16 april till och med den 31 oktober om växterna har sitt ursprung på norra halvklotet samt från och med den 1 november till och med den 15 april om de har sitt ursprung på södra halvklotet.
Detta beslut inverkar inte på senare upptäckter som kan visa att den ovan nämnda organismen förekommer i landet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE. Artikel 1
RÅDETS DIREKTIV av den 21 mars 1991 om ändring för nionde gången i direktiv 76/769/EEG om tillnärmning av medlemsstaternas lagar och andra författningar om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar) (91/173/EEG)
med beaktande av kommissionens förslag(1),
med beaktande av följande: Åtgärder bör vidtas för att stegvis upprätta den inre marknaden under tiden fram till den 31 december 1992. Den inre marknaden skall vara ett område utan inre gränser, inom vilket den fria rörligheten för varor, personer, tjänster och kapital är säkerställd.
Kommissionen kommer att utarbeta en samordnad gemenskapskapsstrategi som avser rätten att släppa ut på marknaden och använda kemiska produkter för träskyddsändamål. Denna strategi utarbetas på grundval av uppgifter som medlemsstaterna lämnar, särskilt om hälso- och miljörisker, och med beaktande av de svårigheter som finns i medlemsstaterna på detta område.
med beaktande av kommissionens förslag (),
Artikel 2
1. Båtförarcertifikat som fortfarande är giltiga och som är upptagna i grupp A i bilaga 1 skall erkännas av alla medlemsstater som giltiga för navigering på de vattenvägar av havskaraktär som är upptagna i bilaga 2, som om de själva hade utfärdat ifrågavarande båtförarcertifikat.
4. En medlemsstats erkännande av ett båtförarcertifikat får begränsas till de kategorier av fartyg för vilka detta certifikat gäller i den medlemsstat som har utfärdat det.
Om så behövs skall kommissionen vidta nödvändiga åtgärder för att anpassa förteckningen över certifikat i bilaga 1 i enlighet med det förfarande som anges i artikel 7.
Artikel 6
2. Kommissionens företrädare skall förelägga kommittén ett förslag till ändring av bilaga 1. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen varvid medlemsstaternas röster skall vägas enligt angivna artikel. Ordföranden får inte rösta.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta om den föreslagna ändringen.
KOMMISSIONENS FÖRORDNING (EEG) nr 147/91 av den 22 januari 1991 om definition och fastställande av toleranser för svinn av jordbruksprodukter i offentlig interventionslagring
med beaktande av rådets förordning (EEG) nr 3492/90 om fastställande av de faktorer som skall beaktas i årsredovisningarna för finansiering av interventionsåtgärder i form av offentlig lagring genom garantisektionen inom Europeiska utvecklings- och garantifonden för jordbruket(1), särskilt artikel 4 i denna, och
Denna tolerans skall fastställas för varje berörd produkt med hjälp av en enkel metod och mot bakgrund av den oidentifierbara kvantitet svinn som konstaterats i samband med lagring under senare år. Toleransnivån bör därför fastställas som en procentsats av det totala lagret.
Tidpunkten för när de finansiella följderna av tillämpningen av toleranser skall beaktas av garantisektionen inom EUGFJ bör fastställas.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från EUGFJ-kommittén.
2. Toleransen skall fastställas som en procentsats av den faktiska vikten utan emballage av de kvantiteter som placeras i lager och övertas under det aktuella räkenskapsåret, med tillägg för kvantiteter i lager i början av det aktuella räkenskapsåret. Den skall för varje produkt beräknas på grundval av de totala kvantiteter som lagras av ett interventionsorgan.
- urbening av nötkött 32 %
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE. Artikel 1
"Artikel 3
B. Slaktkroppar av andra okastrerade djur av hankön.
E. Slaktkroppar av andra djur av honkön.
2. Slaktkroppar av vuxna nötkreatur skall klassificeras genom en bedömning i följdordning av
enligt definitionerna i bilagorna 1 respektive 2.
3. Medlemsstater skall vara bemyndigade att dela upp var och en av de klasser som anges i bilagorna 1 och 2 i högst tre underklasser."
KOMMISSIONENS FÖRORDNING (EEG) nr 1781/91 av den 19 juni 1991 om ändring av förordning (EEG) nr 1014/90 om närmare tillämpningsföreskrifter för definition, beskrivning och presentation av spritdrycker
med beaktande av rådets förordning (EEG) nr 1576/89 av den 29 maj 1989 om allmänna bestämmelser för definition, beskrivning och presentation av spritdrycker(1), särskilt artikel 6.3 i denna, och med beaktande av följande:
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för genomförande av regler om spritdrycker.
2. I linje med situationen vid tiden för den här förordningens ikraftträdande får dock följande sammansatta beteckningar användas vid presentation av likörer som framställts i gemenskapen:
Artikel 2 Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Förvaltningskommittén för fjäderfäkött och ägg har inte yttrat sig inom den tid som dess ordförande bestämt.
Till och med den 31 december 1991 får aktörerna emellertid förpacka produkter som omfattas av denna förordning i förpackningsmaterial som är försett med de uppgifter som anges i gemenskapslagstiftningen eller i den nationella lagstiftning som tillämpades före denna förordnings ikraftträdande. Dessa produkter får sedan saluföras till och med den 31 december 1992."
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, och särskilt artikel 43 i detta,
Mot bakgrund av den positiva utvecklingen i fråga om harmonisering inom veterinärområdet, bör man fastställa nya bestämmelser om datorisering av veterinärförfarandena vid import och beslut 88/192/EEG bör därför upphävas.
Datorisering av veterinärförfarandena vid import bör erbjuda möjligheter för en officiell veterinär som skall avvisa en sändning vid en gränskontrollstation att på ett effektivt sätt förmedla relevanta upplysningar och också omfatta databaser med importvillkor och för import av djur och animaliska produkter.
Kommissionen bör få till uppgift att besluta om nödvändiga tillämpningsföreskrifter.
- Organisation och drift av databaser som innehåller gemenskapens importvillkor för djur och produkter.
Artikel 2
1. Det informationssystem som avses i artikel 1.1 första strecksatsen skall omfatta gränskontrollstationer, medlemsstaternas centrala myndigheter och kommissionen.
1. De databaser som avses i artikel 1 andra strecksatsen skall innehålla alla upplysningar om importvillkor för import till gemenskapen av djur och produkter och särskilt upplysningar om förteckningar över godkända tredje länder, godkända anläggningar, vidtagna skyddsåtgärder och godkända intygsförebilder.
1. De databaser som avses i artikel 1.1 tredje strecksatsen skall innehålla alla upplysningar om varje sändning av djur eller produkter som förs in till gemenskapen, särskilt om de transportvillkor för djur som fastställs i kapitel III i direktiv 91/628/EEG och resultaten av de kontroller som utförs i enlighet med direktiv 90/675/EEG och 91/496/EEG.
Den utrustning som används vid gränskontrollstationer vid tillämpning av detta beslut kan vara den som anges i artikel 2.2 i kommissionens beslut 91/398/EEG av den 19 juli 1991 om ett datoriserat nätverk som länkar samman veterinärmyndigheterna (Animo)(7).
Artikel 8
2. Följande skall läggas till i artikel 8.2:
"Den officiella veterinären skall se till att uppdatering av de databaser som avses i artikel 1 tredje strecksatsen i beslut 92/438/EG utförs."
5. Följande mening skall läggas till artikel 11.4 b:
"- aktivera det informationssystem som avses i artikel 1 första strecksatsen i beslut 92/438/EEG."
"5. Bestämmelserna i beslut 92/438/EEG skall tillämpas."
1. I artikel 4.1 skall följande strecksats läggas till:
"Den officiella veterinären skall se till att all uppdatering av de databaser som avses i artikel 1 tredje strecksatsen i beslut 92/438/EEG utförs."
"- aktivera det informationssystem som avses i artikel 1 första strecksatsen i beslut 92/438/EEG".
"4. Bestämmelserna i beslut 92/438/EEG skall tillämpas."
I artikel 11 i direktiv 91/628/EEG skall följande stycke läggas till:
"Artikel 37 a
Tillämpningsföreskrifter för detta beslut skall vid behov antas i enlighet med det förfarande som fastställs i artikel 13.
2. När det förfarande som anges i denna artikel skall tillämpas skall ordföranden utan dröjsmål hänskjuta ärendet till kommittén antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
b) Om förslaget inte är förenligt med kommitténs yttrande, eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Bestämmelserna i detta beslut skall ses över före den 1 juli 1995 för att ta hänsyn till den tekniska utvecklingen och för att göra nödvändiga förbättringar särskilt med hänsyn till ny utveckling som redan kan ha konstaterats i de mest avancerade medlemsstaterna.
KOMMISSIONENS BESLUT av den 25 september 1992 om fastställande av samarbetsformer mellan Animo datacentrum och medlemsstaterna (92/486/EEG)
med beaktande av rådets beslut 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden(1), senast ändrat genom direktiv 92/60/EEG(2) och särskilt artikel 20.3 i detta, och med beaktande av följande:
Bestämmelserna i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Varje medlemsstat skall i enlighet med sina nationella bestämmelser utse en myndighet som skall vara ansvarig för samordningen mellan de interna myndigheterna i varje enskild medlemsstat.
De behöriga myndigheterna i medlemsstaterna skall säkerställa det kontrakt som avses i artikel 1
- innehåller en klausul om uppsägning med sex månaders varsel,
a) 300 ecu per år per lokal enhet enligt förteckningen i kommissionens beslut 92/175/EEG(6).
Medlemsstaterna förpliktar sig att endast åberopa den uppsägningsklausul som avses i artikel 2 tredje strecksatsen enligt det förfarande som fastställs i artikel 20.3 i direktiv 90/425/EEG.
Artikel 5
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
I enlighet med vad som föreskrivs i artikel 6 i direktiv 89/107/EEG har Vetenskapliga livsmedelskommittén rådfrågats om de föreskrifter som kan förväntas påverka folkhälsan.
Artikel 1
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 juni 1993 och skall genast underrätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
För att skydda människan och miljön från potentiella risker som kan uppstå när nya ämnen släpps ut på marknaden är det nödvändigt att besluta om lämpliga åtgärder och särskilt att ändra och skärpa bestämmelserna i rådets direktiv 67/548/EEG(4) senast ändrat genom direktiv 90/517/EEG(5).
För att kunna bedöma inverkan på människan och miljön bör ämnet göras till föremål för en riskbedömning. Enhetliga principer för denna riskbedömning bör fastställas.
Enligt rådets direktiv 86/609/EEG av den 24 november 1986 om tillnärmning av medlemsstaternas lagar och andra författningar om skydd av djur som används för försök och andra vetenskapliga ändamål(8) är det önskvärt att nedbringa till ett minimum antalet djur som används i djurförsök. Alla lämpliga åtgärder bör vidtas för att undvika att redan gjorda djurförsök upprepas.
Till skydd för allmänheten och särskilt de arbetstagare som använder ämnena bör bestämmelser om klassificering och märkning av ämnen antas på gemenskapsnivå.
Det är önskvärt att införa ännu en farosymbol, "miljöfarligt", som skall anges på förpackningen.
Kommissionen bör ha befogenhet att anpassa samtliga bilagor till direktiv 67/548/EEG till den tekniska utvecklingen.
Direktiv 67/548/EEG ändras på följande sätt:
c) bedömning av de anmälda ämnenas potentiella risker för människan och miljön,
b) Kosmetiska produkter som avses i direktiv 76/768/EEG(3), senast ändrat genom direktiv 86/199/EEG(4).
e) Djurfoder.
h) Andra ämnen eller preparat, för vilka tillämpas gemenskapsförfaranden för anmälan eller godkännande och för vilka kraven är likvärdiga med dem som föreskrivs i detta direktiv.
- transport av farliga ämnen på järnväg, väg eller inre vattenväg, till sjöss eller med flyg,
1. I detta direktiv används följande beteckningar med de betydelser som här anges:
c) polymer: ett ämne bestående av molekyler, som kännetecknas av sammankoppling av en eller fler monomerenheter och utgörs av en enkel viktmajoritet molekyler som innehåller åtminstone tre monomerenheter kovalent bundna till åtminstone en annan monomerenhet eller annan reaktant, och som består av mindre än en enkel viktmajoritet molekyler med samma molekylvikt. Molekylerna skall vara fördelade över en rad molekylvikter, där skillnaden i molekylvikt främst kan hänföras till skillnader i antalet monomerenheter. I denna definition avses med "monomerenhet" en monomers form i en polymer efter reaktionen.
e) släppa ut på marknaden: tillhandahållande till tredje part. I detta direktiv skall import till gemenskapens tullområde likställas med att släppa ut på marknaden.
h) EINECS: (European Inventory of Existing Commercial Substances): Europeisk förteckning över befintliga marknadsförda ämnen. Denna lista utgör en fullständig förteckning över de ämnen som anses finnas på den gemensamma marknaden den 18 september 1981.
b) oxiderande ämnen och preparat: ämnen och preparat som i kontakt med andra ämnen, i synnerhet brandfarliga, ger upphov till en kraftig exoterm reaktion,
- ämnen och preparat som kan bli heta och slutligen fatta eld i kontakt med luft av rumstemperatur utan tillförsel av energi, eller
- ämnen och preparat som i kontakt med vatten eller fuktig luft utvecklar brandfarliga gaser i farliga mängder.
g) Giftiga ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden i små mängder leder till döden eller ger akuta eller kroniska skador.
j) Irriterande ämnen och preparat: ämnen och preparat som ej är frätande men som vid direkt, långvarig eller upprepad kontakt med hud eller slemhinnor kan orsaka inflammation.
m) Mutagena ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan orsaka eller öka förekomsten av ärftliga genetiska defekter.
Artikel 3
För vissa ämnen i EINECS kan det emellertid redan finnas existerande uppgifter som har tagits fram med andra metoder än de som förskrivs i bilaga 5. Huruvida dessa uppgifter är tillräckliga för att ämnet skall kunna klassificeras och märkas eller om produkten måste testas på nytt i enlighet med bilaga 5 avgörs från fall till fall, varvid bland annat beaktas att det är angeläget att begränsa antalet djurförsök med ryggradsdjur.
Artikel 4
2. De allmänna principerna för klassificering och märkning av ämnen och preparat skall tillämpas enligt kriterierna i bilaga 6(1), utom i fall då andra krav för farliga preparat anges i särskilda direktiv.
Medlemsstaternas förpliktelser
- förpackats och märkts i enlighet med artikel 22-25, enligt kriterierna i bilaga 6 och i enlighet med resultaten av de tester som föreskrivs i bilaga 7 och 8, utom i fråga om preparat för vilka det finns särskilda bestämmelser i andra direktiv.
Artikel 6
Artikel 7
- En dokumentation med de uppgifter som krävs för att bedöma de förutsebara risker, såväl omedelbara som fördröjda, som ämnet kan medföra för människan och miljön, tillsammans med all tillgänglig information som är relevant för en sådan bedömning. Som ett minimum skall ingå de uppgifter och de undersökningsresultat som avses i bilaga 7 A, tillsammans med en detaljerad och fullständig beskrivning av de företagna undersökningarna och av de metoder som använts eller litteraturreferenser till dem.
- Endast beträffande farliga ämnen, ett förslag till säkerhetsdatablad enligt artikel 27.
Utöver ovan nämnda uppgifter kan anmälaren också tillhandahålla en preliminär riskbedömning som han gjort i enlighet med principerna i artikel 3.2.
- när den mängd av ämnet som släppts ut på marknaden uppnår 100 ton per år och tillverkare, eller när den totala mängd av ämnet som släppts ut på marknaden uppnår 500 ton per tillverkare, varvid den behöriga myndigheten skall kräva att de kompletterande tester/undersökningar som föreskrivs i bilaga 8 nivå 1 skall utföras inom den tid som den behöriga myndigheten bestämmer, utom i fall då anmälaren kan visa att en viss test/undersökning är olämplig eller att en alternativ test/undersökning är att föredra,
Artikel 8
- En dokumentation med de uppgifter som krävs för en bedömning av de förutsebara risker, såväl omedelbara som fördröjda, som ämnet kan medföra för människan och miljön, tillsammans med all tillgänglig information som är relevant för en sådan bedömning. Som ett minimum skall i dokumentationen ingå de uppgifter och de undersökningsresultat som avses i bilaga 7 B, tillsammans med en detaljerad och fullständig beskrivning av de företagna undersökningarna och av de metoder som använts eller litteraturreferenser till dem, om den medlemsstat där anmälan lämnas så kräver.
3. Om en anmälare har lämnat en begränsad dokumentation enligt punkt 2, skall han, innan den mängd av ämnet som släpps ut på marknaden uppnår 100 kg per år och tillverkare eller den totala mängd som släpps ut på marknaden per tillverkare uppnår 500 kg, förse den behöriga myndigheten med de kompletterande uppgifter som krävs för att rapporten skall motsvara kraven i bilaga 7 B.
Artikel 9
Artikel 10
Om den behöriga myndigheten anser att dokumentationen inte uppfyller kraven i direktivet och meddelar anmälaren detta enligt artikel 16.2, får ämnet släppas ut på marknaden tidigast 60 dagar efter det att myndigheten mottagit de uppgifter som behövs för att anmälan skall överensstämma med direktivet.
Artikel 11
Artikel 12
Artikel 13
- Ämnen som finns upptagna i EINECS.
- Aktiva ingredienser som endast används i de farmaceutiska produkter som avses i artikel 1.2 a. Som sådana räknas inte kemiska halvfabrikat.
- Polymerer med undantag för sådana som i kombinerad form innehåller minst 2 % av ett ämne som inte finns upptaget i EINECS.
En tillverkare eller importör som begagnar sig av detta undantag måste föra löpande anteckningar av vilka framgår ämnets identitet, märkningsinformation, mängder samt en förteckning över kunder. Dessa uppgifter skall på begäran ställas till förfogande för den behöriga myndigheten i den medlemsstat där tillverkningen, importen eller den vetenskapliga forskningen och utvecklingen sker.
3. De ämnen som avses i punkt 2 skall, i den mån anmälaren rimligen kan förväntas känna till deras farliga egenskaper, förpackas och provisoriskt märkas av tillverkaren eller dennes representant i enlighet med reglerna i artikel 22-25 och enligt kriterierna i bilaga 6.
Kompletterande uppgifter
- nya rön angående ämnets påverkan på människan eller miljön, som han rimligen kan förväntas känna till,
- alla förändringar i hans ställning (tillverkare eller importör).
Ny anmälan av samma ämne och åtgärder för att undvika upprepade tester på ryggradsdjur
a) om det ämne han avser att anmäla redan är anmält, och
b) Ämnet är tidigare anmält.
3. Anmälare av ett ämne som i enlighet med punkt 1 och 2 har kommit överens om utbyte av information enligt bilaga 7 skall också vidta alla nödvändiga åtgärder för att nå en överenskommelse om utbyte av information som erhållits från tester på ryggradsdjur och som lämnats i enlighet med artikel 7.2.
Myndigheternas rättigheter och skyldigheter
Dessutom får de behöriga myndigheterna
- vidta lämpliga åtgärder som hänför sig till en säker användning av ämnet, tills sådana bestämmelser införs på gemenskapsnivå.
Om dokumentationen godtas skall myndigheten samtidigt meddela anmälaren det officiella nummer som tilldelats hans anmälan. Om dokumentationen inte godtas skall myndigheten meddela anmälaren vilka kompletterande uppgifter som krävs för att dokumentationen skall anses överensstämma med detta direktiv.
5. Förfarandet i artikel 28 skall följas när ett förslag till klassificering och märkning fastställs eller ändras.
Kommissionens roll i anmälningsförfarandet
Den riskbedömning som avses i artikel 16.1 eller en sammanfattning av denna bedömning skall vidarebefordras till kommissionen så snart den är tillgänglig.
1. När dokumentation och de uppgifter som avses i artikel 17 kommit in till kommissionen skall den vidarebefordra kopior till medlemsstaterna. Kommissionen kan också om den anser det lämpligt vidarebefordra annat relevant material som den har insamlat i enlighet med detta direktiv.
Sekretess
a) ämnets handelsnamn,
d) möjliga sätt att göra ämnet ofarligt,
i) vad gäller ämnen i bilaga 1, analysmetoder som gör det möjligt att upptäcka ett farligt ämne när det kommit ut i miljön och bestämma direkt exponering hos människor.
Uppgifter som godtagits som konfidentiella av den myndighet som mottagit anmälningshandlingarna från anmälaren skall behandlas som konfidentiella även av andra behöriga myndigheter och av kommissionen.
4. Sekretessbelagda uppgifter som kommer till kommissionens eller en medlemsstats kännedom skall hållas hemliga.
- dock får röjas för sådana personer som är direkt engagerade i administrativa eller rättsliga förfaranden som innefattar sanktioner och som genomförs i syfte att kontrollera ämnen som släppts ut på marknaden, samt för personer som deltar i eller skall höras i samband med lagstiftningsarbete.
1. De uppgifter som lämnats i enlighet med artikel 17 och 18.1 kan vidarebefordras till kommissionen och medlemsstaterna i sammanfattad form.
Artikel 21
Artikel 22
a) Förpackningen skall vara så utformad och konstruerad att allt läckage förhindras. Detta krav skall inte gälla om särskilda säkerhetsanordningar föreskrivs.
d) Återförslutbara stängningsanordningar skall vara så konstruerade att de kan återförslutas upprepade gånger utan att innehållet kan komma ut.
2. Medlemsstaterna kan också föreskriva att förpackningarna ursprungligen skall vara förslutna och plomberade på ett sådant sätt att plomberingen bryts när förpackningen öppnas första gången.
Artikel 23
2. På varje förpackning skall tydligt och outplånligt anges följande:
c) Farosymboler, om sådana fastställts, och upplysning om typen av fara som är förenad med ämnets användning. Farosymbolens utformning och ordalydelsen i faroangivelsen skall följa vad som föreskrivs i bilaga 2(1). Symbolen skall vara tryckt i svart på orangegul botten. Farosymboler och faroangivelser skall överensstämma med dem som anges i bilaga 1. För farliga ämnen som ännu inte finns upptagna i bilaga 1 skall faroangivelser och farobeteckningar tilldelas enligt reglerna i bilaga 6.
- Om symbolen C är obligatorisk behöver inte symbolen X anges.
e) Standardfraser (S-fraser) med skyddsanvisningar för en säker användning av ämnet. S-fraserna skall överensstämma med vad som anges i bilaga 4. De S-fraser som skall användas för varje ämne anges i bilaga 1. För farliga ämnen som ännu inte finns upptagna i bilaga 1 skall S-fraser tilldelas enligt reglerna i bilaga 6.
3. För irriterande, mycket brandfarliga, brandfarliga och oxiderande ämnen behöver R-fraser och S-fraser inte anges om förpackningen inte innehåller mer än 125 ml. Detta gäller också för samma mängd farliga ämnen som inte säljs av detaljister till allmänheten.
Tillämpningen av märkningskraven
3. Etiketten - eller i fall som avses i punkt 2, förpackningen - skall ha sådan färg och utformning att farosymbolen och dess bakgrund framträder tydligt.
5. Medlemsstaterna får föreskriva att farliga ämnen som släpps ut på marknaden i det egna landet skall vara märkta på landets eget eller egna språk.
b) När det bara finns en förpackning
För farliga ämnen som inte lämnar en medlemsstats territorium får märkning ske enligt nationella regler i stället för enligt internationella regler för transport av farliga ämnen.
1. Artikel 22-24 skall inte gälla sådana bestämmelser som avser ammunition eller explosiva varor som släpps ut på marknaden för att vid användningen ge explosioner eller pyrotekniska effekter.
a) tillåta att märkning enligt artikel 23 anbringas på annat lämpligt sätt om förpackningen är för liten eller på annat sätt olämplig för att märkas i enlighet med artikel 24.1 och 24.2,
Detta undantag innebär inte att andra symboler, faroangivelser, R-fraser eller S-fraser än dem som föreskrivs i detta direktiv får användas.
Reklam
Säkerhetsdatablad
2. Allmänna regler för säkerhetsdatabladens utarbetande, distribution, innehåll och utformning skall fastställas i enlighet med förfarandet i artikel 29.4 a.
Nödvändiga ändringar för att anpassa bilagorna till den tekniska utvecklingen skall beslutas i enlighet med förfarandet i artikel 29.
1. Kommissionen skall biträdas av en kommitté bestående av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Artikel 30
Artikel 31
2. Kommissionen skall fatta ett beslut i enlighet med förfarandet i artikel 29.4 a.
Rapporter
2. Artikel 24, 25 och 27 skall betecknas artikel 33, 34 och 35.
- Bilaga 6 del 1 A ersätts av bilaga 2 till detta direktiv.
- I artikel 10.3 och 11 ersätts "artikel 8c" med "artikel 28".
- I artikel 10.3 och 11 ersätts "artikel 8 c" av "artikel 28".
- I artikel 3.3 ersätts "cancerogena, mutagena och teratogena verkningar" med "cancerogena och mutagena egenskaper samt verkningar på fortplantningen".
"o) Preparat skall anses som skadliga för fortplantningen och tilldelas åtminstone farosymbolen och faroangivelsen "giftigt" om de innehåller ett ämne som har sådana verkningar och som tilldelas minst en av de R-fraser enligt bilaga 6 till direktiv 67/548/EEG som betecknar ämnen som skadliga för fortplantningen i kategori 1, i koncentrationer som motsvarar eller överstiger
- Artikel 3.5 p skall ha följande lydelse:
- den koncentration som anges i punkt 6 i bilaga 1 (tabell VI) till detta direktiv, om ämnet inte är upptaget i bilaga 1 till direktiv 67/548/EEG eller förekommer där, men utan angivande av koncentrationsgränser."
- antingen de koncentrationer som anges i bilaga 1 till direktiv 67/548/EEG för ämnet i fråga, eller
- I artikel 6.3 ersätts "artikel 21" av "artikel 28".
- Följande punkt infogas i artikel 8:
- I artikel 10, 14.2 och 15 ersätts "artikel 21" med "artikel 28".
Artikel 3
3. Medlemsstaterna skall till kommissionen överlämna texterna till nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
RÅDETS DIREKTIV 92/77/EEG av den 19 oktober 1992 med tillägg till det gemensamma systemet för mervärdesskatt och med ändring av direktiv 77/388/EEG (harmonisering av mervärdesskattesatser)
med beaktande av kommissionens förslag(),
med beaktande av följande: Fullbordandet av den inre marknaden, vilket är ett av de grundläggande målen för gemenskapen, kräver som ett första steg att tull- och skattekontrollerna vid gränserna avskaffas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 12.3 skall ersättas med följande:
Medlemsstaterna får även tillämpa en eller två reducerade skattesatser. Dessa får inte vara lägre än 5 % och får endast avse tillhandahållande av sådana varor och tjänster som anges i bilaga H.
d) Regler om beskattningen av andra jordbruksprodukter än sådana som tillhör kategori 1 i bilaga H skall enhälligt antas av rådet före den 31 december 1994 på grundval av kommissionens förslag.
Medlemsstaterna kommer från och med den 1 januari 1993 att vidta alla nödvändiga åtgärder för att bekämpa bedrägeri och annan oredlighet på detta område. Dessa åtgärder får inbegripa införandet av ett system för redovisning av mervärdesskatt på tillhandahållande av guld mellan skattskyldiga personer inom samma medlemsstat, vilket låter köparen betala skatt för säljarens räkning och samtidigt ger köparen rätt till avdrag med samma belopp som ingående skatt."
"På grundval av kommissionens rapport skall rådet vartannat år, med början 1994, granska omfattningen av de reducerade skattesatserna. Rådet kan på kommissionens förslag enhälligt besluta att ändra i förteckningen över varor och tjänster i bilaga H."
a) Undantag med återbetalning av skatt som erlagts i föregående led, och reducerade skattesatser som är lägre än den minimiskattesats som lagts fast i artikel 12.3 vad gäller de reducerade skattesatser som var i kraft den 1 januari 1991 och som står i överensstämmelse med gemenskapslagstiftningen och uppfyller de villkor som stadgas i artikel 17 sista strecksatsen i rådets andra direktiv av den 11 april 1967, får bibehållas.
b) Medlemsstater som den 1 januari 1991 på andra varor och tjänster än sådana som anges i bilaga H i överensstämmelse med gemenskapslagstiftningen tillämpade regler om undantag med återbetalning av skatt som erlagts i föregående led eller reducerade skattesatser som var lägre än det minimum som lagts fast i artikel 12.3 vad gäller reducerade skattesatser får tillämpa den reducerade skattesatsen eller den ena av de två reducerade skattesatser som nämns i artikel 12.3 på sådana varor eller tjänster.
e) Medlemsstater som den 1 januari 1991 tillämpade en reducerad skattesats på andra varor och tjänster än sådana som specificeras i bilaga H får tillämpa denna reducerade skattesats eller en av de två reducerade skattesatser som nämns i artikel 12.3 på dessa områden, förutsatt att skattesatsen inte understiger 12 %.
5. Bilaga H i bilagan till detta direktiv skall bifogas.
När medlemsstaterna antar dessa åtgärder, skall besluten innehålla en hänvisning till detta direktiv eller åtföljas av sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Vissa av bestämmelserna skiljer sig mellan de olika språkversionerna. Dessa bestämmelser bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Ett mindre fel i formen (dock inte svullnader eller missbildningar).
- Ett mindre "Haywardmärke" i form av längsgående linjer men utan förhöjning."
2. Under "III. Bestämmelser angående storlekssortering" skall första stycket ha följande lydelse:
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
För att uppnå en effektiv administration är det önskvärt att de upplysningar som skall ingå i en anhållan om fastställande av gränsvärde för farmakologiskt verksamma ämnen i veterinärmedicinska produkter i enlighet med förordning (EEG) nr 2377/90 så mycket som möjligt motsvarar de uppgifter som skall lämnas till medlemsstaterna i en ansökan om tillstånd att släppa ut en veterinärmedicinsk produkt på marknaden, vilken inges i enlighet med artikel 5 i rådets direktiv 81/851/EEG av den 28 september 1981 om tillnärmning av medlemsstaternas lagstiftning om veterinärmedicinska läkemedel(3), ändrat genom direktiv 90/676/EEG(4).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 113 i detta,
I denna resolution fastställs särskilt genomförandet av åtgärder för att främja jordbruksexport från dessa länder till gemenskapen, och närmare bestämmelser för tillämpningen av åtgärderna måste därför definieras.
Artikel 1
3. Som ett resultat av tillämpningen av punkt 1 skall tullarna upphävas helt när de når en nivå på 2 % eller mindre.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 42 och 43 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
Det förefaller därför lämpligt att särskilt erkänna de organisationer som kan påvisa att de är representativa på regional eller interregional nivå eller på gemenskapsnivå och som aktivt strävar efter att förverkliga de ovan nämnda målen. Ett sådant erkännande bör kunna beviljas av medlemsstaten eller av kommissionen, beroende på hur omfattande branschorganisationens verksamhet är.
För att säkerställa att programmet fungerar på ett riktigt sätt bör det etableras ett nära samarbete mellan medlemsstaterna och kommissionen, varvid kommissionen bör ha en stående kontrollbefogenhet, särskilt vad gäller erkännandet av de branschorganisationer som arbetar på regional eller interregional nivå och vad gäller de avtal och de samordnade förfaranden som dessa organisationer tillämpar.
3. bedriver några av följande verksamheter på regional nivå i en eller flera regioner inom gemenskapen eller inom hela gemenskapen, och därvid beaktar konsumentintressena:
c) Förbättrande av kunskapen om och insynen i marknaden.
f) Forskning om metoder som gör det möjligt att begränsa användningen av växtskyddsmedel samtidigt som produktens kvalitet säkerställs och jorden skyddas.
Kommissionen kan inom 60 dagar efter medlemsstatens anmälan motsätta sig ett erkännande.
b) branschorganisationen överträder ett eller flera av de förbud som anges i artikel 7.3, utan att det påverkar tillämpningen av rättsliga förfaranden enligt nationell lagstiftning,
Artikel 4
b) har bildats i överensstämmelse med en medlemsstats lagstiftning eller gemenskapsrätten
Kommissionen skall fatta beslut om erkännande inom tre månader efter det att den har mottagit ansökan och all information.
Kommissionen skall offentliggöra namnen på de branschorganisationer som erkänts i C-serien av Europeiska gemenskapernas officiella tidning och samtidigt ange inom vilken ekonomisk sektor eller geografiskt område de är verksamma och vilka av de i artikel 2 angivna verksamheterna som de bedriver. Återkallanden av erkännanden skall också offentliggöras.
Artikel 7
- avtalen och de samordnade förfarandena anmälts till kommissionen, och
3. Avtal och samordnade förfaranden skall under alla omständigheter förklaras vara oförenliga med gemenskapens bestämmelser om de
- kan medföra en snedvridning av konkurrensen som inte är nödvändig för att uppnå målen för den gemensamma jordbrukspolitik som branschåtgärderna syftar till.
Detta beslut får inte träda i kraft tidigare än det datum då den berörda branschorganisationen underrättats om beslutet, såvida inte branschorganisationen har lämnat felaktiga uppgifter eller missbrukat det undantag som anges i punkt 1.
Branschorganisationerna måste för att få utvidga tillämpningsområdet för sina bestämmelser företräda minst två tredjedelar av den berörda produktionen eller handeln. Om den föreslagna utvidgningen berör flera regioner, måste branschorganisationerna påvisa att de uppnår en viss minsta nivå i fråga om representativitet inom varje näringsgren och varje region.
b) Fastställande av minimikvantiteter.
e) Användande av certifierat utsäde och kontroll av produktkvaliteten.
1. Då det gäller bestämmelser antagna av branschorganisationer som erkänts av medlemsstaterna, svarar medlemsstaterna för att berörda intressenter informeras genom offentliggörande av de avtal och samordnade förfaranden vars tillämpning avses utvidgas till att omfatta enskilda eller grupper som inte tillhör någon branschorganisation i en viss region eller grupp av regioner.
3. Kommissionen skall i C-serien av Europeiska gemenskapernas officiella tidning offentliggöra de bestämmelser för vilka utvidgad tillämpning som begärts av de branschorganisationer som den erkänt enligt artikel 4. Efter offentliggörandet skall medlemsstaterna och de berörda intressenterna ha två månader på sig att lämna sina synpunkter.
5. Kommissionen skall senast tre månader efter medlemsstatens anmälan fatta beslut i enlighet med punkt 2 och, i det fall punkt 3 är tillämplig, senast fem månader efter offentliggörandet av ansökan om utvidgad tillämpning av bestämmelserna i Europeiska gemenskapernas officiella tidning.
- begränsar frihandeln, eller
7. Om bestämmelser i enlighet med denna artikel gjorts bindande för näringsidkare som inte är medlemmar i en branschorganisation, får medlemsstaten eller kommissionen, det som är lämpligast från fall till fall, besluta att enskilda eller grupper som inte är medlemmar skall betala till organisationen hela eller del av medlemsavgiften, utom för den del av avgiften som används för att täcka administrativa kostnader i samband med tillämpningen av bestämmelserna eller de samordnade förfarandena.
2. De verksamheter som avses i denna artikel skall anknyta till något eller några av följande områden:
- Forskning om odlingsmetoder som medger en minskad användning av växtskyddsmedel och garanterar att jorden och miljön skyddas.
Artikel 11
Tillämpningsföreskrifter till denna förordning skall fastställas i enlighet med det förfarande som anges i artikel 23 i förordning (EEG) nr 2075/92(6).
Som ett led i anpassningen av den gemensamma jordbrukspolitiken bör diversifiering av jordbruksproduktionen uppmuntras så att det blir bättre balans mellan tillgång och efterfrågan. Stimulerad efterfrågan på produkter med särskilda egenskaper skulle kunna vara till stort gagn för landsbygdens ekonomi, särskilt i mindre gynnade eller avlägset belägna trakter, genom att denna förbättras och odlarnas inkomster och avfolkning förebyggs i dessa trakter.
Märkningen av jordbruksprodukter och livsmedel är underkastad de allmänna regler som anges i rådets direktiv 79/112/EEG av den 18 december 1978 om tillnärmning av medlemsstaternas lagstiftning om märkning, presentation och reklam i fråga om livsmedel(4). Med hänsyn till den särskilda beskaffenheten hos jordbruksprodukter och livsmedel bör speciella regler införas om jordbruksprodukter och livsmedel från ett särskilt geografiskt område.
De planerade reglerna bör ta hänsyn till redan befintlig gemenskapslagstiftning om vin och spritdrycker som ger högre skyddsnivå.
En jordbruksprodukt eller ett livsmedel som bär en sådan beteckning måste uppfylla vissa villkor som anges i en specifikation.
Med hänsyn till den tekniska utvecklingen bör det finnas förfaranden som gör det möjligt att ändra specifikationen efter det att registrering skett eller att ur registret avföra den geografiska beteckningen eller ursprungsbeteckningen för en jordbruksprodukt eller ett livsmedel om produkten eller livsmedlet inte längre överensstämmer med den specifikation som låg till grund när skyddet beviljades för beteckningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Denna förordning skall dock inte tillämpas på vinprodukter och spritdrycker.
3. Rådets direktiv 83/189/EEG av den 28 mars 1983 om ett informationsförfarande beträffande tekniska standarder och föreskrifter(5) skall inte tillämpas på ursprungsbeteckningar och geografiska beteckningar som omfattas av denna förordning.
b) geografisk beteckning: Namn på en region, en ort eller i undantagsfall ett land, använt för att beskriva en jordbruksprodukt eller ett livsmedel
3. Vissa traditionella geografiska eller icke-geografiska namn på en jordbruksprodukt eller ett livsmedel som härstammar från en viss region eller viss ort och som uppfyller de villkor som avses i andra strecksatsen i punkt 2 a skall också betraktas som ursprungsbeteckningar.
och - särskilda villkor gäller för framställningen av råvarorna,
6. För att kunna behandlas som ursprungsbeteckningar enligt punkt 4 måste beteckningarna i fråga godkännas eller redan vara godkända som ursprungsbeteckningar med nationellt skydd av ifrågavarande medlemsstat eller, om denna stat inte har ett sådant skyddssystem, ha vedertagen traditionell prägel och enastående rykte och anseende.
1. Namn som har blivit generiska får inte registreras.
- förhållandena i den medlemsstat som namnet kommer från och i de områden där produkten eller livsmedlet konsumeras,
När en ansökan om registrering avslås i enlighet med det förfarande som föreskrivs i artikel 6 och 7 av den anledningen att namnet har blivit generiskt, skall kommissionen offentliggöra beslutet i Europeiska gemenskapernas officiella tidning.
Artikel 4
a) Produktens eller livsmedlets benämning, inkl. ursprungsbeteckning eller geografisk beteckning.
d) Uppgifter som styrker att produkten eller livsmedlet härstammar från det geografiska området, i den mening som avses i artikel 2.2 a respektive b.
g) Uppgifter om de kontrollorgan som föreskrivs i artikel 10.
Artikel 5
4. Ansökningen skall inges till den medlemsstat där det ifrågavarande geografiska området är beläget.
1. Inom sex månader skall kommissionen genom en formell granskning kontrollera att registreringsansökningen innehåller alla de uppgifter som föreskrivs i artikel 4.
3. Om ingen invändning framställs till kommissionen i enlighet med artikel 7 skall namnet införas i ett register, "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar", som kommissionen skall föra och som skall uppta namn på de grupper och kontrollorgan som berörs.
- de ändringar i registret som företagits i enlighet med artikel 9 och 11.
Artikel 7
3. Varje lagligen berörd intresserad fysisk eller juridisk person får framställa invändning mot den begärda registreringen genom att inge en vederbörligen underbyggd skrivelse till den behöriga myndigheten i det medlemsstat där han bor eller verkar. Denna myndighet skall vidta de åtgärder som är nödvändiga för att pröva invändningen inom den fastställda tidsfristen.
- Invändningen visar att den föreslagna registreringen skulle äventyra överlevnaden för ett identiskt eller snarlikt namn eller varumärke eller för produkter som lagligen marknadsförs vid den tidpunkt då denna förordning offentliggörs i Europeiska gemenskapernas officiella tidning.
a) Om förlikning har träffats, skall medlemsstaterna i fråga underrätta kommissionen om alla de faktorer som gjorde förlikningen möjlig jämte om sökandens och invändarens yttranden. När ingen ändring gjorts av de uppgifter som kommissionen har erhållit enligt artikel 5, skall kommissionen gå vidare i enlighet med artikel 6.4. Om någon ändring har gjorts skall kommissionen på nytt inleda det förfarande som föreskrivs i artikel 7.
Beteckningarna PDO, PGI eller motsvarande traditionella nationella angivelser för skyddade ursprungsbeteckningar eller skyddade geografiska beteckningar får endast användas på jordbruksprodukter och livsmedel som uppfyller denna förordnings krav.
Artikel 6 skall därvid äga motsvarande tillämpning.
1. Medlemsstaterna skall se till att, inom sex månader från det att denna förordning har trätt i kraft, kontrollorgan har upprättats med uppgift att säkerställa att jordbruksprodukter och livsmedel som bär en skyddad beteckning uppfyller de krav som fastställts i produktspecifikationen.
Om ett kontrollorgan anlitar ett annat organ för vissa kontrollåtgärder, måste detta senare kunna ge samma garantier. I sådana fall skall den utsedda myndigheter respektive det godkända privata organet fortfarande vara ansvarigt gentemot medlemsstaten för alla kontrollåtgärder.
5. En medlemsstat måste dra tillbaka godkännandet av ett kontrollorgan om de kriterier som avses i punkt 2 och 3 inte längre är uppfyllda. Medlemsstaten skall underrätta kommissionen härom, och denna skall i Europeiska gemenskapernas officiella tidning offentliggöra en reviderad förteckning över godkända kontrollorgan.
Artikel 11
3. Om avvikelser från produktspecifikationen upprepas och medlemsstaterna i fråga inte kunnat träffa förlikning skall en underbyggd ansökan inges till kommissionen.
1. Utan att påverka tillämpningen av internationella överenskommelser kan denna förordning också tillämpas på en jordbruksprodukt eller ett livsmedel från tredje land under följande förutsättningar:
Bruk av sådana beteckningar skall vara tillåtet endast om produktens ursprungsland är klart och tydligt angivet i märkningen.
a) Varje direkt eller indirekt kommersiellt bruk av den skyddade beteckningen för produkter som inte omfattas av registreringen i den mån dessa produkter är jämförbara med de produkter som har registrerats under beteckningen i fråga eller detta bruk av den skyddade beteckningen innebär att dennas anseende exploateras.
d) Annat beteende som är ägnat att vilseleda allmänheten om produktens verkliga ursprung.
- att produkterna lagligen har marknadsförts med användning av sådana uttryck under minst fem år före den dag denna förordning offentliggörs, och
3. Skyddade beteckningar får inte bli generiska.
Varumärkesregistrering som har skett i strid med vad som sägs i föregående stycke skall förklaras ogiltig.
Kommissionen skall biträdas av en kommitté som skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Detaljregler för tillämpningen av denna förordning skall fastställas enligt det förfarande som föreskrivs i artikel 15.
2. I enlighet med det förfarande som föreskrivs i artikel 15 skall kommissionen registrera de av de beteckningar som avses i punkt 1 vilka uppfyller kraven i artikel 2 och 4. Artikel 7 skall inte vara tillämplig. Generiska beteckningar skall dock inte registrerats.
Denna förordning träder i kraft tolv månader efter det att den har publicerats i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: I kommissionens förordning (EEG) nr 1124/77(5), senast ändrad genom förordning (EEG) nr 3049/89(6), fastställs de destinationszoner som skall användas vid fastställandet av exportbidrag och avgifter vid export av spannmål och ris.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
I bilagan till denna förordning anges de destinationszoner som skall användas vid fastställande av differentierade exportbidrag och exportavgifter för de produkter som förtecknas i artikel 1 punkt a, b och c i förordning (EEG) nr 2727/75 och i artikel 1 punkt a och b i förordning (EEG) nr 1418/76.
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Erfarenheten har visat att bestämmelserna om frivillig angivelse av värpdagen bör ändras. Det bör entydigt klargöras att då värpdag anges, skall denna anges både på äggen och på förpackningarna. De villkor på vilka förpackningsanläggningar, som får äggen från produktionsenheter belägna på samma ställe, får ange värpdag bör bringas i överensstämmelse med de villkor som gäller för andra förpackningsanläggningar om man använder slutna behållare. Bestämmelser bör införas om märkning av ägg med värpdag då denna inte infaller på en arbetsdag.
Bestämmelserna om användningen av termen "extra" bör ändras i syfte att specificera villkoren för att denna term ska få förekomma på förpackningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Utöver förpackningsdagen får aktören vid förpackningstillfället ange rekommenderad sista försäljningsdag eller bäst före-dag på äggen eller på förpackningen, eller på bådadera.
4. De datum som avses i denna artikel skall anges med två siffergrupper som i följande ordning utvisar:
Om värpdagen anges på ägg och äggförpackningar i enlighet med bestämmelserna i artikel 15, skall följande villkor gälla:
- på begäran av denna myndighet, antalet värphönor som respektive producent håller.
- den dagliga äggproduktionen från varje hönshus,
- värpdagen,
4 De behållare som avses i punkt 3 skall öppnas på förpackningsanläggningen omedelbart innan klassificeringen påbörjas. Alla ägg från en enskild behållare skall klassificeras och förpackas utan avbrott. För ägg som skall märkas med värpdagen gäller att detta datum skall stämplas på äggen vid klassificeringen eller omedelbart efter denna.
- klassificeras och förpackas i enlighet med föreskrifterna i artikel 1.6, eller
6 Förpackningsanläggningar skall föra separata register över
- antalet sålda ägg och/eller vikten på dessa, uppdelade efter viktklass och köpare, med angivande av köparens namn och adress.
- I punkt 1 skall inledningsfrasen ersättas med följande:
- Punkt 6 skall ersättas med följande:
"c) märkningen 'ÄGG TILL LIVSMEDELSINDUSTRIN', skriven med 2 cm höga bokstäver på ett eller flera av gemenskapens språk."
3. Stora förpackningar som innehåller små förpackningar märks med texten `FÖRPACKNING INNEHÅLLANDE SMÅ FÖRPACKNINGAR MED "EXTRA" ÄGG`, med 2 cm höga versala bokstäver på ett eller flera av gemenskapens språk."
8 Bilaga 1 skall ersättas med bilagan till denna förordning.
KOMMISSIONENS FÖRORDNING (EEG) nr 3224/92 av den 4 november 1992 om rättelse av förordning (EEG) nr 2342/92 om import av renrasiga avelsdjur av nötkreatur från tredje land och beviljande av exportbidrag för detta samt om upphävande av förordning (EEG) nr 1544/79
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött(1), senast ändrad genom förordning (EEG) nr 2066/92(2), särskilt artiklarna 10.5 och 18.6 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR BESLUTAT FÖLJANDE
Artikel 3
Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
Större öppenhet krävs beträffande de beståndsdelar som används i kosmetiska produkter för att dessa skall kunna släppas ut på marknaden utan något föregående förfarande, för att de nödvändiga uppgifterna om slutprodukterna endast skall behövas finnas tillgängliga på tillverkningsstället eller på den plats dit de först importeras inom gemenskapen samt för att ge konsumenterna ökad information. En sådan öppenhet bör kunna uppnås om en kosmetisk produkts användningsområde och beståndsdelar anges på förpackningen. Om det av praktiska skäl är omöjligt att återge beståndsdelar och eventuella varningstexter beträffande användningen på behållaren eller den yttre förpackningen bör dessa uppgifter bifogas, så att konsumenterna får tillgång till all nödvändig information.
Kommissionen bör ha befogenhet att ändra bilagorna 1 och 8 till direktiv 76/768/EEG med hänsyn till dessas informativa och tekniska karaktär.
Direktiv 76/768/EEG ändras på följande sätt:
Kosmetiska produkter som släpps ut på marknaden inom gemenskapen får inte kunna skada människors hälsa vid normal eller rimligen förutsebar användning, varvid följande särskilt skall beaktas: presentationen av produkten, märkning, eventuella bruksanvisningar och anvisningar för kvittblivning samt eventuella andra anvisningar eller upplysningar som lämnas av tillverkaren eller hans representant eller av annan person som är ansvarig för att produkten släpps ut på gemenskapsmarknaden.
"i) beståndsdelar eller kombinationer av beståndsdelar som utprovats på djur efter den 1 januari 1998 för att uppfylla kraven i detta direktiv.
4. Följande artikel skall införas:
I denna artikel avses med beståndsdel i kosmetika varje kemiskt ämne eller beredning av syntetiskt eller naturligt ursprung, med undantag av parfym och aromatiska blandningar, som används i sammansättningen av kosmetiska produkter.
- varje beståndsdels identitet, särskilt dess kemiska benämning, CTFA-benämning, benämning i Europeiska farmakopén, den internationella generiska benämning som rekommenderas av världshälsoorganisationen, Einecs-, IUPAC-, CAS- och färgindexnummer samt den generiska benämning som avses i artikel 7.2,
3. Kommissionen skall offentliggöra inventeringen och uppdatera den regelbundet med det förfarande som fastställs i artikel 10. Inventeringen skall vara vägledande, d. v. s. inte betraktas som en uttömmande förteckning över de ämnen som är godkända för användning i kosmetiska produkter."
6. Artikel 6.1 d skall ersättas med följande:
"f) Produktens funktion, om detta inte tydligt framgår av presentationen av produkten.
- Föroreningar i de använda råvarorna.
Parfym, aromatiska sammansättningar och råvaror till dessa skall betecknas med orden "parfym" eller "aromämne". Beståndsdelar som förekommer i lägre koncentrationer än 1 % får nämnas i valfri ordning efter de beståndsdelar som förekommer i högre koncentrationer. Färgämnen får upptas i valfri ordning efter övriga beståndsdelar med de färgindexnummer eller benämningar som används i bilaga 4.
Kommissionen skall senast den 14 december 1994 i enlighet med förfarande i artikel 10 fastställa på vilka kriterier och villkor en tillverkare för att bevara affärshemligheter får ansöka om att befrias från kravet att uppta en eller flera beståndsdelar i den nämnda förteckningen."
I fråga om tvål, kulor med badskum och andra små produkter vilkas storlek eller form gör det omöjligt att uppta de uppgifter som avses i g på en etikett, remsa, tejp eller kort eller på en bipacksedel skall dessa uppgifter skyltas i omedelbar närhet av den kosmetiska produktens säljbehållare."
10. Artikel 7.2 skall ersättas med följande:
"3. Dessutom kan en medlemsstat kräva att snar och adekvat medicinsk behandling i händelse av betänkligheter skall göras möjlig genom att lämplig och tillräcklig information om vilka ämnen som ingår i den kosmetiska produkten finns tillgänglig för den behöriga myndigheten, som skall garantera att informationen endast används för att underlätta sådan medicinsk behandling.
"Artikel 7a
b) Fysikaliskkemiska och mikrobiologiska specifikationer för råvarorna och slutprodukten och renhetskriterier och kriterier för mikrobiologisk kontroll avseende den kosmetiska produkten.
Om samma produkt tillverkas på flera platser inom gemenskapen får tillverkaren välja att hålla informationen tillgänglig endast på en av dessa platser. Om så sker, samt om en begäran om detta riktas till honom i kontrollsyfte, skall han vara skyldig att ange den plats han valt till den eller de berörda tillsynsmyndigheterna.
g) Bevisning för den verkan som den kosmetiska produkten uppges ha, om detta är motiverat med hänsyn till arten av denna verkan eller av produkt.
4. Tillverkaren eller dennes representant eller den person för vars räkning en kosmetisk produkt tillverkas eller den som är ansvarig för att en importerad kosmetisk produkt släpps ut på gemenskapsmarknaden skall till den behöriga myndigheten i medlemsstaten meddela adressen till den plats där de kosmetiska produkterna tillverkas eller dit de först importeras inom gemenskapen, innan dessa produkter får släppas ut på gemenskapsmarknaden.
"2. Den gemensamma nomenklaturen för beståndsdelar i kosmetiska produkter och de ändringar som, efter samråd med Vetenskapliga kosmetologikommittén, har bedömts nödvändiga för att anpassa bilagorna med hänsyn till den tekniska utvecklingen skall fastställas på lämpligt sätt med samma förfarande."
1. Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att säkerställa att, från och med den 1 januari 1997, varken tillverkare eller importörer som är etablerade inom gemenskapen släpper ut kosmetiska produkter, som inte uppfyller kraven i detta direktiv, på marknaden.
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 14 juni 1995. De skall genast underrätta kommissionen om detta.
Artikel 4
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
i samarbete med Europaparlamentet(2),
Direktiv 93/39/EEG(7) innehåller bestämmelser för den fortsatta administrationen av godkännanden för försäljning, som medlemsstaterna har meddelat efter yttrande från Kommittén för farmaceutiska specialiteter enligt direktiv 87/22/EEG.
I rättssäkerhetens intresse bör bestämmelser fastställas för den fortsatta granskningen av ansökningar om godkännande för försäljning, som före den 1 januari 1995 föreläggs Kommittén för farmaceutiska specialiteter eller Kommittén för veterinärmedicinska läkemedel enligt direktiv 87/22/EEG.
Direktiv 87/22/EEG skall upphöra att gälla med verkan från och med den 1 januari 1995.
Artikel 3
Artikel 4
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av yttrandet från Ekonomiska och sociala kommittén(3), och
Nationella lagar om skydd av djur vid tidpunkten för slakt eller avlivning påverkar konkurrensvillkoren och följaktligen också hur den gemensamma marknaden för jordbruksprodukter fungerar.
Det är emellertid nödvändigt att tillåta att tekniska och vetenskapliga experiment utförs samt att ta hänsyn till de särskilda krav som vissa religiösa ceremonier ställer.
I samband med detta skall gemenskapens handlande vara i enlighet med subsidiarietsprincipen i artikel 3b i fördraget.
2. Det skall inte gälla för
- vilda djur som avlivas i enlighet med artikel 3 i direktiv 92/45/EEG.
6. Avlivning: Varje metod som leder till att ett djur avlider.
Den religiösa myndigheten i en medlemsstat för vars räkning slakt utförs skall emellertid ha befogenhet att tillämpa och övervaka särskilda bestämmelser i samband med slakt enligt vissa religiösa ceremonier. I fråga om dessa bestämmelser skall denna myndighet vara underställd den officiella veterinären, enligt definitionen i artikel 2 i direktiv 64/433/EEG.
KAPITEL II Krav för slakterier
Artikel 5
b) fasthållas i enlighet med bilaga B,
2. Kraven i punkt 1 c skall inte tillämpas beträffande djur som slaktas med särskilda metoder som krävs i samband med vissa religiösa ceremonier.
1. Instrument, fasthållningsanordningar och annan utrustning och anläggningar som används vid bedövning och avlivning skall utformas, konstrueras, underhållas och användas på ett sådant sätt att bedövningen eller avlivningen sker snabbt och effektivt i enlighet med bestämmelserna i detta direktiv. Den behöriga myndigheten skall kontrollera att instrument, fasthållningsanordningar och annan utrustning som används vid bedövning eller avlivning är i överensstämmelse med ovanstående principer och skall regelbundet kontrollera att de är i gott skick och kan uppfylla denna målsättning.
Förflyttning, uppstallning, fasthållning, slakt eller avlivning av djur får endast utföras av personer som har nödvändiga kunskaper och yrkesskicklighet för att utföra arbetet humant och effektivt i enlighet med kraven i detta direktiv.
Den behöriga myndigheten skall ansvara för att det utförs besiktningar och kontroller av slakterier och skall vid alla tidpunkter ha fritt tillträde till slakteriernas alla delar för att säkerställa att bestämmelserna i detta direktiv efterlevs. Besiktningarna och kontrollerna får dock genomföras samtidigt som kontroller som genomförs i andra syften.
1. När de djur som avses i artikel 5.1 slaktas utanför slakterier skall artikel 5.1 b, 5.1 c och 5.1 d tillämpas.
1. När de djur som avses i artikel 5.1 skall slaktas eller avlivas vid sjukdomsbekämpning skall detta utföras i enlighet med bilaga E.
Artikel 11
Skadade eller sjuka djur måste slaktas eller avlivas på stället. Den behöriga myndigheten kan emellertid tillåta transport av skadade eller sjuka djur för slakt eller avlivning under förutsättning att detta inte innebär ytterligare lidande för djuren.
1. Rådet skall, om nödvändigt, genom kvalificerad majoritet på kommissionens förslag anta andra bestämmelser om skydd av djur vid tidpunkten för slakt eller avlivning än de som omfattas av detta direktiv.
- pistol med skarp ammunition, där kulan drivs in i hjärnan, eller andra gaser än de som avses i bilaga C eller kombinationer av dessa som används vid bedövning, särskilt koldioxid vid bedövning av fjäderfä,
Rådet skall ta ställning till dessa förslag med kvalificerad majoritet.
ii) nödvändig gaskoncentration och exponeringstid vid bedövning av de olika berörda arterna.
1. Kommissionens experter får, i den mån detta är nödvändigt för att säkerställa en enhetlig tillämpning av detta direktiv, utföra kontroller på plats. De kan i detta syfte kontrollera ett representativt urval av anläggningar för att säkerställa att den behöriga myndigheten kontrollerar att dessa anläggningar uppfyller kraven i detta direktiv.
3. Den medlemsstat på vars område kontrollen genomförs skall ge experterna all nödvändig hjälp i deras tjänsteutövning.
Vid besiktning av slakterier eller anläggningar i tredje land vilka har bemyndigats eller skall bemyndigas att exportera till gemenskapen i enlighet med gemenskapsbestämmelser, skall kommissionens experter säkerställa att de djur som avses i artikel 5 har slaktats under villkor som minst garanterar samma humana behandling som den som fastställs i detta direktiv.
1. Vid hänvisning till det förfarande som fastställs i denna artikel skall frågan utan dröjsmål hänskjutas till Ständiga veterinärkommittén av dess ordförande, antingen på dennes eget initiativ eller på anmodan av en representant för en medlemsstat.
b) Om de avsedda åtgärderna inte är förenliga med kommitténs yttrande, eller om inget yttrande avges, skall kommissionen utan dröjsmål förelägga rådet ett förslag om de åtgärder som skall vidtas. Rådet skall fatta beslut med kvalificerad majoritet.
Direktiv 74/577/EEG skall upphöra att gälla från och med den 1 januari 1995.
När medlemsstaterna antar dessa lagar och andra författningar skall de innehålla en hänvisning till detta direktiv eller vid offentliggörandet åtföljas av en sådan hänvisning. Närmare regler för denna hänvisning skall fastställas av medlemsstaterna.
Artikel 19
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
efter samråd med Rådgivande kommittén för kulturföremål, och
Exportlicenser måste upprättas på ett av gemenskapens officiella språk.
2. Användning av exportlicens får inte på något sätt påverka de förpliktelser som är förbundna med exportformaliteter eller därtill knutna handlingar.
2. Formulären skall vara 210 × 297 mm.
- för att låta trycka formulären som skall vara försedda med tryckeriets namn och adress eller identifieringsmärke,
Användning av licens
2. I punkt 1 förstås med sändning antingen ett enda kulturföremål eller ett antal kulturföremål.
Formulären skall bestå av tre exemplar, varav
- ett exemplar märkt nr 3 skall återsändas till den utfärdande myndigheten.
2. Ansökan skall åtföljas av
4. Om tillämpningen av punkterna 2 och 3 orsakar kostnader skall dessa bäras av den som ansöker om exportlicens.
Följande skall framläggas till stöd för exportdeklarationen:
Artikel 8
Artikel 9
3. När en exportlicens löper ut utan att ha använts skall innehavaren omedelbart återsända de exemplar han har i sin ägo till den utfärdande myndigheten.
Artikel 11
KOMMISSIONENS FÖRORDNING (EEG) nr 1785/93 av den 30 juni 1993 om de avgörande faktorerna för tillämpning av jordbruksomräkningskurser inom textilsektorn
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas avseende den gemensamma jordbrukspolitiken(1), särskilt artikel 6.2 i denna, och
Enligt artikel 10.1 och 10.2 i förordning (EEG) nr 1068/93 skall de avgörande faktorerna för minimipriset och för stödet till bomull vara de som anges i artikel 15 i förordning (EEG) nr 1201/89. Det bör dock ges möjlighet att förutfastställa jordbruksomräkningskurserna för stödet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 3
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
I rådets förordning (EEG) nr 1600/92(6), ändrad genom kommissionens förordning (EEG) nr 3714/92(7), fastställs ett stöd för den lokala produktionen av matpotatis på Madeira och för sättpotatis och endiver på Azorerna. Dessa stödbelopp bör justeras enligt ovan nämnda bestämmelser.
Artikel 1
RÅDETS FÖRORDNING (EEG) nr 2617/93 av den 21 september 1993 om ändring av förordning (EEG) nr 1907/90 om vissa handelsnormer för ägg
med beaktande av rådets förordning (EEG) nr 2771/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för ägg(1), särskilt artikel 2.2 i denna,
Bestämmelserna i fråga om direkta leveranser från producenter till förpackningsanläggningar, vissa marknader och livsmedelsindustriföretag bör också gälla sådana leveranser till andra industriföretag.
Erfarenheten har visat att bestämmelserna om datummärkning på ägg av klass A och på de äggförpackningar som innehåller sådana ägg bör ändras så att det krävs ett obligatoriskt angivande av datum för minsta hållbarhetstid på samma sätt som för andra livsmedel, i överensstämmelse med rådets direktiv 79/112/EEG av den 18 december 1978 om tillnärmning av medlemsstaternas lagstiftning om märkning, presentation och reklam i fråga om livsmedel(4). I syfte att underlätta kontroll bör även förpackningen till importerade ägg av klass A ha en märkning som anger förpackningsdatum.
Förordning (EEG) nr 1907/90 ändras på följande sätt:
3. I artiklarna 6.1 och 8.3 skall ordet "livsmedelsindustri" ersättas med "livsmedelsindustriföretag som godkänts i enlighet med direktiv 89/437/EEG."
5. Artikel 10.1 a skall ersättas med följande:
"e) Datum för minsta hållbarhetstid 'bäst-före-datum` åtföljt av lämpliga förvaringsinstruktioner för ägg av klass A, och förpackningsdag för ägg av andra klasser."
8. Artikel 13.2 skall ersättas med följande:
Kommissionen skall i enlighet med förfarandet i artikel 17 i förordning (EEG) nr 2771/75 föreskriva de övergångs-bestämmelser som behövs för genomförandet av den här förordningen, särskilt i fråga om de bestämmelser som gäller användningen av befintligt förpackningsmaterial.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
Även om det i första hand är medlemsstaterna som ansvarar för kontrollen, bör kommissionen också försöka se till att medlemsstaterna opartiskt kontrollerar och förebygger överträdelser. Kommissionen bör därför ges de finansiella medel samt rättskipnings- och lagstiftningsmedel som tillåter den att utföra detta uppdrag så effektivt som möjligt.
Politiken avseende förvaltning av fiskeresurserna, som särskilt bygger på totala tillåtna fångstmängder (TAC), fångstkvoter och tekniska åtgärder bör också omfatta förvaltning av fiskeansträngningen, som innebär att fiskeverksamheten och fiskekapaciteten övervakas.
I samband med införandet av den gemensamma fiskeripolitiken är det nödvändigt med åtgärder för att kontrollera de fartyg som för ett tredje lands flagg och befinner sig i gemenskapens farvatten. Det behövs särskilt ett system som gör det möjligt att följa fartygens rörelser och motta meddelanden om vilka arter som fartyget har ombord, utan att detta påverkar rätten till oskadlig genomfart genom territorialvattnet och friheten att navigera i fiskezonen om 200 sjömil.
Landningsmedlemsstaten måste kunna övervaka landningarna på sitt territorium; därför bör de fiskefartyg som är registrerade i andra medlemsstater informera landningsmedlemsstaten om sin avsikt att landa på dess territorium.
För att säkerställa att gemenskapens handelsåtgärder och åtgärder för bevarande respekteras bör alla fiskeprodukter som importeras till gemenskapen eller landas där, fram till dess att den första försäljningen äger rum, åtföljas av ett transportdokument som anger deras ursprung.
Medlemsstaterna måste hållas underrättade om resultaten av sina fartygs verksamhet i vatten som lyder under tredje lands jurisdiktion eller på internationellt vatten. Skyldigheten att föra loggbok och avge landnings- och omlastningsdeklaration bör därför också gälla för befälhavarna på dessa fartyg. De uppgifter som medlemsstaterna samlar in bör översändas till kommissionen.
När en medlemsstats kvot förbrukats, eller när själva TAC:en är förbrukad, måste kommissionen fatta beslut om förbud mot fiske.
För att säkerställa att de åtgärder som vidtagits förvaltas effektivt är det nödvändigt att införa en deklarationsordning som överensstämmer med de mål och strategier som fastställs i artikel 8 i förordning (EEG) nr 3760/92, vilken är tillämplig på en medlemsstat som överskridit sin kvot.
För att säkerställa granskningens objektivitet är det viktigt att gemenskapens inspektörer under vissa omständigheter får göra självständiga inspektioner utan att förvarna för att granska de kontroller som gjorts av de behöriga myndigheterna i medlemsstaterna. Sådana inspektioner får aldrig omfatta kontroll av privatpersoner.
Medlemsstaterna bör regelbundet avlägga rapport till kommissionen om sin inspektionsverksamhet och om vilka åtgärder som vidtas vid brott mot gemenskapens bestämmelser.
Denna förordning bör inte inverka på sådana nationella kontrollbestämmelser som, även om de hör till dennas tillämpningsområde, sträcker sig utanför förordningens minimiföreskrifter, förutsatt att de nationella bestämmelserna är förenliga med gemenskapsrätten.
Bestämmelserna i vissa artiklar bör träda i kraft den 1 januari 1999 i den mån de berör fisket i Medelhavet, där den gemensamma fiskeripolitiken ännu inte är helt genomförd.
- strukturåtgärderna,
2. I detta syfte skall varje medlemsstat i enlighet med gemenskapsbestämmelserna vidta nödvändiga åtgärder för att säkerställa systemets effektivitet. Den skall ställa tillräckliga medel till sina behöriga myndigheters förfogande, så att de kan genomföra den inspektion och kontroll som fastställs i denna förordning.
2. De fiskefartyg som kan bedriva fiske under ett tredje lands flagg och fiska i vatten som lyder under en medlemsstats överhöghet eller jurisdiktion skall ingå i ett system, där fartygets rörelser kan följas och uppgifter kan fås om vilka fångster som finns ombord.
4. För att inspektionen skall bli så effektiv och ekonomisk som möjligt skall medlemsstaterna samordna sin kontrollverksamhet. De kan därför utarbeta gemensamma inspektionsprogram som gör det möjligt att kontrollera gemenskapens fiskefartyg i de i punkterna 1 och 3 nämnda farvattnen. Medlemsstaterna skall vidta sådana åtgärder som gör det möjligt för deras behöriga myndigheter och kommissionen att regelbundet och ömsesidigt hålla varandra underrättade om den erfarenhet som vunnits.
2. För att utvärdera vilken teknik som skall användas och vilka fartyg som skall omfattas av nämnda system skall medlemsstaterna i samarbete med kommissionen genomföra vissa pilotprojekt före den 30 juni 1995. Medlemsstaterna skall därför se till att ett system för fortlöpande lokalisering av vissa kategorier av fiskefartyg inom gemenskapen införs, som arbetar från en land- eller satellitbaserad basstation och använder sig av satellitkommunikation för dataöverföringen.
Om fiskefartygen befinner sig i farvatten som lyder under en annan medlemsstats överhöghet eller jurisdiktion skall flaggmedlemsstaten se till att de behöriga myndigheterna i den berörda medlemsstaten omgående underrättas om detta.
2. De ansvariga för de fiskefartyg, lokaler eller transportmedel som skall inspekteras skall medverka till att underlätta den inspektion som skall genomföras i överensstämmelse med punkt 1.
a) identifiering av officiellt utsedda inspektörer, inspektionsfartyg och andra liknande inspektionsmedel som en medlemsstat kan utnyttja,
d) den rapport som inspektörerna skall sammanställa efter varje inspektion ombord,
g) registrering av uppgifter rörande fiskefartygens position och överföring av dessa uppgifter till medlemsstaterna och kommissionen,
1. Befälhavarna på sådana fiskefartyg inom gemenskapen som fiskar arter ur ett bestånd eller en grupp av bestånd skall föra loggbok, i vilken de skall ange vilka fångstmängder som finns ombord av varje art, datum och plats (statistisk rektangel ICES) för dessa fångster och vilken typ av fiskeredskap som använts.
4. Befälhavarna på gemenskapens fiskefartyg skall undantas från kraven i punkterna 1 och 3 om fartygets största längd understiger 10 m.
Varje medlemsstat skall därför utarbeta en provtagningsplan, som skall lämnas till kommissionen. Resultaten av de kontroller som görs skall regelbundet meddelas kommissionen.
Artikel 7
- vilka mängder av varje art som skall landas.
Artikel 8
3. Varje medlemsstat skall genom stickprovskontroller övervaka den verksamhet som bedrivs av de fiskefartyg som är undantagna från kraven i punkt 1 för att säkerställa att dessa fartyg följer gällande bestämmelser inom gemenskapen.
Artikel 9
3. De avräkningsnotor som avses i punkterna 1 och 2 skall minst innehålla följande uppgifter:
- Destinationen för de eventuella produkter som dragits tillbaka från marknaden (biprodukter, mänsklig komsumtion, förädling).
4. Dessa avräkningsnotor skall fyllas i och översändas i enlighet med landningsmedlemsstatens lagstiftning på sådant sätt och enligt sådana försäljningsvillkor att följande uppgifter kan inkluderas:
- Hamn och datum för landningen.
7. Kommissionen kan i enlighet med förfarandet i artikel 36 bevilja undantag från skyldigheten att presentera avräkningsnotan för medlemsstaternas behöriga myndigheter eller andra behöriga organ för de fiskprodukter som landats från vissa kategorier av gemenskapens fiskefartyg med en största längd av mindre än 10 m.
9. Närmare bestämmelser för tillämpningen av denna artikel skall antas i enlighet med det förfarande som anges i artikel 36.
b) Varje medlemsstat skall se till att befälhavaren på ett fiskefartyg som för ett tredje lands flagg eller är registrerat i ett tredje land, eller dennes ställföreträdare, vid landningen lämnar in en deklaration till myndigheterna i den medlemsstat vars landningsplatser han utnyttjar med uppgift om landade mängder och datum och plats för varje fångst; för deklarationens riktighet ansvarar befälhavaren eller dennes ställföreträdare.
Medlemsstaterna skall fastställa tillämpningsföreskrifter för punkt 1 c och anmäla dem till kommissionen.
Artikel 11
- direktlandar sådana fångstmängder utanför gemenskapens territorium,
Befälhavaren på mottagarfartyget skall förvara uppgifterna om storleken på de fångster ur ett bestånd eller en grupp av bestånd inom en TAC eller kvot vilka tagits emot vid en omlastning, datumet när de togs emot och fartyget som lastade om fångsterna till mottagarfartyget. Denna skyldighet skall anses vara uppfylld när kopior förvaras av de omlastningsdeklarationer som är utfärdade i enlighet med de närmare bestämmelserna om medlemsstaternas registrering av uppgifter om fiskefångster.
Befälhavarna på mottagarfartyget och ovannämnda tredje fartyg skall låta de behöriga myndigheterna kontrollera riktigheten av de uppgifter som krävs enligt denna punkt.
Artikel 12
1. Alla fiskeprodukter som importeras till gemenskapen eller landas där, såväl icke beredda som beredda ombord, vilka transporteras till en annan plats än landnings- eller införselplatsen, skall åtföljas av ett dokument utfärdat av transportören fram till dess att den första försäljningen ägt rum.
b) försändelsens eller försändelsernas destination och transportmedlet,
4. Transportföretaget skall undantas från sin skyldighet enligt punkt 1 om något av följande villkor är uppfyllt:
5. En medlemsstats behöriga myndigheter kan bevilja undantag från skyldigheten enligt punkt 1 om fiskmängderna transporteras innanför hamnområdet eller högst 20 km från landningsplatsen.
Artikel 14
3. Undantag kan göras från skyldigheten att behandla uppgifter om vilka mängder som landats av vissa kategorier av fartyg som omfattas av undantagen i artiklarna 7 och 8 eller vilka mängder som landats i hamnar som inte har en tillräckligt utvecklad administrativ struktur för att kunna registrera landningarna om en medlemsstat lämnar in en begäran om detta till kommissionen inom tolv månader efter det att denna förordning trätt i kraft. Ett sådant undantag kan beviljas om registreringen av dessa data skulle vara en oproportionerligt stor belastning för de nationella myndigheterna i förhållande till de totala mängder som landats, och om de landade arterna säljs lokalt. Varje medlemsstat skall upprätta en förteckning över de hamnar och fartyg som uppfyller kraven för ett sådant undantag och sända denna till kommissionen.
1. Före den 15 i varje månad skall varje medlemsstat genom dataöverföring anmäla till kommissionen vilka mängder ur varje bestånd eller grupp av bestånd som omfattas av en TAC eller kvot som landats under föregående månad, samt ge kommissionen alla de upplysningar som erhållits enligt artiklarna 11 och 12.
När fångsterna ur bestånd eller grupper av bestånd som omfattas av TAC:er eller kvoter riskerar att nå nivån för gällande TAC:er eller kvoter skall medlemsstaterna på kommissionens begäran lämna mer ingående upplysningar eller lämna sådana oftare än vad som krävs enligt denna punkt.
4. Varje medlemsstat skall före utgången av den första månaden i varje kvartal genom dataöverföring anmäla till kommissionen vilka mängder som landats under föregående kvartal av andra bestånd än de som avses i punkt 1.
Denna information skall bestå av ifrågavarande fartygs namn och distriktsbeteckning, vilka fiskmängder per bestånd eller grupp av bestånd som detta fartyg landat, bjudit ut till försäljning eller lastat om samt dagen och platsen för landningen, den första utbjudningen till försäljning eller omlastningen. Denna information skall överlämnas inom fyra arbetsdagar räknat från medlemsstatens förfrågan, eller inom en längre tidsfrist, som denna medlemsstat eller landningsmedlemsstaten kan fastställa.
1. Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa att fångsterna av sådana arter som deras fartyg tar såväl i farvatten som lyder under ett tredje lands överhöghet eller jurisdiktion som på internationellt vatten utanför zongränserna övervakas, och att omlastningar och landningar av sådana fångster granskas och registreras.
- Under landning i gemenskapens hamnar skall en landningsdeklaration lämnas in till myndigheterna i den medlemsstat där landningen äger rum.
Artikel 18
Fångster som tas på internationellt vatten utanför zongränserna skall anmälas med hänvisning till det minsta statistiska område som fastställs i den internationella konventionen om fångstplats för varje art eller grupp av arter för alla bestånd som ingår i ifrågavarande fiskeverksamhet.
1. För att säkerställa att de förpliktelser som fastställs i artiklarna 3, 6, 8, 9, 10, 14 och 17 uppfylls skall varje medlemsstat införa ett system för giltighetskontroll, som skall omfatta dubbelkontroller och granskning av de uppgifter som kommit in till följd av dessa förpliktelser.
3. Om en medlemsstat inte omedelbart kan uppfylla kraven i punkt 2 med avseende på delar av eller hela sitt fiske kan kommissionen på denna medlemsstats begäran besluta att i enlighet med förfarandet i artikel 36 bevilja den en övergångsperiod på högst tre år räknat från den dag denna förordning träder i kraft.
6. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 36.
Nätredskap som finns ombord men inte används skall stuvas undan så att de inte kan användas utan vidare i enlighet med följande bestämmelser:
2. Om fångsterna ombord på något av gemenskapens fiskefartyg tagits med nät med olika minsta maskstorlek under samma resa skall artsammansättningen beräknas för varje del av den fångst som tagits under olika förhållanden.
a) inget av gemenskapens fiskefartyg som deltar i speciella typer av fiske får medföra nät med olika minsta maskstorlek under samma resa,
1. Alla fångster ur ett kvoterat bestånd eller en kvoterad grupp av bestånd, som tas av gemenskapens fiskefartyg skall skrivas av från den kvot som tilldelats flaggmedlemsstaten för gällande bestånd eller grupp av bestånd, oberoende av landningsplatsen.
I samband med bedömningen av den situation som avses i första stycket skall kommissionen informera de berörda medlemsstaterna om sannolikheten av ett fiskestopp till följd av att en TAC är förbrukad.
Om den skada som en medlemsstat lidit genom att fisket förbjudits innan dess kvot förbrukats inte avhjälpts i enlighet med artikel 9.2 i förordning nr 3760/92, skall åtgärder beslutas på det sätt som anges i artikel 36 i syfte att på ett lämpligt sätt reparera den skada som förorsakats. Dessa åtgärder kan innebära att det görs avdrag för den medlemsstat som överskridit sin kvot, tilldelning eller andel, och att de mängder som dras av på ett lämpligt sätt delas ut till de medlemsstater vars fiske stoppats innan deras kvot förbrukats. Dessa avdrag och efterföljande tilldelningar skall göras med hänsyn till i första hand de arter och zoner för vilka kvoterna, tilldelningarna eller de årliga andelarna fastställts. Dessa avdrag eller tilldelningar kan göras under det år skadan uppstår eller under något av de följande åren.
1. Om en medlemsstats behöriga myndigheter finner att ett av gemenskapens fiskefartyg allvarligt eller upprepade gånger brutit mot denna förordning kan flaggmedlemsstaten underkasta fartyget ytterligare kontroll.
1. Om kommissionen konstaterat att en medlemsstat överskridit sin kvot, tilldelning eller andel av ett bestånd eller en grupp av bestånd skall kommissionen göra avdrag från den årliga kvot, tilldelning eller andel som den medlemsstaten förfogar över. Dessa avdrag skall fastställas i enlighet med förfarandet i artikel 36.
- Eventuella fall av överfiske av samma bestånd under de föregående åren.
För att säkerställa att de mål och strategier som fastläggs av rådet i enlighet med artikel 11 i förordning (EEG) nr 3760/92 följs, särskilt mängdmålen avseende fiskekapaciteten hos gemenskapens fiskeflotta och anpassningen av fiskeflottans verksamhet, skall varje medlemsstat på sitt territorium och i de farvatten som lyder under dess överhöghet eller jurisdiktion göra regelbundna kontroller hos alla dem som berörs av genomförandet av ovan nämnda mål.
a) Omstrukturering, förnyelse och modernisering av fiskeflottan.
d) Begränsning av fiskeredskapens utformning och antal, samt deras användningssätt.
Artikel 26
b) fiskefartygens registertonnage,
2. Medlemsstaterna skall omgående meddela kommissionen vilka kontrollmetoder som används samt namn och adress till de organ som svarar för kontrollen.
- den loggbok som avses i artikel 6,
2. För detta ändamål skall medlemsstaterna upprätta databaser eller bygga ut redan existerande databaser med relevant information om fiskeflottans kapacitet och verksamhet.
Artikel 28
a) handelsstandarder, särskilt minsta storlekar,
- lagring och/eller bearbetning av produkter som återtagits från marknaden.
Kommissionen och medlemsstaternas behöriga myndigheter, samt tjänstemän och andra ombud, får inte sprida sådan information som samlas in genom tillämpningen av denna artikel som omfattas av tystnadsplikt.
1. Kommissionen skall kontrollera att medlemsstaterna tillämpar denna förordning genom att granska dokument och göra besök på platsen. Om kommissionen finner det lämpligt kan den företa granskningar utan förvarning.
a) Medlemsstaterna skall samarbeta med kommissionen för att underlätta för denna att genomföra sina uppdrag. De skall särskilt vidta alla nödvändiga åtgärder för att inspektionerna inte skall offentliggöras, vilket skulle kunna störa genomförandet av inspektionen och kontrollen.
c) Vid inspektion till havs eller från luften skall medlemsstaternas myndigheter i de fall de nationella behöriga organen skall tillvarata andra viktiga uppgifter, särskilt i samband med försvaret eller säkerheten till sjöss, ha rätt att skjuta upp eller omdirigera de inspektioner som kommissionen planerat att närvara vid. I sådana fall skall medlemsstaten samarbeta med kommissionen för att vidta alternativa åtgärder.
När gemenskapens inspektörer granskar tillämpningen av detta program är medlemsstatens ombud alltid ansvariga för dess genomförande. Gemenskapens inspektörer kan inte på eget initiativ använda sig av de inspektionsbefogenheter som anförtrotts de nationella ombuden. Dessa inspektörer har bara tillgång till fartyg eller lokaler om de ledsagas av en medlemsstats ombud.
5. Inom ramen för de besök som nämns i punkterna 2 och 3 skall kommissionens behöriga inspektörer i de ansvariga organens närvaro på platsen få tillträde till hela eller delar av informationen i de specificerade databaserna och få granska alla de dokument som är relevanta för tillämpningen av denna förordning.
1. Medlemsstaterna skall till kommissionen på dennas begäran överlämna all information om tillämpningen av denna förordning. Om kommissionen begär information skall den ange en rimlig tid inom vilken denna skall lämnas.
För att kunna delta i de inspektioner som avses i denna punkt skall kommissionens tjänstemän visa fram en skriftlig fullmakt, av vilken deras identitet och tjänstebeteckning framgår.
4. Denna artikel påverkar inte de nationella bestämmelserna om sekretess vid rättsligt förfarande.
2. De rättsliga åtgärder som vidtas med stöd av punkt 1 skall vara av sådan art att de i enlighet med tillämpliga bestämmelser i den nationella lagstiftningen effektivt berövar de ansvariga det ekonomiska utbytet av överträdelsen eller framkallar effekter som står i proportion till överträdelsens allvar, i syfte att avskräcka från ytterligare överträdelser av samma slag.
- beslag av förbjudna fiskeredskap och fångster,
- återkallande av licensen.
1. Om de behöriga myndigheterna i landnings- eller omlastningsmedlemsstaten konstaterar att en överträdelse skett mot denna förordning skall de vidta lämpliga åtgärder i enlighet med artikel 31 mot ifrågavarande fartygs befälhavare eller mot någon annan person som är ansvarig för överträdelsen.
Om landnings- eller omlastningsmedlemsstaten inte längre har motsvarande kvot till sitt förfogande skall artikel 21.4 också tillämpas, och de olovligen landade eller omlastade fiskmängderna anses motsvara omfånget av den skada som registreringsmedlemsstaten lidit på det sätt som anges i den artikeln.
2. Efter en överlåtelse av den rättsliga uppföljningen i enlighet med artikel 31.4 skall flagg- eller registreringsmedlemsstaten vidta varje sådan lämplig åtgärd som avses i artikel 31.
1. Medlemsstaterna skall till kommissionen anmäla vilka lagar och andra författningar de antagit för att förebygga och beivra lagöverträdelser.
3. Kommissionen skall förse medlemsstaterna med ett sammandrag av de upplysningar som den erhållit i enlighet med punkterna 1 och 2.
Artikel 36
Kommissionen skall besluta med omedelbar verkan. Om beslutet inte är förenligt med kommitténs yttrande skall kommissionen emellertid genast underrätta rådet. I sådana fall får kommissionen uppskjuta verkställandet av de beslutade åtgärderna under en tid som inte överstiger en månad från dagen då rådet underrättats.
1. Medlemsstaterna och kommissionen skall vidta alla nödvändiga åtgärder för att säkerställa att de uppgifter som tas emot inom ramen för denna förordning behandlas konfidentiellt.
3. Uppgifterna som utväxlas mellan medlemsstaterna och kommissionen får bara lämnas vidare till de personer i medlemsstaternas och gemenskapens institutioner vars uppgifter kräver att de har tillgång till dem; om de lämnas till andra personer skall de medlemsstater som lämnat uppgifterna uttryckligen ha givit sitt samtycke till det.
6. Bestämmelserna i punkt 1 5 får inte tolkas som ett hinder mot att de uppgifter som erhålls genom tillämpningen av denna förordning används inom ramen för sådana rättsliga åtgärder som vidtas senare på grund av att gemenskapens fiskelagstiftning inte följts. De behöriga myndigheterna i den medlemsstat som lämnar uppgifterna skall informeras om alla de fall i vilka uppgifterna används i detta syfte.
8. Bestämmelserna i punkt 1 5 får inte tolkas som ett hinder mot att allmänna upplysningar eller undersökningar offentliggörs, som inte nämner enskilda fysiska eller juridiska personer.
Artikel 38
Artikel 39
Artikel 40
Medlemsstaterna skall fram till den 1 januari 1999 undantas från skyldigheten att tillämpa bestämmelserna i artiklarna 6, 8 och 19 i fråga om fiske i Medelhavet.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av följande: I artikel 12 i förordning (EEG) nr 2019/93 föreskrivs att stöd skall beviljas de mindre Egeiska öarna för produktion av kvalitetshonung som innehåller en stor andel timjanhonung. Tillämpningsföreskrifter bör antas för förvaltning av ord-ningen och för kontroll av de villkor som rådet har uppställt.
Med hänsyn till genomförandet av denna stödordning bör undantag fastställas vad gäller sista ansökningsdag och sista utbetalningsdag för stöd för 1993 års produktion.
Artikel 1
Artikel 2
- Upprätthållande av avkastningen genom att gamla drottningar två gånger om året byts ut mot hybrider som är anpassade till området.
Artikel 3
2. Stödansökan skall minst innehålla följande uppgifter:
- Den mängd honung med stor andel timjanhonung som producerats under den period för vilken det ansöks om stöd.
Grekland skall betala ut stödet senast den 31 december under den period för vilken stöd beviljas, i proportion till den faktiska graden av genomförande av initiativprogrammet. Stöd skall inte utbetalas om genomförandegraden under-stiger 50 %.
Grekland skall, senast den 31 januari varje år, meddela kommissionen följande:
- Den sänkningskoefficient som eventuellt tillämpas.
För år 1993 får dessa uppgifter emellertid överlämnas senast den 15 mars 1994.
- Genomförandet av inititativprogrammet.
RÅDETS FÖRORDNING (EEG) nr 3089/93 av den 29 oktober 1993 om ändring av förordning (EEG) nr 2299/89 om en uppförandekod för datoriserade bokningssystem
med beaktande av kommissionens förslag (),
med beaktande av följande: Förordning (EEG) nr 2299/89 () utgör ett viktigt led i avskaffandet av snedvriden konkurrens mellan lufttrafikföretag och mellan datoriserade bokningssystem, och skyddar därigenom konsumenternas intressen.
Enligt kommissionens förordning (EEG) nr 83/91 () är fördragets artikel 85.1 inte tillämplig på överenskommelser om gemensamma inköp, gemensam utveckling och drift av datoriserade bokningssystem.
I princip konkurrerar "seat-only" eller separata lufttransportprodukter på icke-regelbunden lufttrafik direkt med de lufttransportprodukter som erbjuds på regelbundna flygningar.
De konsumenter som söker efter olika produkter bör ges möjlighet att begära textbilder för enbart regelbunden eller icke-regelbunden lufttrafik.
Det är lämpligt med en klar åtskillnad mellan ett avtal om deltagande i eller som tillåter användning av ett system och leveransen av den tekniska utrustningen, varvid leveransen omfattas av sedvanlig avtalsrätt vilket ger systemleverantören rätt att kräva att få sina direkta kostnader täckta i de fall då ett avtal om deltagande eller abonnemang sägs upp enligt bestämmelserna i denna förordning.
Konkurrensmässig likhet kommer att ökas genom att man säkerställer att de datoriserade bokningssystemen har separat juridisk identitet.
Det är önskvärt att utförliga upplysningar om avsättning, bokning och försäljning görs tillgängliga för deltagande lufttrafikföretag på ett icke diskriminerande sätt och med samma skyndsamhet. Identifiering av eller personlig information om en passagerare eller ett företag måste förbli konfidentiell. Därför skall en systemleverantör genom tekniska hjälpmedel och lämpliga säkerhetskrav, åtminstone vad gäller mjukvara, säkerställa att otillåtet tillträde till information inte kan äga rum.
Systemleverantören skall säkerställa att principerna om teknisk överensstämmelse med bestämmelserna om likhet i funktion och datasäkerhet övervakas av en oberoende kontrollant.
Förordning (EEG) nr 2299/89 ändras på följande sätt:
P varifrån den utnyttjade informationen kommer eller var den centrala databehandlingsanläggningen i fråga är belägen,
I denna förordning används följande beteckningar med de betydelser som här anges:
c) lufttransportprodukt: både separata lufttransportprodukter och kombinerade lufttransportprodukter.
P Den bedrivs så att den betjänar trafiken mellan samma, två eller flera, orter antingen
e) biljettpris: det pris som skall betalas för separata lufttransportprodukter och villkoren för när detta pris är tillämpligt.
P platstillgång,
med eller utan möjligheter till
av sådan omfattning att några av eller samtliga dessa tjänster ställs till förfogande för abonnenterna.
i) moderföretag: ett lufttrafikföretag som direkt eller indirekt, ensamt eller tillsammans med andra, äger eller effektivt kontrollerar en systemleverantör, såväl som varje lufttrafikföretag som det äger eller effektivt kontrollerar.
P rättigheter eller avtal som ger ett avgörande inflytande över sammansättningen hos företagets organ, omröstning eller andra beslut, eller som på annat sätt ger ett avgörande inflytande över driften av ett företag.
m) konsument: varje person som önskar upplysning om eller har för avsikt att köpa en lufttransportprodukt.
p) serviceförbättring: varje produkt eller tjänst som inte är en distributionstjänst och som en systemleverantör på egna vägnar erbjuder abonnenter i anslutning till ett datoriserat bokningssystem.
fordra att tilläggsvillkor godtas, som genom sin karaktär eller enligt affärssed inte har något samband med deltagandet i leverantörens datoriserade bokningssystem, och skall tillämpa samma villkor för samma servicenivå.
I sådana fall skall en systemleverantör bara ha rätt att få tillbaka de direkta kostnaderna för uppsägningen av avtalet.
"Artikel 3a
1. c) Moderföretaget skall ha rätt att utföra kontroller för att säkerställa att artikel 5.1 respekteras av det konkurrerande datoriserade bokningssystemet.
"Artikel 4
1. a) Ett datoriserat bokningssystem skall ge en textbild som är klar och som inte är diskriminerande.
1. b) En konsument skall ges möjlighet att begära primära textbilder för enbart regelbunden eller icke-regelbunden lufttrafik.
1. e) De normer som används för att rangordna informationen får inte baseras på någon faktor som direkt eller indirekt har samband med lufttrafikföretagets identitet och inte tillämpas på ett sätt som diskriminerar något deltagande lufttrafikföretag.
5. Ett datoriserat bokningssystem anses inte bryta mot bestämmelserna i denna förordning i den utsträckning som det förändrar en textbild för att tillmötesgå en konsuments specifika förfrågningar.
a) Information om enskilda bokningar skall ställas till förfogande på lika villkor för det eller de lufttrafikföretag som deltar i utförandet av den tjänst som bokningen avser och för de abonnenter som berörs av bokningen.
ii) Att sådana uppgifter får, och skall på begäran, omfatta alla deltagande lufttrafikföretag och abonnenter, men skall inte identifiera eller ge personlig information om en passagerare eller ett företag.
3. Systemleverantören skall säkerställa att bestämmelserna i punkt 1 och 2 uppfylls genom tekniska medel eller lämpliga säkerhetskrav avseende åtminstone mjukvara, på ett sådant sätt att ett eller flera av moderföretagen inte på något sätt kan få tillgång till information som ges av eller skapas för lufttrafikföretag, utom vad som tillåts enligt denna artikel.
6. I artikel 7 skall punkterna 1 och 2 ersättas med följande:
"5. a) När det konstateras allvarlig diskriminering enligt punkterna 1 och 2 får kommissionen besluta om att de datoriserade bokningssystemen skall instrueras att ändra sina metoder så att diskrimineringen upphör. Kommissionen skall genast informera medlemsstaterna om ett sådant beslut.
2. Ett moderföretag får varken direkt eller indirekt kräva att en abonnent använder ett visst datoriserat bokningssystem för att sälja eller utställa biljetter för en lufttransportprodukt som företaget självt direkt eller indirekt levererar.
"4. a) En systemleverantör får inte ställa upp oskäliga villkor i ett avtal med en abonnent om användning av dess datoriserade bokningssystem, och i synnerhet får en abonnent alltid säga upp sitt avtal med en systemleverantör med en uppsägningstid som inte behöver överstiga tre månader, dock att den tidigast får löpa ut vid utgången av det första avtalsåret.
5. En systemleverantör skall i varje abonnentavtal fastställa
6. En systemleverantör får inte ålägga en abonnent någon skyldighet att acceptera ett erbjudande om teknisk utrustning eller mjukvara, men får kräva att en utrustning eller mjukvara som är kompatibel med hans eget system används."
Fakturorna för det datoriserade bokningssystemets tjänster skall vara tillräckligt informativa för att de deltagande lufttrafikföretagen och abonnenterna skall kunna se exakt vilka tjänster de utnyttjat och avgifterna för dem. Fakturor för bokningsavgifter skall minst innehålla följande uppgifter för varje sträcka:
P Stat.
P De två orterna eller sträckan.
P Linjenummer.
P Boknings-/avbokningsindikator.
2. En systemleverantör skall på begäran lämna intresserade parter uppgifter om tillämpade metoder och avgifter, om erbjudna systemtjänster, inklusive gränssnitt, samt om de kriterier för redigering och textbildspresentation som används. Denna bestämmelse förpliktar emellertid inte en systemleverantör att lämna information som är äganderättsligt skyddad, till exempel programvara."
Bestämmelserna i artikel 5, artikel 9.5 och i bilagan till denna förordning skall inte tillämpas på ett datoriserat bokningssystem som används av ett lufttrafikföretag eller en grupp av lufttrafikföretag i dess eget (deras egna) klart markerade kontor och försäljningsdiskar."
1. Systemleverantören skall säkerställa att en oberoende kontrollant övervakar att dess datoriserade bokningssystem är tekniskt förenligt med artiklarna 4a och 6. För detta ändamål skall kontrollanten vid varje tidpunkt beviljas tillträde till de program, metoder, förfaranden och säkerhetskrav som används i de datorer eller datorsystem genom vilka systemleverantören erbjuder sina distributionstjänster. Varje systemleverantör skall minst en gång per år till kommissionen lämna sin kontrollants inspektionsrapport och slutsatser. Denna rapport skall granskas av kommissionen för att utröna om det behöver vidtas åtgärder enligt artikel 11.1.
"Artikel 22
14. Artikel 23 skall ersättas med följande:
2. Rådet skall se över tillämpningen av artiklarna 4a och 6.3 på grundval av en rapport som kommissionen skall lämna senast vid utgången av 1994."
1. Denna förordning träder i kraft den trettionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av artikel 132 i konventionen om tillämpning a
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113 i förening med artikel 228.2 i detta,
med beaktande av följande: Kommissionen har på gemenskapens vägnar förhandlat fram ett tilläggsprotokoll till interimsavtalet om handel och handelsfrågor och till Europaavtalet med Rumänien.
Artikel 1
Artikel 2
KOMMISSIONENS BESLUT av den 7 februari 1994 om ändring av rådets beslut 90/424/EEG om vissa utgifter på veterinärområdet (84/77/EG)
med beaktande av rådets beslut 90/424/EEG av den 26 juni 1990 om vissa utgifter på veterinärområdet(1), senast ändrat genom beslut 93/439/EEG(2), särskilt artikel 24.1 i detta, och med beaktande av följande:
Med hänsyn till den särskilda hälsosituationen i de franska utomeuropeiska departementen är det motiverat att lägga till nämnda sjukdomar i bilagan till beslut 90/424/EEG.
Artikel 1
- Babesios, som överförs av smittbärande insekter i de franska utomeuropeiska departementen,
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De åtgärder som föreskrivs i det här direktivet är förenliga med yttrandet från Ständiga veterinärkommittén.
Bilagorna till direktiv 89/556/EEG skall ändras enligt vad som framgår av bilagan till detta beslut.
Beslutet skall inte tillämpas på embryon som samlas, hanteras och förvaras före den 1 mars 1994.
KOMMISSIONENS BESLUT av den 23 februari 1994 om inrättande av en rådgivande samordningskommitté för förebyggande av bedrägerier (94/140/EG)
med beaktande av följande: En sund förvaltning av gemenskapens finanser förutsätter att bedrägerier som skadar gemenskapens budget motarbetas effektivt.
Kommissionen har även ett stort ansvar som ett led i sin generella uppgift att se till att gemenskapens budget tillämpas korrekt och att fördragets bestämmelser genomförs.
Eftersom kommittén kommer att behandla alla aspekter av bedrägeriproblematiken och alla medlemsstater har behov av en representation på rätt nivå som avspeglar strukturen i den egna förvaltningen, bör det läggas fast att kommittén skall bestå av två företrädare från varje medlemsstat.
1. Kommittén skall bestå av två företrädare för varje medlemsstat, vilka får biträdas av två tjänstemän från de berörda myndigheterna.
2. Kommissionen kan när den begär ett yttrande från kommittén fastställa en tidsfrist för avgivande av yttrandet.
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av ramen för den gemensamma åtgärd som Europeiska rådet enades om den 10 och 11 december 1993, och
Artikel 1
- använda sitt inflytande för att uppmuntra alla parter att ovillkorligt stödja fredsprocessen på grundval av inbjudningar till Madrid-konferensen och arbeta för att stärka demokratin och respekten för de mänskliga rättigheterna,
- utveckla sin roll i den särskilda sambandskommitté som ansvarar för samordningen av internationellt stöd till de ockuperade områdena,
c) Europeiska unionen skall
- följa utvecklingen vad avser israeliska bosättningar inom samtliga ockuperade områden och fortsätta att rikta demarscher till Israel i denna fråga.
- ett snabbt genomförande av biståndsprogrammen för utveckling av de ockuperade områdena och en palestinsk driftsbudget, i nära samråd med palestinierna och en lika nära samverkan med andra biståndsgivare,
För att aktivt och snabbt bidra till att en palestinsk polisstyrka upprättas skall
c) ett belopp på högst 10 miljoner ecu från gemenskapens budget som en brådskande åtgärd ställas till förfogande som bistånd till upprättandet av en palestinsk polisstyrka.
De praktiska arrangemangen och den finansiering som följer av denna artikel skall behandlas i ett särskilt, separat beslut.
Artikel 6
Detta beslut skall ha verkan från och med denna dag.
KOMMISSIONENS BESLUT av den 25 maj 1994 om tillämpningsföreskrifter till rådets direktiv 90/425/EEG vad avser provtagningen i samband med veterinärkontroller på bestämmelseorten (94/338/EG)
med beaktande av rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden(1), senast ändrat genom direktiv 92/118/EEG(2), särskilt artikel 5.3 i detta, och med beaktande av följande:
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Artikel 4
EUROPEISKA GEMENSKAPERNAS RÅD HAR FATTAT DETTA BESLUT
med beaktande av kommissionens förslag, och
Beslut om utsträckning av skyddet bör i största möjliga omfattning fattas av gemenskapen som helhet.
I avtalet om handelsrelaterade aspekter på immateriella rättigheter, som är ett av förhandlingsresultaten i de multilaterala handelsförhandlingarna under Uruguay-rundan och ingår i Marrakesh-slutakten av den 15 april 1994, krävs det att medlemmarna skall ge skydd åt mönster i integrerade kretsar enligt bestämmelserna i det avtalet och bestämmelserna i konventionen om skydd av immateriella rättigheter beträffande integrerade kretsar, till vilket avtalet hänvisar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) Fysiska personer som är medborgare i Canada eller som har sin vanliga vistelseort inom Canadas territorium skall behandlas som om de vore medborgare i en medlemsstat.
Detta beslut skall tillämpas från och med den 1 november 1994.
KOMMISSIONENS BESLUT av den 30 november 1994 om särskilda villkor för import av levande tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar med ursprung i Turkiet (Text av betydelse för EES) (94/777/EG)
med beaktande av rådets direktiv 91/492/EEG av den 15 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av levande tvåskaliga blötdjur(1), särskilt artikel 9 i detta, och
Ministry of Agriculture and Rural Affairs och dess laboratorier kan effektivt kontrollera tillämpningen av gällande lagar i Turkiet.
Turkiet kan tas upp i den förteckning över tredje länder som uppfyller de bestämmelser om likvärdighet som anges i artikel 9.3 a i direktiv 91/492/EEG.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
4. Varje förpackning skall ha en beständig hälsomärkning som innehåller minst följande uppgifter:
- Uppgift om upptagningsområdets och leveransanläggningens godkännandenummer.
1. Intygen enligt artikel 2.1 skall vara utfärdade på minst ett officiellt språk i den medlemsstat där kontrollerna görs.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
1. Förpackningsanläggningar som endast plockar samman produkter utan att ta bort innerförpackningen skall uppfylla tillämpliga villkor enligt bilaga B, kapitel VII punkt 1 till direktiv 77/99/EEG.
1. Produkter från de förpackningsanläggningar som avses i artikel 1.1 skall bibehålla kontrollmärket från det ursprungliga produktionsföretaget.
2. Förpackningsanläggningar skall upprätta ett särskilt registreringssystem som gör det möjligt för den behöriga myndigheten att spåra en ompaketerad produkt till ursprungsföretaget.
KOMMISSIONENS BESLUT av den 28 december 1994 om godkännande av Finlands operativa program för bekämpning av salmonella hos vissa levande djur och i animaliska produkter (94/968/EG)
med beaktande av rådets direktiv 64/432/EEG av den 26 juni 1964 om djurhälsoproblem som påverkar handeln inom gemenskapen med nötkreatur och svin(1), ändrat genom del 1 kapitel 2 avsnitt A punkt 1. h i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 10a andra stycket i detta,
med beaktande av rådets direktiv 71/118/EEG av den 15 februari 1971 om hälsoproblem som påverkar handeln med färskt fjäderfäkött(4), ändrat genom del 1 kapitel 3 punkt 3. b i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 5.4 i detta,
Detta operativa program omfattar alla de åtgärder som Finland från och med dagen för ikraftträdandet av anslutningsfördraget har åtagit sig att vidta för att bekämpa salmonella hos nötkreatur och svin för avel, produktion och slakt, avelsfjäderfä, daggamla kycklingar som skall ingå i flockar av avelsfjäderfä eller flockar av produktionsfjäderfä, värphöns (produktionsfjäderfä som föds upp för att producera konsumtionsägg), slaktfjäderfä, nötkött och griskött, fjäderfäkött och ägg till direkt konsumtion som livsmedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Det finska programmets åtgärder avseende värphöns (produktionsfjäderfä som föds upp för att producera konsumtionsägg) godkänns.
Artikel 5
Det finska programmets åtgärder avseende fjäderfäkött godkänns.
Artikel 8
Detta beslut träder i kraft om och på samma dag som anslutningsfördraget för Norge, Österrike, Finland och Sverige träder i kraft.
RÅDETS FÖRORDNING (EEG) nr 163/94 av den 24 januari 1994 om ändring av förordning (EEG) nr 386/90 om kontroll i samband med export av jordbruksprodukter som berättigar till exportbidrag eller andra belopp
med beaktande av kommissionens förslag(1),
Det framgår klart av denna rapport och av tilläggsrapporten att den bristande smidigheten hos vissa regler kan motverka förbättringar av effektiviteten i kontrollerna; riskanalyser kan komma till bättre användning om kontrollorganen har större frihet att själva bestämma på vilka områden det särskilt skall genomföras kontroller.
För att minska risken för utbyte av produkter, särskilt när det gäller exportdeklarationer som framläggs och godkänns inne i medlemsstaten eller i exportörens lokaler måste det fastställas en lägsta procentsats av representativa fysiska stickprovskontroller som skall genomföras vid utförseltullkontoret.
Artikel 1
- per kalenderår, och,
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovanstående förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
Om inte annat följer av de åtgärder som är i kraft i gemenskapen beträffande system med dubbelkontroll och med övervakning i för- och efterhand av import av textilprodukter till gemenskapen, är det lämpligt att de bindande klassificeringsbesked som getts ut av medlemsstaternas tullmyndigheter rörande klassificeringen av varor i Kombinerade nomenklaturen och som inte överensstämmer med denna förordning, fortsatt får åberopas av mottagaren under en tid av 60 dagar, enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för anpassning till tekniska framsteg av direktiven om avskaffande av tekniska handelshinder inom sektorn veterinärmedicinska läkemedel.
Bilagorna 1, 2, 3 och 4 till förordning (EEG) nr 2377/90 ändras på det sätt som anges i bilagan till den här förordningen.
KOMMISSIONENS FÖRORDNING (EG) nr 3129/94 av den 20 december 1994 om ändring av förordning (EEG) nr 2273/93 om fastställande av interventionsorter för spannmål till följd av Österrikes, Finlands och Sveriges anslutning
med beaktande av Anslutningsakten för Norge, Österrike, Finland och Sverige(1), särskilt artikel 169.2 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
KOMMISSIONENS BESLUT av den 10 februari 1995 om fastställande av särskilda villkor för import av fiskeri- och vattenbruksprodukter från Marocko (Text av betydelse för EES) (95/30/EG)
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av fiskeriprodukter (1), särskilt artikel 11.1 i detta, och med beaktande av följande:
Direction de l'élevage, ministère de l'agriculture (DEMA) i Marocko är i stånd att på ett effektivt sätt kontrollera tillämpningen av den gällande lagstiftningen.
I enlighet med artikel 11.4 c i direktiv 91/493/EEG är det viktigt att fastställa en förteckning över godkända anläggningar. Denna förteckning bör fastställas på grundval av ett meddelande till kommissionen från DEMA. Det åligger således DEMA att förvissa sig om att de villkor som fastställs för detta ändamål i artikel 11.4 i direktiv 91/493/EEG uppfylls.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Artikel 1
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I överensstämmelse med förordning (EEG) nr 2377/90 måste gränsvärden fortlöpande fastställas för högsta tillåtna restmängder för alla i gemenskapen använda farmakologiskt verkande substanser i veterinärmedicinska läkemedel avsedda att tillföras livsmedelsproducerande djur.
För kontrollen av restmängder bör vanligtvis gränsvärden för högsta tillåtna restmängder för målvävnaderna lever eller njure fastställas, för vilket är ombesörjt i tillämplig gemenskapslagstiftning; och med hänsyn till att levern och njuren emellertid ofta avlägsnas från djurkroppen vid transport inom internationell handel, bör gränsvärden för högsta tillåtna restmängder alltid fastställas även för muskel- eller fettvävnad.
Lecirelin, natrium dikloroisocyanurat, dinoprost trometamin, saltsyra, äpplesyra, l-vinsyra och dess en- och tvåbasiska salter av natrium, kalium och kalcium, bensylalkohol, etanol, n-butanol bör bilaga II tillföras till förordning (EEG) nr 2377/90.
Då det förefaller som om resthalter av MRL, vid vilken nivå som helst, i livsmedel av animaliskt ursprung utgör hälsorisk för konsumenten, bör furazolidon därför föras till bilaga IV i förordning (EEG) nr 2377/90,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
Med stöd av förordning (EEG) nr 2309/93, skall kommissionen anta de bestämmelser som krävs för det skriftliga förfarandet som avses i artiklarna 10.3 och 32.3 i den förordningen.
Artikel 1
Ordföranden skall hänskjuta ärenden till kommittén med stöd tillämpliga bestämmelser i förordning (EEG) nr 2309/93, direktiv 75/319/EEG eller direktiv 81/851/EEG.
Inom trettio dagar efter överlämnandet av förslaget till beslut skall medlemsstaterna meddela ordföranden sitt beslut att godkänna förslaget, underkänna det eller avstå från att yttra sig Medlemsstaterna kan komplettera sina beslut med skriftliga anmärkningar. En medlemsstat som inte har meddelat sina invändningar eller sitt beslut att avstå från att yttra sig inom de trettio dagarna anses ha givit förslaget sitt godkännande.
Om kommissionen finner att de skriftliga anmärkningar som lämnats av en medlemsstat inom ramen för förfarandet i artikel 3 väcker betydelsefulla nya frågor av vetenskaplig eller teknisk natur vilka inte har behandlats i Europeiska läkemedelsmyndighetens yttrande, skall ordföranden avbryta förfarandet och kommissionen hänskjuta förslaget till myndigheten för vidare behandling. Ordföranden skall underrätta kommitténs medlemmar om detta.
När en medlemsstat har tillämpat det förfarande som föreskrivs i artikel 18.4 eller 40.4 i förordning (EEG) nr 2309/93 om brådskande tillfälligt förbud mot användning av ett läkemedel inom sitt territorium, skall den tidsfrist som anges i artikel 3 förkortas till femton dagar.
Dessa handlingar måste nå adressaterna senast tio dagar före sammanträdesdagen eller, i fall enligt artikel 2 andra stycket, en månad före denna dag.
Artikel 8
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100c.3 i detta,
med beaktande av följande: Enligt artikel 100c.3 i Romfördraget skall rådet besluta om åtgärder som syftar till en enhetlig utformning av visumhandlingar före den 1 januari 1996.
Denna förordning fastställer endast de specifikationer som inte är av konfidentiell art. Dessa specifikationer skall kompletteras med andra som skall förbli hemliga för att förebygga risken för efterbildningar och förfalskningar och som inte får innefatta personliga uppgifter eller hänvisning till sådana. Behörigheten att fastställa andra specifikationer bör tillkomma kommissionen.
När det gäller de personuppgifter som skall förekomma på den enhetliga visumhandlingen enligt bilagan till denna förordning, skall hänsyn tas till medlemsstaternas bestämmelser om skydd av personuppgifter och till gemenskapslagstiftningen på området.
De visum som beviljas av medlemsstaterna i enlighet med artikel 5 utformas enligt en modell (klistermärke). De skall uppfylla specifikationerna enligt bilagan.
Artikel 3
Artikel 4
Artikel 5
- en resa genom territoriet eller transitzonen på en flygplats i denna medlemsstat eller flera medlemsstater.
2. Kommissionen skall biträdas av en kommitté bestående av företrädare för medlemsstaterna med en företrädare för kommissionen som ordförande.
b) Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om medlemsstaterna använder modellen för visumhandling för andra ändamål än dem som omfattas av artikel 5 skall de åtgärder vidtas som behövs för att undvika all förväxling med den visumhandling som beskrivs i artikel 5.
RÅDETS FÖRORDNING (EG) nr 1935/95 av den 22 juni 1995 om ändring i förordning (EEG) nr 2092/91 om ekologisk produktion av jordbruksprodukter och uppgifter därom på jordbruksprodukter och livsmedel
med beaktande av kommissionens förslag (1),
med beaktande av följande: Kommissionen har inom ramen för förordning (EEG) nr 2092/91 (4), fått ett särskilt uppdrag att före den 1 juli 1994 göra en förnyad granskning av vissa bestämmelser i nämnda förordning samt att lägga fram lämpliga förslag med tanke på dess eventuella revidering.
Den förnyade granskningen har visat att bestämmelserna om märkning av livsmedel som endast till viss del beretts med hjälp av ingredienser med jordbruksursprung som producerats med ekologiska metoder bör förbättras för att åstadkomma bättre möjligheter att framhäva den ekologiskt producerade beståndsdelen i sådana livsmedel.
Konventionellt erhållna plantor avsedda för växtproduktion bör av samma anledning kunna få användas under en övergångsperiod.
Förordning (EEG) nr 2092/91 ändras på följande sätt:
"2. `produktion`: verksamheter på gården med avseende på framställning, förpackning och ursprunglig märkning som ekologiskt producerade produkter av jordbruksprodukter som produceras på den gården."
4. Artikel 6.4 ersätts med följande text:
"9. `färdigförpackat livsmedel`: saluförd enhet såsom den definieras i artikel 1.3 b i direktiv 79/112/EEG,
7. Följande punkt läggs till artikel 5.1:
9. Artikel 5.3 med följande text:
b) alla andra ingredienser av jordbruksursprung omfattas av bilaga VI punkt C eller har godkänts provisoriskt av ett medlemsland i enlighet med någon av de vidtagna genomförandeåtgärderna, vilken, i förekommande fall, antagits i enlighet med punkt 7,
e) produkten eller dess ingredienser har inte behandlats med joniserande strålning,
Uppgifter som hänvisar till ekologisk produktion skall klart visa att de gäller en produktionsmetod inom jordbruket och skall åtföljas av en hänvisning till de åsyftade ingredienserna av jordbruksursprung om detta inte klart framgår av ingrediensförteckningen."
11. Artikel 5.5 ersätts med följande text:
b) en omställningsperiod om minst 12 månader före skörd har iakttagits,
e) för produkter som beretts efter den 1 januari 1997 skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som den leverantör som har utfört den sista beredningsåtgärden är underställd. Valet av om namn eller kodnummer skall användas åligger medlemsstaten som skall meddela sitt beslut till kommissionen."
a) minst 70 % av produktens ingredienser av jordbruksursprung är produkter eller härrör från produkter som erhållits i enlighet med de regler som anges i artikel 6 eller är importerade från tredje land inom ramen för den ordning som anges i artikel 11,
d) produkten innehåller enbart ämnen som finns förtecknade i bilaga VI, punkt A i egenskap av ingredienser som inte är av jordbruksursprung,
g) produkten har beretts eller importerats av en leverantör som är underkastad den kontroll som anges i artiklarna 8 och 9,
"6. Under en övergångsperiod som går ut den 31 december 1997, får märkning av och reklam för en produkt som anges i artikel 1.1 b och som delvis erhållits från ingredienser som inte uppfyller kraven i punkt 3 a hänvisa till ekologisk produktion om följande villkor är uppfyllda:
c) de uppgifter som hänvisar till ekologisk produktion:
d) ingredienserna och deras andelar anges i fallande storleksordning efter vikt i ingrediensförteckningen,
"8. Sådana begränsande förteckningar över de ämnen och produkter som avses i punkt 3 b, c och d, samt i punkt 5 a, b, d och e skall upprättas i enlighet med det förfarande som fastställs i artikel 14 och omfattas av punkterna A, B och C i bilaga VI."
10. En produkt som anges i artikel 1.1 får inte innehålla både en ingrediens som har erhållits i enlighet med reglerna i artikel 6 och samma ingrediens som har erhållits enligt andra regler.
"Artikel 6
b) endast produkter som består av ämnen som finns förtecknade i bilagorna I och II får användas som växtskyddsmedel, tvätt- och rengöringsmedel, gödningsmedel eller markberedningsmedel eller för varje annat ändamål som med avseende på vissa ämnen anges i bilaga II. De får endast användas på de särskilda villkor som anges i bilagorna I och II i den mån deras motsvarande användning är tillåten i vanligt jordbruk i de berörda medlemsländerna i enlighet med tillämpningen av gemenskapsbestämmelser eller enligt nationella bestämmelser som överensstämmer med gemenskapslagstiftningen,
3. a) Trots vad som sägs i punkt 1 c får utsäde och vegetativt förökningsmaterial som inte har erhållits i enlighet med den ekologiska produktionsmetoden användas under en övergångsperiod fram till den 31 december 2000 med godkännande från den behöriga myndigheten i medlemsstaten under förutsättning att användarna av sådant förökningsmaterial på ett för medlemsstatens kontrollmyndighet eller kontrollorgan tillfredsställande sätt kan visa att de på gemenskapsmarknaden inte har kunnat erhålla ett förökningsmaterial för en lämplig sort av ifrågavarande art som uppfyller kraven i stycke 2. I detta fall skall ett förökningsmaterial som inte har behandlats med andra produkter än de som anges i bilaga II punkt B användas, under förutsättning att sådant material finns på gemenskapsmarknaden. Medlemsstaterna skall anmäla godkännanden som lämnats enligt detta stycke till de andra medlemsstaterna och till kommissionen,
- bibehållande, efter den 31 december 2000, av det i a angivna undantaget i fråga om vissa arter och/eller typer av förökningsmaterial för hela eller delar av gemenskapens område,
17. Följande artikel införs efter artikel 6:
2. Den ekologiska produktionsmetoden innebär att plantor som används för produktion också skall ha producerats i enlighet med bestämmelserna i artikel 6.
b) plantorna har efter sådden inte behandlats med andra produkter än de som räknas upp i bilaga II, delarna A och B,
e) märkningen av produkter som innehåller ingredienser som härrör från sådana plantor får inte innehålla den uppgift som anges i artikel 10,
- datum för godkännandet,
- trolig varaktighet för bristsituationen,
4. c) På begäran av en medlemsstat eller på kommissionens initiativ, skall ärendet föreläggas den kommitté som avses i artikel 14. I enlighet med det förfarande som avses i artikel 14 kan beslut fattas om att återkalla eller förkorta godkännandets giltighetstid."
19. I artikel 9.1 skall orden "leverantörerna av produkter av det slag som anges i artikel 1" ersättas med orden "leverantörer som producerar, bereder eller från tredje land importerar produkter av det slag som anges i artikel 1."
22. I artikel 9.6 d ersätts orden "punkt 7-9" med orden "punkterna 7, 8, 9 och 11".
24. Följande stycke skall införas i artikel 9:
"1. Uppgift och/eller logotyp utvisande att produkterna omfattas av ett särskilt kontrollsystem som visas i bilaga V, får uteslutande ingå i märkningen av produkter av det slag som avses i artikel 1 när sådana produkter
c) säljs direkt i slutna förpackningar av producent eller beredare till slutlig konsument, eller släpps ut på marknaden som färdigförpackade livsmedel. Vid direktförsäljning av producent eller beredare till slutlig konsument är slutna förpackningar inte nödvändiga när det av märkningen klart och tydligt framgår vilken produkt det är fråga om,
27. Artikel 10.5, 10.6 och 10.7 ersätts med följande text:
1. När en medlemsstat med avseende på en produkt som härrör från en annan medlemsstat och som är försedd med de uppgifter som anges i artikel 2 och/eller bilaga V konstaterar avvikelser eller överträdelser rörande tillämpningen av denna förordning, skall den informera den medlemsstat som har utsett kontrollmyndigheten eller godkänt kontrollorganet och kommissionen om detta.
29. I artikel 11.6 a ersätts datumet den 31 juli 1995 med datumet den 31 december 2002.
31. I artikel 11 läggs följande punkt till:
"- tillämpningsföreskrifter för denna förordning."
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt motsvarande KN-nummer som anges i kolumn 2 med de motiveringar som ges i kolumn 3.
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
Förhållandena i den internationella handeln eller vissa marknaders särskilda krav kan göra det nödvändigt att differentiera bidraget med hänsyn till en bestämd produkts användning eller destination.
1. De exportbidrag som avses i artikel 55 i förordning (EEG) nr 822/87 fastställs i bilagan till den här förordningen.
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2777/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för fjäderfäkött (5), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94, särskilt artiklarna 5.4 och 8.12 i denna,
med beaktande av rådets förordning (EG) nr 3491/93 av den 13 december 1993 om vissa förfaranden vid tillämpning av Europaavtalen om upprättandet av en associering mellan Europeiska gemenskaperna och dess medlemsstater å ena sidan och Ungern, å andra sidan (9), senast ändrad genom förordning (EG) nr 3379/94 (10), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 3297/94 av den 19 december 1994 om vissa förfaranden för tillämpning av Europaavtalet om associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Slovakien, å andra sidan (13), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 3641/93 av den 20 december 1993 om vissa förfaranden vid tillämpning av interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Bulgarien, å andra sidan (18), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 1276/95 av den 29 maj 1995 om vissa förfaranden för tillämpningen av avtalet om frihandel och vissa handelsrelaterade frågor mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Lettland, å andra sidan (21), särskilt artikel 1 i denna,
Artikel 1
- i artikel 1 i kommissionens förordning (EEG) nr 109/80 (24).
- i artikel 6.2 i rådets förordning (EEG) nr 715/90,
- kommissionens förordning (EEG) nr 2699/93 (28),
- kommissionens förordning (EG) nr 1474/95 (31),
6. Artikel 1 i rådets förordning (EEG) nr 2783/75 skall ersättas med följande:
Artikel 2
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 84.2 i detta,
i enlighet med det i artikel 189c i fördraget angivna förfarandet (3), och
Detta utgör en av en serie åtgärder för att förbättra säkerheten till sjöss. ISM-koden har ännu inte tvingande utan endast rekommenderande karaktär.
I sin resolution av den 22 december 1994 om säkerheten på ro-ro-passagerarfartyg (4) uppmanade rådet kommissionen att lägga fram ett förslag om ett påskyndat tvingande genomförande av ISM-koden för alla ro-ro-passagerarfartyg som bedriver reguljär trafik till eller från europeiska hamnar, i överensstämmelse med internationell rätt.
För det tvingande och påskyndade genomförandet av ISM-koden för alla ro-ro-passagerarfartyg, oavsett deras flagg, beaktas även anmodan enligt punkt 2 i IMO:s resolution A.741(18), vilken är en kraftfull uppmaning till regeringarna att införa ISM-koden snarast möjligt, i första hand för passagerarfartyg.
Det är nödvändigt att ange de krav som uppställs för att säkerställa genomförandet av ISM-koden och att definiera villkoren för utfärdande och kontroll av dokumentet om godkänd säkerhetsorganisation och av certifikatet om godkänd säkerhetsorganisation.
Ett förenklat förfarande som omfattar en kommitté med föreskrivande uppgifter är nödvändigt för att ändra denna förordning under beaktande av utvecklingen på internationell nivå.
Artikel 1
- att administrationerna i flagg- och hamnstaterna kontrollerar dessa.
a) ro-ro-passagerarfartyg: ett havsgående passagerarfartyg som är utrustat med anordningar som gör det möjligt för väg- eller järnvägsfordon att rulla på och av fartyget, och som medför fler än 12 passagerare,
2. med resor som företas så regelbundet eller så ofta att de utgör en uppenbar, systematisk serie.
e) ISM-koden: de internationella organisationsreglerna för säker drift av fartyg och för förhindrande av förorening, som antogs av IMO genom församlingens resolution A.741(18) av den 4 november 1993 och som utgör en bilaga till denna förordning,
h) certifikat om godkänd säkerhetsorganisation: det certifikat som i enlighet med punkt 13.4 i ISM-koden utfärdas till ro-ro-passagerarfartyg,
Denna förordning skall tillämpas på alla företag som bedriver reguljär trafik med minst ett ro-ro-passagerarfartyg till eller från en hamn i en medlemsstat inom den Europeiska gemenskapen, oavsett fartygets flagg.
2. Utan hinder av bestämmelserna i punkt 1 får företag som bedriver reguljär trafik med ett eller flera ro-ro-passagerarfartyg enbart i skyddade vatten mellan hamnar som är belägna i en och samma medlemsstat uppskjuta efterlevnaden av bestämmelserna i denna förordning till den 1 juli 1997.
2. För tillämpningen av punkt 1 får medlemsstaterna endast godkänna, eller helt eller delvis förlita sig på, en erkänd organisation.
4. Certifikatet om godkänd säkerhetsorganisation skall endast gälla i fem år från dagen för dess utfärdande, under förutsättning att en mellanliggande kontroll görs åtminstone var trettionde månad eller oftare för att bekräfta att säkerhetsorganisationssystemet fungerar väl och att eventuella ändringar som gjorts sedan den senaste kontrollen överensstämmer med ISM-kodens bestämmelser.
Dokument om godkänd säkerhetsorganisation och certifikat om godkänd säkerhetsorganisation som utfärdats för administrationer i tredje land får endast erkännas om de har utfärdats av en erkänd organisation.
Artikel 7
Artikel 8
För att ta hänsyn till utvecklingen på det internationella planet och särskilt inom IMO får följande ändras, särskilt för att i bilagan införa riktlinjer för administrationer för genomförande av ISM-koden, i enlighet med förfarandet i artikel 10.2:
c) Bilagan.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag från kommissionen. Medlemsstaternas röster skall vägas enligt bestämmelserna i samma artikel. Ordföranden får inte rösta.
c) Om rådet inte har fattat något beslut vid utgången av en period på 40 dagar från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av rådets beslut 93/464/EEG av den 22 juli 1993 om ramprogram för prioriterade åtgärder för statistik information 1993 1997 (3), särskilt artikel 4 a i detta, och med beaktande av följande:
Bland dessa förändringar återfinns de huvudområden där det är möjligt att göra besparingar och där det finns nya eller växande behov. Förändringarna bör vara i överensstämmelse med de överenskomna allmänna principerna.
b) eventuella nödvändiga ändringar i rådets lagstiftning i god tid kan identifieras, förberedas och föreslås av kommissionen samt dessutom att kommissionen kan anta genomförandebestämmelser till rådets lagstiftning i god tid,
e) gemenskapens ekonomiska resurser till stöd för detta program utnyttjas så effektivt som möjligt som ett komplement till andra nationella resurser.
För att uppnå önskade besparingar kan det bli nödvändigt med anpassningar av det tekniska genomförandet av vissa undersökningar. Innan dessa anpassningar beviljas bör de undergå lämpliga säkerhetskontroller.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
För att jordbruksstatistiken bättre skall tillfredsställa det informationsbehov som reformen av den gemensamma jordbrukspolitiken leder till, skall medlemsstaterna, inom ramen för tillgängliga resurser, vidta lämpliga åtgärder för att anpassa sina nationella system för jordbruksstatistik. Medlemsstaterna skall härvidlag beakta de arbetsområden som anges i bilagorna I och II till detta beslut samt de mål, variabler och kriterier som anges i bilaga III.
Kommissionen skall i samråd med medlemsstaterna
c) fastställa och genomföra åtgärder på gemenskapsnivå som är betydelsefulla för syftet med detta beslut.
Den anpassningsprocess för gemenskapens jordbruksstatistik som avses i artikel 1 skall samordnas av kommissionen med hjälp av tekniska handlingsplaner i enlighet med vad som anges i artikel 4. Efter denna period kan rådet besluta om en förlängning i enlighet med kommissionens förslag i artikel 11.
1. Kommissionen skall varje år fastställa en teknisk handlingsplan för jordbruksstatistiken i enlighet med förfarandet i artikel 10. Dessa planer skall omfatta de åtgärder som medlemsstaterna skall genomföra i enlighet med artikel 1. Disponibla resurser skall användas på ett sådant sätt att största möjliga förbättring av den gemensamma jordbruksstatistikens kostnadseffektivitet sker när kraven från gemenskapslagstiftningen, de informella avtalen och de nya informationsbehoven skall uppfyllas.
b) Skriftlig information som medlemsstaterna skall lämna enligt artikel 5 b och 5 c.
Medlemsstaternas rapporter
b) en kortfattad beskrivning av de åtgärder som anges i planen för det kommande året (år n + 1),
I enlighet med det förfarande som anges i artikel 10 kommer kommissionen att utarbeta förenklade modeller för att underlätta utarbetandet av dessa rapporter.
1. Kommissionen skall bidra till medlemsstaternas kostnader för att anpassa sina nationella system för jordbruksstatistik eller till kostnaderna för de förberedande arbeten som hänger samman med nya eller växande behov och som utgör en del av en teknisk handlingsplan.
Artikel 7
Artikel 8
Artikel 9
a) Medlemsstaternas rapporter om genomförandet av åtgärderna under det föregående året.
d) Gemenskapens finansiella bidrag enligt artikel 6.
Nödvändiga åtgärder för tillämpningen
Kommissionen skall själv anta de föreslagna åtgärderna om de är förenliga med kommitténs yttrande.
Artikel 11
Artikel 12
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
I artikel 10 till 18 i direktiv 90/220/EEG fastställs ett gemenskapsförfarande som bemyndigar en medlemsstats behöriga myndighet att medge utsläppande på marknaden av levande produkter som består av genetiskt modifierade organismer.
Enligt artikel 13.3 skall kommissionen därför besluta enligt förfarandet i artikel 21 i direktiv 90/220/EEG.
- Tillstånd till utsläppande på marknaden av denna produkt bör inte omfatta dess användning som livsmedel eller djurfoder, eftersom den anmälan som ingått omfattar dessa aspekter.
Tillstånd för användning av kemiska herbicider på växter, samt utvärderingen av deras inverkan på människors hälsa och på miljön är underkastade rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande på marknaden av växtskyddsprodukter (3), senast ändrat genom kommissionens direktiv 96/12/EG (4), och faller därför inte under tillämpningsområdet för direktiv 90/220/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Produkten består av frön och plantor från cikorialinjerna Cichorium intybus L. subspecies radicchio rosso (RM3-3, RM3-4 och RM3-6) som framställts med hjälp av Agrobacterium tumefaciens-modifierad Ti-plasmid och som innehåller följande inom T-DNA-gränserna:
iii) Neo-genen från Escherichia coli (neomycinfosfotransferas II) med promotorn från nopalinsyntasgenen från Agrobacterium tumefaciens och octopinsyntasgenterminatorn från Agrobacterium tumefaciens.
4. Utan att det påverkar bestämmelserna om etikettering och märkning i övrig gemenskapslagstiftning skall det på etiketten till varje utsädesförpackning anges att produkten
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
En expertdelegation utsänd av kommissionen har kommit tillbaka från Mauretanien efter att ha förvissat sig om villkoren för produktion, lagring och transport av fiskeriprodukter med gemenskapen som destination.
Villkoren för det intyg som avses i artikel 11.4 a i direktiv 91/493/EEG omfattar fastställande av en mall för intyget, vilket eller vilka språk intyget skall vara avfattat på och vilken ställning den som undertecknar intyget skall ha.
MPEM - CNROP - DVIS har officiellt gett försäkringar i fråga om efterlevnaden av de regler som anges i kapitel V i bilagan till direktiv 91/493/EEG och i fråga om krav som är likvärdiga med dem som föreskrivs i det direktivet för godkännande av anläggningar och frysfartyg.
1. Det intyg som avses i artikel 2.1 skall utfärdas på minst ett av de officiella språken i den medlemsstat där kontrollen äger rum.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Föreskrifterna i Elfenbenskustens lagstiftning i fråga om inspektion och hygienkontroll av fiskeriprodukter kan betraktas som likvärdiga med dem som fastställs genom direktiv 91/493/EEG.
Det är lämpligt att i enlighet med artikel 11.4 b i direktiv 91/493/EEG anbringa ett märke med uppgifter om det tredje landets namn och ursprungsanläggningens godkännandenummer på förpackningen för fiskeriprodukterna.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
2. I intyget skall finnas namn och tjänstebeteckning på representanten för MARA-DGRA, dennes namnteckning samt den officiella stämpeln för MARA-DGRA; allt detta skall vara i en annan färg än övriga uppgifter i intyget.
RÅDETS DIREKTIV 96/22/EG av den 29 april 1996 om förbud mot användning av vissa ämnen med hormonell och tyreostatisk verkan samt av â-agonister vid animalieproduktion och om upphävande av direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG
med beaktande av kommissionens förslag (1),
med beaktande av följande: 1. Genom rådets direktiv 81/602/EEG (4) förbjöds vissa ämnen med hormonell eller tyreostatisk verkan och genom direktiv 88/146/EEG (5) förbjöds användningen av vissa ämnen med hormonell verkan i animalieproduktion men tilläts samtidigt vissa undantag.
4. Nya ämnen med anabol verkan såsom â-agonister används illegalt vid uppfödning i syfte att stimulera djurens tillväxt och produktivitet.
7. Tillförsel av läkemedel baserade på â-agonister kan emellertid tillåtas i noggrant definierade terapeutiska syften för vissa kategorier nötkreatur, hästdjur och sällskapsdjur.
10. Bristande harmonisering på gemenskapsnivå beträffande karenstid och de stora skillnader som föreligger mellan medlemsstater, särskilt beträffande godkända veterinärmedicinska läkemedel som innehåller hormonella substanser eller â-agonister, gör att maximala karenstider för dessa läkemedel i harmoniseringssyfte bör bestämmas.
13. Effektiv kontroll av tillämpningen av bestämmelserna i detta direktiv bör säkerställas.
16. Den 18 januari 1996 uppmanades kommissionen och rådet av Europaparlamentet att fortsätta att motsätta sig import av hormonbehandlat kött till gemenskapen; parlamentet önskade att totalförbudet mot användning av tillväxtbefrämjande medel i uppfödningen skulle kvarstå och uppmanade i detta syfte rådet att snarast anta kommissionens förslag om vilket parlamentet yttrat sig den 19 april 1994.
1. I detta direktiv tillämpas de definitioner för kött och köttprodukter som återfinns i direktiv 64/433/EEG (7), 71/118/EEG (8), 77/99/EEG (9), 91/495/EEG (10) för vattenbruksprodukter som återfinns i direktiv 91/493/EEG (11), samt de definitioner för veterinärmedicinska läkemedel som återfinns i direktiv 81/851/EEG (12) och 81/852/EEG (13).
b) terapeutisk behandling: tillförsel av godkända ämnen genom tillämpning av artikel 4 i det här direktivet, till ett enstaka husdjur i syfte att, efter undersökning av en veterinär, behandla fertilitetsstörningar inklusive avbrytande av oönskad dräktighet och när det gäller â-agonister, för att motverka livmoderkontraktioner hos kor vid kalvning samt behandla andningssvårigheter och motverka livmoderkontraktioner hos hästdjur som uppfötts av andra skäl än för köttproduktion,
ii) till vattenbruksdjur, till en avelsgrupp i syfte att erhålla inverterat kön, efter förskrivning av veterinär och på dennes ansvar,
Medlemsstaterna skall säkerställa att följande förbjuds:
c) Avyttring av vattenbruksdjur, som livsmedel, om djuren tillförts ämnen som avses i a, samt bearbetade produkter av dessa djur.
Artikel 4
- slag av behandling,
- behandlade djurs identititet.
i) trenbolon allyl som skall intas oralt eller â-agonister till hästdjur eller sällskapsdjur under förutsättning att de används enligt tillverkarens specifikationer,
Innehav av veterinärmedicinska läkemedel som innehåller â-agonister vilka kan användas för att motverka livmoderkontraktioner är förbjuden.
Trots artikel 3 a och utan att det påverkar tillämpningen av artikel 2, kan medlemsstaterna i zootekniskt syfte tillåta tillförsel till husdjur av veterinärmedicinska läkemedel med östrogen, androgen eller gestagen verkan, godkända enligt direktiv 81/851/EEG och 81/852/EEG. Tillförseln skall utföras av en veterinär till noggrant identifierade djur och behandlingen skall registreras av den ansvarige veterinären enligt artikel 4.1.
I de fall som avses i denna artikel, skall veterinären utfärda ett recept som inte kan förnyas, i vilket den aktuella behandlingen skall specificeras och nödvändig mängd av produkten anges, och veterinären skall också registrera förskrivna produkter.
1. Hormonprodukter och â-agonister vars tillförsel till husdjur enligt artikel 4 och 5 är tillåten, skall motsvara kraven i direktiv 81/851/EEG och 81/852/EEG.
i) Produkter med depåeffekt.
- som är godkända enligt de bestämmelser som var i kraft före ändringen genom förordning (EEG) nr 2309/93 (14),
b) Veterinärmedicinska läkemedel som innehåller â-agonister med en karenstid som överstiger 28 dygn efter avslutad behandling.
Handel med hästar med högt värde, särskilt kapplöpningshästar, tävlingshästar, cirkushästar eller hästar avsedda för betäckning eller utställning, inklusive registrerade hästdjur som tillförts veterinärmedicinska läkemedel innehållande trenbolon allyl eller â-agonister i de syften som anges i artikel 4, kan emellertid äga rum innan karenstiden är över, under förutsättning att villkoren för tillförsel har uppfyllts och att slag av behandling samt datum för behandling anges på det intyg eller pass som följer med dessa djur.
Medlemsstaterna skall säkerställa följande:
a) om förbjudna ämnen eller produkter som är avsedda för tillförsel till djur i tillväxtbefrämjande syfte enligt artikel 2 innehas eller förekommer,
d) om restriktionerna i artikel 4 och 5 för användning av vissa substanser eller produkter respekteras.
4) Att när kontrollerna enligt punkt 2 och 3
Artikel 9
Artikel 10
1. Tredje länder vilkas lagstiftning tillåter avyttring och tillförsel av stilbener, stilbenderivat, deras salter eller estrar samt tyreostatiska medel i syfte att tillföra dem till alla djurarter, får inte finnas på någon lista som enligt gemenskapslagstiftningen reglerar från vilka länder medlemsländerna har tillstånd att importera husdjur eller vattenbruksdjur eller kött eller produkter från sådana djur.
i) som på något sätt tillförts produkter eller ämnen som avses i artikel 2 a,
3. Djur avsedda för avel, uttjänta avelsdjur, eller deras kött, vilka härrör från tredje land, får emellertid importeras under förutsättning att de uppfyller garantier som minst motsvarar dem som anges i detta direktiv och som inrättats enligt förfarandet i artikel 33 i rådets direktiv 96/23/EG, och med tillämpning av kapitel V i det direktivet.
Rådet får, på förslag av kommissionen och med kvalificerad majoritet, anta nödvändiga övergångsåtgärder innan den ordning som föreskrivs i detta direktiv trätt i kraft.
2. Hänvisningar till de upphävda direktiven skall läsas som hänvisningar till detta direktiv och skall läsas enligt jämförelsetabellen i bilagan.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter för hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 15
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100a i detta,
I direktiv 76/116/EEG fastställs bestämmelser för saluföring av gödselmedel på den inre marknaden.
Åtgärderna i detta direktiv är förenliga med yttrandet från Kommittén för anpassning till teknisk utveckling av direktiven om avskaffandet av tekniska hinder för handel med gödselmedel.
Bilaga I till direktiv 76/116/EEG ändras på följande sätt:
>Plats för tabell>
2. Medlemsstaterna skall underrätta kommissionen om de nationella bestämmelser de antar inom det område som omfattas av detta direktiv.
RÅDETS DIREKTIV 96/42/EG av den 25 juni 1996 om ändring av direktiv 77/388/EEG om ett gemensamt system för mervärdeskatt
med beaktande av kommissionens förslag,
med beaktande av följande: I artikel 12.3 d i direktiv 77/388/EEG (3), anges att de regler som gäller beskattningen av andra jordbruksprodukter än dem som tillhör kategori 1 i bilaga H enhälligt skall antas av rådet på kommissionens förslag senast den 31 december 1994. Till och med denna dag tilläts de medlemsstater som redan tillämpade en reducerad skattesats behålla denna medan de som tillämpade normalskattesatsen inte fick använda en reducerad skattesats. Denna bestämmelse tillät en senareläggning av tillämpningen av normalskattesatsen med två år.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 12.3 skall punkt d utgå.
Artikel 2
Detta direktiv gäller från och med den 1 januari 1995.
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 96/57/EG av den 3 september 1996 om energieffektivitetskrav för elektriska kylskåp och frysar (även i kombination) för hushållsbruk
med beaktande av kommissionens förslag (1),
med beaktande av följande: 1. Det är viktig att främja åtgärder som syftar till att den inre marknaden fungerar väl.
4. Några medlemsstater står i begrepp att anta bestämmelser om energieffektiviteten hos kylskåp och frysar för hushållsbruk, vilka bestämmelser är av sådant slag att de kan medföra handelshinder för dessa produkter inom gemenskapen.
7. I artikel 130r i fördraget föreskrivs dessutom att gemenskapens miljöpolitik skall bidra till bland annat målen att skydda och förbättra miljön samt att utnyttja naturresurserna varsamt och rationellt. Produktion och förbrukning av elektricitet bidrar till ungefär 30 % av koldioxidutsläpp (CO2) förorsakade av människor och motsvarar ungefär 35 % av gemenskapens bruttoenergiförbrukning och denna andel ökar.
10. Genom rådets beslut 91/565/EEG (6) upprättades ett program för att främja effektiv energianvänding i gemenskapen (Save-programmet).
13. Direktiv 92/75/EEG (7) (ramdirektivet) och kommissionens direktiv 94/2/EG (8) (om genomförandet av direktiv 92/75/EEG) som föreskriver obligatorisk märkning av apparater och andra former av upplysningar om energiförbrukning kommer att öka konsumenternas medvetenhet om energieffektivitet hos kylskåp och frysar för hushållsbruk. Denna åtgärd kommer följaktligen även att leda till att de konkurrerande tillverkarna erbjuder apparater med högre energieffektivitet än vad som föreskrivs i direktivets normer. I konsumentupplysningarna bör normerna ändå anges för att de ska bli så effektiva som möjligt och leda till en verklig förbättring av de sålda apparaternas genomsnittliga samlade effektivitet.
16. Hänsyn bör tas till beslut 93/465/EEG av den 22 juli 1993 om moduler för olika stadier i förfaranden vid bedömning av överensstämmelse samt regler inför anbringande och användning av CE-märkning om överensstämmelse, avsedda att användas i tekniska harmoniseringsdirektiv (10).
19. Detta direktiv omfattar inte kylskåp och frysar som tillverkats enligt särskilda specifikationer utan endast nätanslutna kylskåp och frysar för hushållsbruk, avsedda för livsmedel. Kyl- och frysanläggningar för kommersiellt bruk är avsevärt mer varierade och kan därför inte omfattas av detta direktiv.
Detta direktiv skall tillämpas på nya nätanslutna kylskåp, frysfack och frysar, även i kombination, för hushållsbruk, enligt bilaga I, nedan kallade "kyl- och frysapparater". Apparater som även kan utnyttja andra energikällor, t.ex. batterier, samt kyl- och frysapparater för hushållsbruk som bygger på absorptionsprincipen och apparater som tillverkats enligt särskilda specifikationer omfattas inte av direktivet.
2. Tillverkaren av en kyl- och frysapparat som omfattas av detta direktiv, dennes i gemenskapen etablerade ombud eller den person som ansvarar för att apparaten släpps ut på marknaden inom gemenskapen åläggs att se till att varje apparat som släppts ut på marknaden uppfyller kravet som avses i punkt 1.
2. Om det inte finns bevis om motsatsen skall medlemsstaterna utgå från att kyl- och frysapparater med EG-märkning enligt artikel 5 överensstämmer med samtliga bestämmelser i detta direktiv.
Artikel 4
1. Apparaterna skall, då de släpps ut på marknaden, vara försedda med EG-märkning. Denna skall bestå av bokstäverna "CE". Den utformning som skall användas visas i bilaga III. EG-märkningen skall vara väl synlig, läsbar och outplånligt anbringad på kyl- och frysapparaterna samt vid behov på emballaget.
1. Om en medlemsstat konstaterar att EG-märkningen har använts på ett oriktigt sätt är tillverkaren eller dennes i gemenskapen etablerade ombud skyldig att anpassa produkten till bestämmelserna och upphöra med överträdelsen på de villkor som medlemsstaten föreskriver. Om varken tillverkaren eller dennes ombud är etablerade i gemenskapen åligger denna skyldighet den person som ansvarar för att kyl- och frysapparaten släpps ut på marknaden i gemenskapen.
1. Alla beslut som fattas enligt detta direktiv och som innehåller inskränkningar av villkoren för att släppa ut kyl- och frysapparater på marknaden skall noga ange på vilka grunder beslutet är fattat. Den berörda parten skall omedelbart underrättas om beslutet och samtidigt få information om vilka möjligheter till överklagande som gäller i den berörda medlemsstaten och inom vilken tid detta skall äga rum.
Senast fyra år efter det att detta direktiv har antagits skall kommissionen utvärdera de resultat som uppnåtts i förhållande till de förväntade resultaten. Med sikte på att gå vidare med nästa steg i förbättringen av energieffektiviteten skall kommissionen därefter i samråd med de berörda parterna undersöka om det finns behov av att upprätta ytterligare en rad lämpliga åtgärder för att på ett märkbart sätt förbättra energieffektiviteten för kyl- och frysapparater för hushållsbruk. Om så är fallet skall åtgärderna och tidpunkten för deras ikraftträdande grundas på energieffektivitetsnivåer som är ekonomiskt och tekniskt motiverade med hänsyn till de omständigheter som råder vid det tillfället. Andra åtgärder som har bedömts vara lämpliga för att förbättra effektiviteten för kyl- och frysapparater för hushållsbruk kommer också att beaktas.
Medlemsstaterna skall tillämpa sådana bestämmelser tre år efter antagandet av detta direktiv.
3. Under en tid av tre år efter antagandet av detta direktiv skall medlemsstaterna tillåta att sådana kyl- och frysapparater släpps ut på marknaden som är godkända i respektive medlemsstat vid den tidpunkt detta direktiv antas.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
Bromsprovningstestet kan förbättras genom att medelretardationen ersätts med en formel som anger bromssträckan som en funktion av hastigheten. Denna ändring kommer att följas av ytterligare ändringar i syfte att öka säkerheten för traktorer och de element som berör deras användning.
Artikel 1
1. Från och med den 1 oktober 1997 får medlemsstaterna inte
- inte längre bevilja EG-typgodkännande eller ett sådant dokument som avses i artikel 10.1 sista strecksatsen i direktiv 74/150/EEG, och
Artikel 3
3. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
Europaparlamentets och rådets direktiv 96/74/EG av den 16 december 1996 om benämningar på textilier (5) föreskriver obligatorisk märkning för att ange vilka fibrer som ingår i textilvaror. Att märkningarna överensstämmer med innehållet i varorna kontrolleras genom analyser.
Den tekniska utvecklingen gör det nödvändigt att med täta mellanrum anpassa de tekniska specifikationer som definieras i särdirektiven om metoder för analys av textilier. För att underlätta genomförandet av de åtgärder som krävs för detta bör ett förfarande fastställas som upprättar ett nära samarbete mellan medlemsstaterna och kommissionen, i Kommittén för direktiv om benämningen och märkningen av textilier.
Detta direktiv skall inte påverka medlemsstaternas skyldigheter att överföra direktiven inom de tidsfrister som anges i bilaga III del B.
Detta direktiv gäller metoder för kvantitativ analys av vissa binära textilfiberblandningar, inklusive framtagning av analysprov och provexemplar.
Provexemplar avser den del av analysprovet som behövs för ett enskilt provningsresultat.
Artikel 4
1. Härmed inrättas en kommitté för direktiv om benämningen och märkningen av textilier (nedan kallad "kommittén"). Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
Artikel 6
3. a) Kommissionen skall anta de föreslagna åtgärderna om det är förenligt med kommitténs yttrande.
c) Om rådet inte har fattat något beslut inom tre månader från det att förslaget har mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 8
Artikel 9
RÅDETS DIREKTIV 96/75/EG av den 19 november 1996 om system för befraktning och prissättning inom området nationella och internationella transporter av varor på inre vattenvägar inom gemenskapen
med beaktande av kommissionens förslag (1),
med beaktande av följande: De tilltagande problem som rör överbelastning av vägtrafikleder och järnvägslinjer, transportsäkerheten, miljön, energisparande och medborgarnas livskvalitet kräver i allmänhetens intresse en längre driven utveckling och ett bättre utnyttjande av transportmöjligheterna på inre vattenvägar, genom bland annat förbättrad konkurrenskraft för dessa transporter.
För detta ändamål bör en övergångsperiod föreskrivas med en successiv begränsning av tillämpningsområdet för systemet med befraktning i turordning för att transportörerna skall kunna anpassa sig till den fria marknadens villkor och i förekommande fall genomföra former för kommersiella sammanslutningar som är bättre anpassade till avlastarnas logistiska behov.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) system med befraktning i turordning: ett system som består i att transportförfrågningar från kundkretsen fördelas i en befraktningspool till fastställda priser och enligt offentliggjorda villkor, i den ordning som fartygen blir tillgängliga efter lossning. Transportörerna erbjuds, i den ordning de anmält sig till turordningen, att välja ut en transport bland dem som bjuds ut. De som inte väljer behåller likväl sin plats i turordningen,
d) allvarlig marknadsstörning: uppträdande på marknaden för varutransport på inre vattenvägar av specifika problem av ett slag som kan medföra ett allvarligt och eventuellt bestående överskott av utbud i förhållande till efterfrågan och som innebär ett allvarligt hot mot den ekonomiska stabiliteten och överlevnaden för ett betydande antal företag som transporterar varor på inre vattenvägar, under förutsättning att de kort- och medellångsiktiga prognoserna på den aktuella marknaden inte visar betydande och varaktiga förbättringar.
Artikel 3
- att systemen med befraktning i turordning och de fastställda priserna är fritt tillgängliga på samma villkor för alla transportörer i medlemsstaterna.
a) Transporter av olja och gas, flytande och torr last i bulk, specialtransporter av tungt och odelbart gods, containertransporter, transporter inom hamnområden, alla slags transporter för egen räkning samt alla slags transporter som redan utförs utanför systemet med befraktning i turordning.
- kombinerade transporter, det vill säga transporter med flera olika transportmedel där de huvudsakliga sträckorna utgörs av inre vattenvägar och där de inledande och/eller avslutande sträckorna, som skall vara så korta som möjligt, antingen utgör väg eller järnväg.
- föreskriva möjlighet för avlastarna att ingå avtal om flera transporter, det vill säga en serie på varandra följande transporter utförda av ett och samma fartyg,
Inom en frist på två år från och med ikraftträdandet av detta direktiv skall de medlemsstater som berörs av systemen med befraktning i turordning vidta nödvändiga åtgärder för att avlastarna fritt skall kunna välja mellan följande tre slag av avtal:
- Avtal om enstaka eller upprepade transporter.
2. Om en medlemsstat begär lämpliga åtgärder, skall beslut fattas inom tre månader efter det att begäran har mottagits.
- uppgift om i vilken grad lastutrymmet har utnyttjats,
4. De beslut som fattas i enlighet med denna artikel, vilka inte får gälla längre än störningen på marknaden varar, skall medlemsstaterna utan dröjsmål underrättas om.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är, i förekommande fall genom omröstning.
Artikel 9
2. Medlemsstaterna skall genast till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
Det är lämpligt att bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning förfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen (3) ändrad genom Kommissionens förordning (EEG) nr 2454/93 (4), under en period av tre månader.
Artikel 1
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan förfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
KOMMISSIONENS FÖRORDNING (EG) nr 569/96 av den 29 mars 1996 om ändring av förordningarna (EEG) nr 1362/87 och (EEG) nr 1158/91 vad gäller interventionsuppköp och beviljande av stöd för privat lagring av skummjölkspulver och förordning (EEG) nr 1756/93 om avgörande faktorer för den jordbruksomräkningskurs som tillämpas för mjölk och mjölkprodukter
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter (1), senast ändrad genom kommissionens förordning (EG) nr 2931/95 (2), särskilt artiklarna 7.5 och 28 i denna,
I kommissionens förordning (EEG) nr 1362/87 av den 18 maj 1987 om tillämpningsföreskrifter till rådets förordning (EEG) nr 777/87 med avseende på uppköp och beviljandet av stöd för privat lagring av skummjölkspulver (11), senast ändrad genom förordning (EG) nr 1137/94 (12), kommissionens förordning (EEG) nr 1158/91 av den 3 maj 1991 om interventionsorgans uppköp av skummjölkspulver genom anbud (13), senast ändrad genom förordning (EG) nr 1802/95, och kommissionens förordning (EEG) nr 1756/93 (14), senast ändrad genom förordning (EG) nr 315/96 (15), görs det hänvisningar till förordningarna (EEG) nr 1014/68 och (EEG) nr 625/78. I dessa förordningar bör det istället hänvisas till förordning (EG) nr 322/96. Dessutom bör förordning (EEG) nr 1158/91 ändras för att närmare fastställa sättet att beräkna uppköpspriset i förhållande till proteinhalten i skummjölkspulver.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) Punkt a skall ersättas med följande:
3. Artikel 5 skall utgå.
2. I artikel 3 skall punkt 1 ersättas med följande:
- om de skriftligen åtar sig att följa artikel 4.6 i förordning (EG) nr 322/96."
4. Artikel 9 skall ersättas med följande:
Uppköpspriset skall beräknas på följande sätt:
d = anbudspriset × [(0,356 - proteinhalten) × 1,75].
Artikel 3
Artikel 4
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande (1), och
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
För att på ett korrekt sätt kunna bedöma situationen när det gäller socker som köpts eller sålts med stöd av de regler om interventionsåtgärder som fastställts i förordning (EEG) nr 1785/81 måste relevant information finnas, särskilt i fråga om de kvantiteter som hålls av interventionsorganen, samt om fördelningen av dessa kvantiteter på lager som godkänts i enlighet med artikel 1.2 i rådets förordning (EEG) nr 447/68 av den 9 april 1968 om allmänna bestämmelser för interventionsköp av socker (5), senast ändrad genom förordning (EEG) nr 1359/77 (6). För att kunna följa tillämpningen av interventionssystemet är det också viktigt att regelbundet få information om de kvantiteter socker som blivit otjänliga för konsumtion och de kvantiteter som har använts för att tillverka vissa kemiska produkter, varvid också måste anges de kvantiteter socker som antingen har denaturerats i enlighet med någon av de processer som beskrivs i bilagan till kommissionens förordning (EEG) nr 100/72 av den 14 januari 1972 om föreskrifter för denaturering av socker till foderändamål (7), senast ändrad genom förordning (EG) nr 260/96 (8), eller som använts vid tillverkning av de kemiska produkter som räknas upp i bilagan till rådets förordning (EEG) nr 1010/86 av den 25 mars 1986 om allmänna bestämmelser om produktionsbidrag för vissa sockerprodukter som används i den kemiska industrin (9), senast ändrad genom förordning (EG) nr 1101/95, samt de produkter som räknas upp i bilagan till kommissionens förordning (EEG) nr 1729/78 av den 24 juli 1978 om tillämpningsföreskrifter för produktionsbidrag för socker som används i den kemiska industrin (10), senast ändrad genom förordning (EG) nr 260/96.
De personer som berörs skall försäkras om att information som rör enskilda företag omfattas av tystnadsplikt.
Artikel 1
b) de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som tagits över av interventionsorganet,
På begäran av kommissionen skall varje medlemsstat överlämna en förteckning till kommissionen över de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som tagits över av interventionsorganet, samt över fördelningen av dessa kvantiteter på godkända lager.
1. Varje vecka, med avseende på närmast föregående vecka, anmäla de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, för vilka en licens om denatureringsbidrag har utfärdats.
Vad gäller interventionsåtgärder som vidtagits i enlighet med artikel 9.3 i förordning (EEG) nr 1785/81 skall varje medlemsstat till kommissionen anmäla följande:
b) ett produktionsbidrag har utbetalats.
b) ett produktionsbidrag har utbetalats.
Vad gäller export till tredje land skall varje medlemsstat till kommissionen anmäla följande:
- vitsocker KN-nr 1701 91 00, 1701 99 10, 1701 99 90,
- isoglukos uttryckt som torrsubstans KN-nr 1702 40 10, 1702 60 10, 1702 90 30 och 2106 90 30,
c) de kvantiteter C-vitsocker, C-råsocker, C-isoglukos, C-inulinsirap, uttryckta som vitsocker, torrsubstans respektive som socker/isoglukos ekvivalent, för vilka exportlicens har utfärdats,
3. För varje kalendermånad och senast vid utgången av den tredje månaden efter den kalendermånad som anmälan avser:
c) de kvantiteter socker och sackarossirap uttryckt som vitsocker, samt isoglukos uttryckt som torrsubstans, som exporterats obearbetat i enlighet med artikel 2a andra stycket i förordning (EEG) nr 3665/87 med angivande av motsvarande bidrag,
De uppgifter som avses i d och e ovan skall lämnas var för sig till kommissionen i enlighet med de bestämmelser som gäller för respektive bearbetad produkt.
1. Varje vecka, med avseende på närmast föregående vecka, de kvantiteter vitsocker och råsocker angivna i icke omräknad vikt, förutom, förmånssocker, sirap, isoglukos och inulinsirap, för vilka importlicens har utfärdats.
b) importerats från eller exporterats till en annan medlemsstat i obearbetat skick eller i form av bearbetade produkter.
1. Varje vecka, med avseende på närmast föregående vecka, de kvantiteter vitsocker och råsocker angivna i icke omräknad vikt, för vilka import- eller exportlicens utfärdats i enlighet med artikel 10 i förordning (EG) nr 1464/95.
Vad gäller import av förmånssocker åligger följande varje medlemsstat:
a) kopior av relevanta varucertifikat EUR.1,
De dokument som avses i a och b ovan skall förutom de uppgifter som anges i artiklarna 6 och 7 i förordning (EEG) nr 2782/76 innehålla uppgift, med en noggrannhet av sex decimaler, om graden av polarisering av varje importerad kvantitet.
b) den totala kvantiteten råsocker, angiven i ton i icke omräknad vikt,
Artikel 9
2. Senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, anmäla produktionen av isoglukos, fastställd i enlighet med artikel 3.2 och punkt 2a i förordning (EEG) nr 1443/82, vid vart och ett av de isoglukosproducerande företagen på dess territorium. De kvantiteter isoglukos som varje månad producerats inom ramen för bestämmelserna om aktiv förädling skall redovisas separat.
Varje medlemsstat skall varje kalendermånad, med avseende på den närmast föregående kalendermånaden, och allt efter vad som är lämpligt uttryckt som vitsocker, torrsubstans eller som socker/isoglukos ekvivalent, anmäla följande:
Artikel 11
Varje medlemsstat skall till kommissionen anmäla följande:
Emellertid:
Varje medlemsstat skall till kommissionen anmäla följande:
a) de kvantiteter som avses i artikel 4.2 i förordning (EEG) nr 1358/77,
Varje medlemsstat skall till kommissionen anmäla följande:
Artikel 15
I denna förordning avses med
c) närmast föregående produktionsår: referensperioden från och med den 1 oktober ett kalenderår till och med den 30 september påföljande kalenderår.
Om informationen innehåller upplysningar som rör ett enskilt företag, dess tekniska installationer eller arten och omfattningen av dess produktion, eller upplysningar som kunde göra det möjligt att rekonstruera sådana fakta, skall emellertid informationen endast lämnas till de personer som inom kommissionen är ansvariga för marknadsfrågor i sockersektorn. Sådan information får inte lämnas ut till tredje man.
Denna förordning träder i kraft den 1 juli 1996.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Varje medlemsstat anmodas, enligt artikel 5,1 b i förordning (EG) nr 2494/95, att ta fram ett harmoniserat konsumentprisindex (HIKP) där ett första index skall gälla för januari 1997.
Det är nödvändigt att vidta åtgärder för att säkerställa att HIKP blir jämförbara enligt artikel 5.3 i förordning (EG) nr 2494/95.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Målet för denna förordning är att fastställa delindexen till de harmoniserade konsumentprisindexen (HIKP) som varje månad skall beräknas och överlämnas till kommissionen (Eurostat) för vidare spridning.
I denna förordning defineras ett "delindex till HIKP" som ett prisindex för en av de utgiftskategorier som anges i bilaga I och beskrivs i bilaga II till förordningen. De bygger på COICOP/HIKP-klassifikationen (Classification of individual consumption by purpose adopted to the needs of HICPs) (3). "Spridning" avser utlämnande av uppgifter i vilken form som helst.
Medlemsstaterna skall varje månad beräkna och överlämna till kommissionen (Eurostat) alla delindex (bilaga I) som har en vikt som är större än en promille av de totala utgifterna som täcks av HIKP (4). Tillsammans med index för januari 1997 skall medlemsstaterna även till kommissionen (Eurostat) överföra motsvarande uppgifter om vikterna, och därefter vid varje tillfälle som vikterna ändras.
Kommissionen (Eurostat) skall låta sprida delindex av HIKP för de kategorier som anges i bilaga I till denna förordning där index för 1996=100.
Medlemsstaterna skall till kommissionen (Eurostat), på dess begäran, lämna information om fördelningen av varor och tjänster på de olika utgiftskategorierna i bilagorna I och II i tillräcklig omfattning för att kunna utvärdera att förordningen följs.
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Identifieringssystemet kommer regelbundet att ses över och kommer, vid behov, att ändras genom det förfarande som fastställts i artikel 21 i direktiv 94/62/EG.
Artikel 1
I detta beslut skall följande gälla:
Artikel 3
Beslut om att införa ett obligatoriskt identifieringssystem för något av materialen får antas enligt det förfarande som anges i artikel 21 i direktiv 94/62/EG.
KOMMISSIONENS BESLUT av den 12 februari 1997 om precisering av principer för inkomst från institut för kollektiv investering, för tillämpning av rådets direktiv 89/130/EEG, Euratom om harmonisering av beräkningen av bruttonationalinkomst till marknadspris (Text av betydelse för EES) (97/157/EG, Euratom)
med beaktande av Fördraget om upprättandet av Europeiska atomenergigemenskapen,
I nuvarande upplaga av ENS beskrivs inte närmare hur inkomst från institut för kollektiv investering skall bokföras, och detta gäller i synnerhet för ej utdelad inkomst.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Om utdelning sker, skall denna inkomst föras till aktieägarnas inkomstfördelningskonto som kapital- och företagarinkomster (post R40 i gällande ENS).
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Enligt artikel 13.4 i direktiv 89/106/EEG krävs att det förfarande som sålunda bestämts anges i uppdragen och i de tekniska specifikationerna. Det är därför önskvärt att definiera de produkter eller produktgrupper som används i uppdragen och i de tekniska specifikationerna.
Det åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga byggkommittén.
För de produkter och produktgrupper som anges i bilaga I skall överensstämmelsen bestyrkas genom ett förfarande där tillverkaren ensam ansvarar för ett tillverkningskontrollsystem i fabriken som säkerställer att produkten överensstämmer med de relevanta tekniska specifikationerna.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, och
Enda artikel
"Medlemmarna skall utses för en period på tre år."
3. Artikel 9 skall ersättas med följande:
KOMMISSIONENS BESLUT av den 11 december 1997 om upphävande av kommissionens beslut 97/613/EG och om införande av särskilda villkor för import av pistaschmandlar och vissa produkter som är framställda av dessa, som har sitt ursprung i eller försänds från Iran (Text av betydelse för EES) (97/830/EG)
med beaktande av rådets direktiv 93/43/EEG (1) av den 14 juni 1993 om livsmedelshygien, särskilt artikel 10.1 i detta, och med beaktande av följande:
Vetenskapliga livsmedelskommittén har konstaterat att aflatoxin B1, även i mycket små mängder, orsakar levercancer och att ämnet dessutom är genotoxiskt.
Pistaschmandlar och produkter som är framställda av dessa, som har sitt ursprung i eller försänds från Iran får importeras under förutsättning att dessa särskilda villkor uppfylls.
Partier med pistaschmandlar som har sitt ursprung i eller försänds från andra länder utanför EU bör underkastas analyser för att fastställa pistaschmandlarnas halter av aflatoxin B1 och den totala aflatoxinhalten, oberoende av varifrån pistaschmandlarna kommer. De samordnade programmen för officiell kontroll av livsmedel bör därför kompletteras.
Artikel 1
1. Medlemsstaterna får importera
som har sitt ursprung i eller som försänds från Iran, under förutsättning att sändningen åtföljs av officiella provtagnings- och analysresultat samt av ett hälsointyg enligt bilaga I, ifyllt, undertecknat och kontrollerat av en företrädare för det iranska hälsoministeriet.
4. De behöriga myndigheter i varje medlemsstat skall säkerställa att importerade pistaschmandlar som har sitt ursprung i, eller sänds från Iran, underkastas dokumentkontroller i syfte att säkerställa att sändningarna överensstämmer med de krav för hälsointyg och provtagningsresultat som avses i punkt 1.
Detta beslut skall tas upp till förnyad behandling senast den 31 oktober 1998, för att bedöma huruvida de särskilda villkor som avses i artikel 2 ger ett tillräckligt skydd av folkhälsan i gemenskapen. Vid översynen skall också fastställas om det finns fortsatt behov av de särskilda villkoren.
Artikel 5
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av följande: Textilprodukter får endast införas på gemenskapsmarknaden om de uppfyller direktivets bestämmelser.
Detta direktivs bestämmelser är i enlighet med det yttrande som Kommittén för direktiv om benämningen och märkningen av textilier har avgett.
Bilaga I till direktiv 96/74/EG ändras på följande sätt:
- I kolumnen "beskrivning" läggs "kashgoraget" (en korsning mellan kashmirget och angoraget) till efter "guanaco".
3) Numren 31-41 ersätts med 34-44.
5) Ett nytt nr 32 införs enligt följande:
"fiber av regenererad cellulosa som fås genom upplösning och en spinnprocess i organiskt lösningsmedel utan att derivats bildas".
"fiber av regenererad cellulosa som erhålls genom en ändrad viskosprocess och som har en hög hållfasthet och en hög våtmodul. Hållfastheten (BC) i konditionerat provningstillstånd och den dragkraft (BM) som krävs för att åstadkomma en förlängning om 5 % i vått tillstånd är följande:
1) Numren 31-41 ersätts med 34-44.
>Plats för tabell>
>Plats för tabell>
>Plats för tabell>
De skall genast underrätta kommissionen om detta.
Artikel 4
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
2. Genom direktiven 92/50/EEG (5), 93/36/EEG (6) och 93/37/EEG (7) samordnades de nationella förfarandena vid tilldelning av offentliga tjänstekontrakt, varukontrakt respektive bygg- och anläggningskontrakt för att införa rättvisa konkurrensvillkor för sådana kontrakt i alla medlemsstater.
5. Vissa av avtalets bestämmelser medför fördelaktigare villkor för anbudsgivande företag än de som framgår av direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG.
8. Tillämpningen av dessa direktiv måste förenklas samtidigt som jämvikten i gemenskapens gällande lagstiftning om offentlig upphandling måste bibehållas så långt det är möjligt.
11. Kommissionen bör tillhandahålla små och medelstora företag utbildnings- och informationsunderlag för att göra det möjligt för dem att fullt ut delta i det ändrade upphandlingsförfarandet.
A) ersätts punkterna 1 och 2 med följande text:
- de offentliga kontrakt avseende sådana tjänster som avses i bilaga I A, med undantag för tjänster i kategori 8 och telekommunikationstjänster i kategori 5, med CPD-referensnumren 7524, 7525 och 7526,
b) Motvärdena i ecu och nationella valutor för de tröskelvärden som fastställs i a skall i princip revideras vartannat år med verkan från den 1 januari 1996. Beräkningen av detta motvärde skall grundas på den genomsnittliga dagskursen för dessa valutor uttryck i ecu och för ecun uttryckt i SDR under de sista 24 månaderna fram till den sista augusti som föregår revisionen per den 1 januari.
2. Vid beräkning av det uppskattade värdet av ett kontrakt skall den upphandlande myndigheten inkludera den uppskattade, sammanlagda ersättningen till tjänsteleverantören med beaktande av bestämmelserna i punkterna 3 7."
"1. Den upphandlande myndigheten skall inom 15 dagar efter att ha mottagit en skriftlig begäran underrätta varje anbudssökande eller anbudsgivare vars ansökan eller anbud har förkastats om orsakerna till att hans ansökan eller anbud förkastats samt underrätta varje anbudsgivare som lämnat ett godtagbart anbud om utformningen av och de relativa fördelarna med det antagna anbudet samt namnet på den anbudsgivare som tilldelats kontraktet.
3. Artikel 13.1 och 13.2 ersätts med följande text:
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen i för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG, eller
- det tröskelvärde som avses i artikel 7.1 a första strecksatsen för de tjänster som avses i bilaga I B, tjänsterna i kategori 8 i bilaga I A och telekommunikationstjänsterna i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, eller
4. Artikel 18.2 ersätts med följande text:
"4. Tidsfristen för mottagande av anbud enligt punkt 3 får förkortas till 26 dagar om de upphandlande myndigheterna har avsänt det preliminära förhandsmeddelande som avses i artikel 15.1, utformat enligt förlagan i bilaga III A (förhandsinformation), till Europeiska gemenskapernas officiella tidning minst 52 dagar och högst tolv månader före dagen för insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 15.2, och om det preliminära förhandsmeddelandet dessutom innehåller minst den information som föreskrivs i förlagan i bilaga III C (selektivt förfarande) eller, beroende på omständigheterna, i bilaga III D (förhandlat förfarande,) förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
- att varje anbud innehåller de upplysningar som krävs för att utvärdera det,
- att öppnande av anbuden äger rum efter utgången av den tidsfrist som bestäms för avgivande av dessa."
1. För att möjliggöra bedömning av resultatet av tillämpningen av det här direktivet skall medlemsstaterna till kommissionen sända en statistisk rapport rörande de tjänstekontrakt som under föregående år tilldelats av de upphandlande myndigheterna, senast den 31 oktober 1997 och därefter senast den 31 oktober varje år.
- det uppskattade sammanlagda värdet för kontrakt som av varje upphandlande myndighet tilldelas under tröskelvärdet,
c) När det gäller de upphandlande myndigheter som framgår av bilaga I till direktiv 93/36/EEG, antal och sammanlagt värde för kontrakt som tilldelas av varje upphandlande myndighet enligt undantagen från avtalet. När det gäller övriga upphandlande myndigheter som omfattas av detta direktiv, det sammanlagda värdet för kontrakt som tilldelats av varje upphandlande myndighet enligt undantagen från avtalet.
3. Kommissionen skall enligt det förfarande som anges i artikel 40.3 bestämma arten av de statistiska upplysningar som krävs enligt det här direktivet."
Direktiv 93/36/EEG ändras på följande sätt:
"1. a) Avdelningarna II, III och IV samt artiklarna 6 och 7 skall gälla offentliga varukontrakt som tilldelas av
b) Det här direktivet gäller offentlig upphandling av varor vilkas uppskattade värde är lika med eller högre än det tröskelvärde som gäller vid tidpunkten för offentliggörande av meddelandet enligt artikel 9.2.
d) De tröskelvärden som avses i a och deras motvärden uttryckta i ecu och nationella valutor skall regelbundet offentliggöras i Europeiska gemenskapernas officiella tidning i början av november efter den revision som avses i c första stycket."
2. Artikel 7.1 och 7.2 ersätts med följande text:
2. De upphandlande myndigheterna skall så snart som möjligt underrätta de anbudssökande och anbudsgivarna om de beslut som fattas rörande tilldelningen av kontrakt, inklusive skälen till att de har beslutat att avstå från en upphandling för vilken anbud begärts eller att upprepa förfarandet; dessa upplysningar skall på begäran lämnas skriftligen. Myndigheterna skall även underrätta Byrån för Europeiska gemenskapernas officiella publikationer om dessa beslut."
4. I artikel 11 skall följande punkt föras in:
"3. Anbud skall avges skriftligen, direkt eller per post. Medlemsstaterna får tillåta avgivande av anbud på alla andra sätt som gör det möjligt att säkerställa
- om det är nödvändigt av bevisskäl, att anbud så snart som möjligt bekräftas skriftligen eller genom översändande av en bestyrkt kopia,
2. Kommissionen skall se över detta direktiv och varje ny åtgärd som kan ha tillkommit enligt vad som sägs i punkt 1, med hänsyn till resultaten av de nya förhandlingar som avses i artikel XXIV.7 i avtalet om offentlig upphandling, som ingåtts inom ramen för de multilaterala förhandlingarna i Uruguayrundan (*), nedan kallat "avtalet`, och den skall i förekommande fall lägga fram lämpliga förslag för rådet.
2. Den statistiska rapporten skall innehålla åtminstone följande:
- antal och värden för kontrakt som av varje upphandlande myndighet tilldelas över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, varukategori i enlighet med den terminologi som avses i artikel 9.1 och nationalitet för den varuleverantör som tilldelas kontraktet samt, i fråga om förhandlade förfaranden, med uppdelning enligt artikel 6 med uppgift om antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
d) Alla andra statistiska upplysningar som skall bestämmas i enlighet med förfarandet i artikel 32.2 och som begärs i enlighet med avtalet.
Artikel 3
A) ersätts punkterna 1 och 2 med följande text:
b) offentliga bygg- och anläggningsarbeten som avses i artikel 2.1 när det uppskattade värdet exklusive mervärdesskatt uppgår till minst 5 000 000 ecu.
b) Den beräkningsmetod som anges under a skall på förslag av kommissionen ses över av Rådgivande kommittén för offentlig upphandling i princip två år efter dess första tillämpning."
2. Artikel 8.1 och 8.2 ersätts med följande text:
2. De upphandlande myndigheterna skall så snart som möjligt underrätta de anbudssökande och anbudsgivarna om de beslut som fattats rörande tilldelningen av kontrakt, inklusive skälen till att de har beslutat att avstå från en upphandling för vilken anbud begärts eller att upprepa förfarandet; dessa upplysningar skall på begäran lämnas skriftligen. Myndigheterna skall även underrätta Byrån för Europeiska gemenskapernas officiella publikationer om dessa beslut."
4. Artikel 13.4 ersätts med följande text:
"2. Anbud skall avges skriftligen, direkt eller per post. Medlemsstaterna får tillåta avgivande av anbud på alla andra sätt som gör det möjligt att säkerställa
- om det är nödvändigt av bevisskäl, att anbud så snart som möjligt bekräftas skriftligen eller genom översändande av en bestyrkt kopia,
"Artikel 33a
a) När det gäller de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG
b) När det gäller de upphandlande myndigheter som omfattas av detta direktiv antal och värde för kontrakt som tilldelats av varje kategori av upphandlande myndigheter över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, kategori av bygg- och anläggningsarbeten i enlighet med den terminologi som används i bilaga II och nationaliteten för det företag som tilldelats kontraktet samt, i fråga om förhandlande förfaranden, med uppdelning enligt artikel 7 med uppgift om antal och värden för de kontrakt som tilldelats varje medlemsstat och tredje land.
3. Kommissionen skall enligt det förfarande som föreskrivs i artikel 35.3 bestämma arten av de statistiska upplysningar som krävs enligt detta direktiv."
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 13 oktober 1998. De skall genast underrätta kommissionen om detta.
Artikel 5
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
Kommissionen har behov av relevanta uppgifter om vissa ämnen för att kunna inleda de förfaranden för översyn som avses i artiklarna 69, 84 och 112 i anslutningsfördraget för bestämmelser som ännu inte tillämpas i de nya medlemsstaterna. Dessa upplysningar måste finnas tillgängliga innan alla de upplysningar som avses i artiklarna 3 och 4 i förordning (EEG) nr 793/93 finns att tillgå.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som inrättats i enlighet med artikel 15 i förordning (EEG) nr 793/93.
De som tillverkar eller importerar ämnen som ingår i förteckningen i bilagan till denna förordning skall inom fyra månader efter det att förordningen träder i kraft till kommissionen lämna all relevant tillgänglig information om exponering av människor eller miljö för dessa ämnen.
- delar av miljön omfattar vatten, mark och luft, vilket också innefattar information om ämnets fördelning och omvandling i reningsverk och dess ackumulering i näringskedjan och
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av kommissionens förslag (3),
med beaktande av följande: Enligt förordning (EG) nr 3281/94 och förordning (EG) nr 1256/96 omfattas Unionen Myanmar (nedan kallad Myanmar) av allmänna tullförmåner.
Den 2 januari 1997 anmälde ICFTU och ETUC till kommissionen att de utvidgade omfattningen av det gemensamma klagomål som de ingivit enligt förordning (EG) nr 3281/94 i syfte att det tillfälliga upphävandet av gemenskapens system med förmåner för Myanmar även görs enligt förordning (EG) nr 1256/96.
De skriftliga och muntliga uppgifter som kommissionen har inhämtat i samband med undersökningen som genomfördes i samråd med kommittén för förvaltningen av allmänna tullförmåner stödjer de påståenden som anges i klagomålet. Det framgår att myndigheterna i Myanmar rutinmässigt med tillgripande av tvång och upprepade våldsamma straffåtgärder har tillämpat tvångsarbete inte endast för militära operationer utan även för civila och militära infrastrukturbyggprojekt.
Av de tillgängliga uppgifterna framgår alltså att det finns tillräckliga skäl att dra slutsatsen att ett upphävande av systemet med allmänna tullförmåner som har beviljats Myanmar är berättigat.
Mot bakgrund av detta bör tillämpningen av allmänna tullförmåner för industriprodukter och jordbruksprodukter med ursprung i Myanmar tillfälligt upphävas till dess det fastställts att metoderna i fråga har upphört.
Artikel 1
Rådet skall, med kvalificerad majoritet, på förslag av kommissionen, låta upphäva tillämpningen av denna förordning då det på grundval av en rapport om tvångsarbete i Myanmar från kommissionen kan visas att de metoder som avses i artikel 9.1 första strecksatsen i förordning (EG) nr 3281/94 och artikel 9.1 första strecksatsen i förordning (EG) nr 1256/96 som har orsakat upphävandet av allmänna tullförmåner för Myanmar inte längre förekommer.
KOMMISSIONENS FÖRORDNING (EG) nr 659/97 av den 16 april 1997 om tillämpningsföreskrifter för förordning (EG) nr 2200/96 med avseende på interventionsordningen för frukt och grönsaker
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker (1), särskilt artiklarna 30.6, 48 och 57 i denna, och
Det är nödvändigt att fastställa regleringsår för de produkter som anges i bilaga II till förordning (EG) nr 2200/96.
I artikel 26 i förordning (EG) nr 2200/96 fastställs gemenskapskompensationen för återtagande av de produkter som anges i bilaga II till den förordningen. Det är lämpligt att föreskriva ett system för utbetalning för att på så sätt hela tiden iaktta de begränsningar som föreskrivs i artikel 23 i förordning (EG) nr 2200/96.
I artikel 30.1 a första andra och tredje strecksatsen i ovannämnda förordning föreskrivs att frukt och grönsaker som återtas från marknaden i enlighet med artikel 23.1 i den förordningen och som förblivit osålda, får delas ut gratis, både inom gemenskapen och utom gemenskapen, som humanitärt bistånd till vissa nödlidande befolkningskategorier med hjälp av välgörenhetsorganisationer. Det är i detta syfte lämpligt att föreskriva att dessa välgörenhetsorganisationer skall godkännas på förhand.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 3
b) den produktion som medlemmarna i producentorganisationen sålde direkt enligt de villkor som avses i artikel 11.1 c 3 första och fjärde strecksatsen i förordning (EG) nr 2200/96,
2. Den saluförda produktion som avses i artikel 23.4 i förordning (EG) nr 2200/96 skall likställas med den saluförda kvantiteten definierad enligt punkt 1.
Regleringsåren för produkter som avses i artikel 1.2 i förordning (EG) nr 2200/96 andra än de som avses i första stycket, sträcker sig från den 1 januari till den 31 december.
a) medlemmarnas produktion som faktiskt sålts genom eller bearbetats av producentorganisationen,
3. Vid behandlingen av varje ansökan skall medlemsstaterna för de sammanlagda kvantiteter som inte saluförts efter inledningen av varje regleringsår i fråga kontrollera att de begränsningar som föreskrivs i artiklarna 23 och 24 i förordning (EG) nr 2200/96 efterlevs. Om ett överskridande sker skall gemenskapskompensation för återtagande endast utgå under förutsättning att dessa begränsningar respekteras med hänsyn till den kompensation som redan utgått. De överskridande kvantiteterna skall återtas vid behandlingen av nästa ansökan.
Artikel 7
Artikel 8
a) De tillgängliga lagren av äpplen och päron den första dagen i varje månad.
1. Före den 10 i varje månad skall medlemsstaterna på elektronisk väg till kommissionen översända en uppskattning fördelad per produkt av de produkter som inte saluförts under föregående månad.
b) senast den 30 november som följer på varje regleringsår för citroner, päron, äpplen, satsumas, clementiner och söta apelsiner.
Artikel 11
a) följa bestämmelserna i denna förordning,
3. Medlemsstaterna skall godkänna välgörenhetsorganisationer i minst en av följande kategorier:
Artikel 12
Medlemsstaterna skall vidta nödvändiga åtgärder för att underlätta kontakter och transaktioner mellan de berörda producentorganisationerna och de välgörenhetsorganisationer som godkänts i enlighet med artikel 11.2.
1. Gratis utdelning som sker utanför gemenskapen inom ramen för humanitärt bistånd skall genomföras av sådana välgörenhetsorganisationer som avses i artikel 11.3 c, enligt punkterna 2 och 3 i denna artikel.
1. Transportkostnader knutna till insatser för gratis utdelning av alla produkter som återtagits från marknaden skall betalas av garantisektionen inom Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) på grundval av schablonbelopp som fastställs utifrån avståndet mellan platsen för återtagandet och leveransplatsen och som anges i bilaga V.
Utbetalningen av beloppen skall ske på villkor att intyg läggs fram som bekräftar
- ett övertagandeintyg utfärdat av välgörenhetsorganisationen,
1. När det gäller återtagna äpplen och citrusfrukter skall sorterings- och förpackningskostnader i samband med gratis utdelning betalas av garantisektionen inom EUGFJ och inom gränsen för de belopp som anges i bilaga V.2, om det rör sig om gratis utdelning inom ramen för ett avtal mellan de berörda producent- och välgörenhetsorganisationerna.
4. Avtalen skall slutas för ett enda regleringsår i den mening som avses i förordning (EG) nr 2200/96 och skall innehålla uppgifter om
- den planerade leveranstakten,
- en uppskattning av antalet stödmottagare per administrativ enhet.
- namnet på de mottagande organisationerna,
- ett övertagandeintyg som utfärdats av välgörenhetsorganisationen.
2. Medlemsstaterna skall minst en gång per regleringsår genomföra fysiska kontroller och dokumentkontroller av alla producentorganisationernas återtagande transaktioner. Dessa kontroller skall för varje produkt gälla minst 20 % av den totala återtagna kvantiteten.
3. Medlemsstaterna skall genomföra dokumentkontroller av interventionerna för att effektivt fastställa att redovisningen utförs på ett korrekt sätt samt att betalningsvillkoren uppfylls för gemenskapskompensation för återtagande eller om finansiering genom driftsfonden, som avses i artikel 15.1 i förordning (EG) nr 2200/96.
Artikel 18
c) produkternas slutliga bestämmelseort.
4. På begäran av medlemsstaten skall kommissionen bistå medlemsstaten vid kontrollen av de gratisutdelningar som genomförs utanför gemenskapen.
a) de produkter som inte saluförts inte överensstämmer med de normer som avses i artikel 2 i förordning (EG) nr 2200/96,
2. De återtagna beloppen samt räntan skall betalas till den behöriga utbetalande organisationen och avräknas de kostnader som finansieras av EUGFJ.
1. Om det vid kontroller i enlighet med artikel 18 konstateras oegentligheter som kan tillskrivas producentorganisationer godkända välgörenhetsorganisationer eller institutionerna som avses i artiklarna 11 och 12 skall bestämmelserna i punkt 2-7 i denna artikel tillämpas.
4. Välgörenhetsorganisationen eller den institution som tagit emot produkten som återtagits från marknaden skall återbetala värdet av de produkter som ställts till dess förfogande ökat med en ränta beräknad på grundval av den tid som förflutit mellan mottagandet av produkten och mottagarens återbetalning.
7. De återtagna beloppen samt räntan skall betalas till det behöriga utbetalande organet och avräknas från de utgifter som finansieras av EUGFJ.
De producentorganisationer som ansökt om godkännande av ett operativt program i enlighet med artiklarna 3 eller 15 i förordning (EG) nr 411/97 får som en tillfällig åtgärd för 1997 på egen risk och i enlighet med artikel 15.3 b i förordning (EG) nr 2200/96 bevilja ett tillägg till gemenskapens ersättning för återtagande.
Artikel 24
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I artikel 2 i förordning (EG) nr 2200/96 fastställs att kommissionen, när den antar normer för färsk frukt och färska grönsaker, skall beakta Ekonomiska kommissionens för Europa (FN) internationella normer.
De förordningar i vilka normer för kronärtskockor, bönor, ärtor, blomkål och vitlök föreskrivs innehåller inga bestämmelser om angivelse av ursprungsland på förpackningen. Bestämmelser av denna art i gällande internationella normer bör införas i dessa förordningar.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för frukt och grönsaker.
Texten i A "Identifiering" skall ersättas med följande:
Texten i C "Produktens ursprung" skall ersättas med följande:
3. Förordning nr 211/66/EEG skall upphöra att gälla.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De allmänna reglerna för hur Kombinerade nomenklaturen skall tolkas har fastställts i förordning (EEG) nr 2658/87. Dessa regler skall också tillämpas på all annan nomenklatur som baseras på denna, även om detta gäller endast delvis eller om underuppdelningar eventuellt gjorts som tillägg till den, och som fastställts genom särskilda gemenskapsbestämmelser för tillämpningen av tullmässiga eller andra åtgärder inom ramen för varuutbytet.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från sektionen för tulltaxe- och statistiknomenklatur inom tullkodexkommittén.
De varor som beskrivs i första kolumnen i tabellen i bilagan hänförs till de nummer i Kombinerade nomenklaturen som anges i andra kolumnen i samma tabell.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I artikel 4 andra strecksatsen i förordning (EG) nr 2027/95 föreskrivs att kommissionen på en medlemsstats begäran skall vidta lämpliga åtgärder så att denna medlemsstat skall kunna utnyttja sina kvoter i enlighet med bestämmelserna i artikel 6.2 tredje stycket i rådets förordning (EG) nr 685/95 av den 27 mars 1995 om administreringen av fiskeinsatsen med avseende på vissa fiskezoner och -resurser i gemenskapen (2).
Förvaltningskommittén för fiskeresurser har avgivit sitt yttrande.
Den årliga maximala fiskeansträngningsnivån för Nederländerna för fiske med släpredskap, bottenlevande arter, som anges i bilaga I till förordning (EG) nr 2027/95 skall anpassas i enlighet med vad som anges i bilagan.
KOMMISSIONENS FÖRORDNING (EG) nr 1365/97 av den 16 juli 1997 om ändring av förordning (EG) nr 716/96 om undantagsåtgärder till stöd för nötköttsmarknaden i Förenade kungariket
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött (1), senast ändrad genom kommissionens förordning (EG) nr 2222/96 (2), särskilt artikel 23 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- 0,8 ecu per kg levande vikt när det gäller kor, och
2. Där det är nödvändigt att väga berörda djur efter slakt för att beräkna vad den levande vikten skulle ha varit, skall man multiplicera slaktvikten efter avblodning, avhudning, urtagning samt avlägsnande av klövar och hud med en koefficient på
3. Gemenskapen skall medfinansiera den utgift som Förenade kungariket haft för de inköp som avses i artikel 1.1 till ett pris av 291 ecu per inköpt ko och 328 ecu per inköpt djur för alla andra djur som har destruerats i enlighet med bestämmelserna i artikel 1.
Producenten eller hans ombud förbinder sig att försäkra att detta bidrag inte har sökts för djuret i fråga.
Artikel 2
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
i enlighet med förfarandet i artikel 189 c i fördraget (2), och med beaktande av följande:
Inom ramen för kampen mot utbudet av narkotika är det synnerligen väsentligt att fattigdomen i söder minskas radikalt och att befolkningen erbjuds ett lagligt alternativ till den olagliga odlingen.
Europaparlamentet avgav ett yttrande om dessa riktlinjer den 15 juni 1995.
Europeiska gemenskapen är part i konventionen från 1988, särskilt i kraft av dess artikel 12, och har antagit gemenskapslagstiftning som syftar till kontroll över handeln med prekursorer, efter rekommendationer från den aktionsgrupp för kemiska produkter (GAPC) som skapades av G7 och ordföranden i EG-kommissionen 1989; en grupp som skulle kunna bli effektivare globalt sett om lämplig lagstiftning och lämpliga förfaranden antogs i andra delar av världen.
Europeiska gemenskapens medlemsstater har skrivit under den politiska deklarationen och det globala åtgärdsprogram som antogs av Förenta nationernas generalförsamling vid dess 17:e extramöte.
Artikel 1
Det bistånd som ges i enlighet med denna artikel skall komplettera och förstärka bistånd som lämnas enligt andra instrument för utvecklingssamarbete.
Att förebygga narkotikamissbruk och att minska efterfrågan bör ingå som åtgärder i en konsekvent politik som innefattar utbildning och objektiv information om följderna av narkotikamissbruk, främst riktad mot de unga.
Gemenskapen skall helst arbeta inom den strategiska ram som har lagts fast i de nationella planerna, och skall även stödja särskilda aktioner med mätbar inverkan (dvs. effektiva och påtagliga resultat inom en i förväg fastställd tidsperiod) på följande områden:
- avtalen mellan gemenskapen och vissa utvecklingsländer skall kunna genomföras, särskilt när det gäller att bekämpa att kemiska prekursorer kommer på avvägar och kampen mot penningtvätt.
- finansiering av studier, seminarier och forum för erfarenhetsutbyte inom ovannämnda områden.
Artikel 5
1. De instrument som skall användas för åtgärderna enligt artiklarna 3 och 4 skall innefatta studier, tekniskt bistånd, utbildning eller andra tjänster, leveranser och anläggningar, liksom även revision samt utvärderings- och övervakningsuppdrag.
4. Ekonomiska bidrag från lokala samarbetsparter, i synnerhet till driftskostnaderna, skall sökas som en prioriterad åtgärd när det gäller projekt med syfte att sätta igång långsiktig verksamhet, för att på så sätt säkerställa att sådana projekt lever vidare då gemenskapsbidragen upphör.
7. För att kunna uppnå fördragets mål om konsekvens och komplementaritet och i syfte att optimera effekten av alla dessa åtgärder kan kommissionen vidta alla de nödvändiga samordningsåtgärderna, i synnerhet
8. I syfte att få största möjliga verkan så väl globalt som nationellt, skall kommissionen tillsammans med medlemsstaterna ta alla initiativ som krävs för att säkerställa god samordning och nära samarbete med mottagarländerna och bidragsgivarna samt andra internationella organ som berörs, i synnerhet de som ingår i Förenta nationernas organisation och då särskilt UNDCP.
Artikel 8
Artikel 9
- Effekten av och möjligheten att genomföra åtgärderna.
- Erfarenheter av åtgärder av samma typ.
4. Kommissionen bemyndigas att, utan dessförinnan höra den kommitté som avses i artikel 10, godkänna de ytterligare åtaganden som kan behövas för att täcka sådana överskridanden som kan förutses eller som har konstaterats i samband med dessa åtgärder om överskridandet uppgår till högst 20 % av det ursprungliga åtagande som fastställdes genom finansieringsbeslutet.
7. Deltagande i anbudsförfaranden och i avtal skall vara öppet på lika villkor för alla fysiska och juridiska personer i medlemsstaterna och mottagarlandet. Det kan utsträckas till andra utvecklingsländer.
- strävan efter kostnadseffektivitet och en varaktig inverkan i samband med att projekten utformas, och
1. Kommissionen skall biträdas av den behöriga geografiska kommittén för utvecklingssamarbete.
Om de planerade åtgärderna inte är förenliga med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Artikel 11
2. Kommissionen skall regelbundet utvärdera de åtgärder som gemenskapen finansierar för att fastställa om de mål som ställdes upp för dessa åtgärder har uppnåtts och för att ange riktlinjer för att förbättra framtida åtgärders effektivitet. Kommissionen skall överlämna en sammanfattning av de utvärderingar som gjorts till den kommitté som avses i artikel 10, vilka denna kommitté i förekommande skall kunna granska. Utvärderingsrapporterna skall finnas tillgängliga för de medlemsstater som önskar ta del av dem.
1. Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av följande: I artikel 17 i direktiv 94/67/EG fastställs att medlemsstaterna skall rapportera om genomförandet av detta direktiv i enlighet med artikel 5 i direktiv 91/692/EEG.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som upprättats i enlighet med artikel 6 i ovan nämnda direktiv.
Det frågeformulär som bifogas detta beslut, och som skall användas i samband med rådets direktiv 94/67/EG om förbränning av farligt avfall, antas härmed.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Att slå vakt om kvaliteten på landsbygdsmiljön är ett av målen för politiken för landsbygdens utveckling.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
av följande skål: Avtalet om ömsesidigt erkännande mellan Europeiska gemenskapen och Kanada, vilket undertecknades i London den 14 maj 1998, har framförhandlats och bör godkännas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Texten till avtalet och bilagorna till det bifogas detta beslut.
Artikel 3
3. I samtliga övriga fall skall gemenskapens ståndpunkt i den gemensamma kommittén eller i de gemensamma sektoriella grupperna fastställas av rådet som skall fatta sina beslut med kvalificerad majoritet på förslag av kommissionen. Samma förfarande skall gälla för beslut som fattas av gemenskapen inom ramen för artiklarna XV.3 och XIX.4 i avtalet.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113 i detta,
(2) Kreditförsäkringar för medellånga och långa exportaffärer spelar en viktig roll för handeln med utvecklingsländer och främjar dessa länders integrering med världsekonomin, vilket är ett mål för gemenskapens utvecklingspolitik.
(5) För att minska befintlig snedvridning av konkurrensen är det önskvärt att de olika statsstödda systemen för exportkreditförsäkringar harmoniseras enligt artikel 112 i fördraget, på grundval av enhetliga principer och på ett sådant sätt att de bildar en integrerad del av den gemensamma handelspolitiken.
(8) En harmonisering skulle gynna samarbete mellan de kreditförsäkrare som agerar på en stats vägnar eller med statligt stöd, och öka samarbetet mellan företag inom gemenskapen enligt artikel 130 i fördraget.
(11) Genom sitt beslut (2) av den 27 september 1960 inrättade rådet en arbetsgrupp för samordning av politiken för kreditförsäkringar, kreditgarantier och finansiella krediter.
(14) Rådets direktiv 70/509/EEG av den 27 oktober 1970 om antagande av gemensamma kreditförsäkringsvillkor för medellånga och långa exportaffärer med offentliga köpare (4), och rådets direktiv 70/510/EEG av den 27 oktober 1970 om antagande av gemensamma kreditförsäkringsvillkor för medellånga och långa exportaffärer med privata köpare (5), bör ersättas med det här direktivet.
Artikel 1
Detta direktiv gäller varken försäkringsskydd för anbud, förskottsbetalning eller fullgörandegarantier och inte heller försäkring för säkerhet för "retention money", så kallad retention payment bond. Det gäller inte heller försäkringsskydd för risker avseende byggutrustning och byggmaterial när dessa används lokalt för att fullgöra ett affärsavtal.
Medlemsstaterna skall se till att alla institut, som direkt eller indirekt erbjuder försäkringsskydd i form av exportkreditförsäkringar, garantier eller refinansiering för medlemsstatens räkning eller med stöd av den medlemsstat som företräder själva regeringen eller som kontrolleras av och/eller handlar enligt bemyndigande av den regering som erbjuder försäkringsskydd, nedan kallade försäkringsgivare, erbjuder försäkringsskydd för affärer avseende export av varor och/eller tjänster i enlighet med bestämmelserna i bilagan, när exportaffärerna görs med länder utanför gemenskapen och finansieras med hjälp av köparkrediter eller leverantörskrediter eller betalas kontant.
De beslut som avses i punkt 46 i bilagan skall fattas av kommissionen i enlighet med det förfarande som avses i artikel 4.
Kommissionen skall biträdas av en kommitté som skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
- Skall kommissionen uppskjuta verkställandet av de beslutade åtgärderna under en tid som inte överstiger en månad från den dag då rådet underrättats.
Rapport och översyn
Förhållande till andra förfaranden
Upphävande
Överföring
RÅDETS DIREKTIV 98/49/EG av den 29 juni 1998 om skydd av kompletterande pensionsrättigheter för anställda och egenföretagare som flyttar inom gemenskapen
med beaktande av kommissionens förslag (1),
av följande skäl: (1) En av de grundläggande friheterna i gemenskapen är fri rörlighet för personer. I fördraget föreskrivs att rådet enhälligt skall besluta om sådana åtgärder inom den sociala trygghetens område som är nödvändiga för att genomföra fri rörlighet för arbetstagare.
(4) Rådet äger stor frihet när det gäller valet av vilka åtgärder som är bäst lämpade för att uppnå målet i artikel 51 i fördraget; det samordningssystem som avses i förordningarna (EEG) nr 1408/71 och (EEG) nr 574/72, och särskilt reglerna för sammanläggning, passar inte för kompletterande pensionssystem, med undantag för system som täcks av begreppet "lagstiftning" enligt definitionen i artikel 1 j första stycket i förordning (EEG) nr 1408/71 eller med avseende på vilka en medlemsstat avger en förklaring enligt den artikeln, och bör därför bli föremål för särskilda åtgärder, av vilka detta direktiv är den första, så att hänsyn kan tas till deras särskilda karaktär och kännetecken och till olikheterna mellan sådana system inom och mellan medlemsstaterna.
(7) Ett bidrag till att nå detta mål kan vara att arbetstagare, som flyttar eller vilkas arbetsplats flyttar från en medlemsstat till en annan, i fråga om skyddet för deras kompletterande pensionsrättigheter garanteras en behandling som är likvärdig med den som ges arbetstagare som stannar kvar eller vilkas arbetsplats stannar kvar inom samma medlemsstat.
(10) För att rätten till fri rörlighet skall kunna utövas på ett effektivt sätt bör arbetstagare och andra berättigade personer ha vissa garantier för lika behandling i fråga om bevarandet av sina intjänade pensionsrättigheter enligt kompletterande pensionssystem.
(13) I detta avseende krävs enligt fördraget inte bara avskaffande av diskriminering av arbetstagare i medlemsstaterna på grund av medborgarskap utan även undanröjande av alla nationella bestämmelser som kan hindra dessa arbetstagares utövande av, eller göra det mindre attraktivt för dem att utöva, de grundläggande friheter som garanteras i fördraget, enligt Europeiska gemenskapernas domstols tolkning i flera på varandra följande domar.
(16) På grund av mångfalden av kompletterande system för social trygghet bör gemenskapen endast ställa upp allmänna mål och därför är ett direktiv det lämpliga rättsliga instrumentet.
KAPITEL I
Syftet med detta direktiv är att skydda rättigheterna för de försäkringstagare som omfattas av kompletterande pensionssystem och som flyttar från en medlemsstat till en annan och att därigenom bidra till att undanröja hinder för den fria rörligheten för anställda och egenföretagare inom gemenskapen. Detta skydd avser pensionsrättigheter enligt både frivilliga och obligatoriska kompletterande pensionssystem, med undantag av de system som omfattas av förordning (EEG) nr 1408/71.
KAPITEL II
I detta direktiv används följande beteckningar med de betydelser som här anges:
c) pensionsrättigheter: alla förmåner som försäkringstagare och andra berättigade personer har rätt till enligt bestämmelserna i ett kompletterande pensionssystem och, i förekommande fall, enligt nationell lagstiftning,
f) avgift: alla betalningar som gjorts eller anses ha gjorts till ett kompletterande pensionssystem.
Artikel 4
Artikel 5
Artikel 6
2. Om avgifter fortsatt betalas in till ett kompletterande pensionssystem i en medlemsstat i enlighet med punkt 1, skall den utsända arbetstagaren och, i förekommande fall, dennas arbetsgivare, vara undantagen från alla förpliktelser att betala in avgifter till ett kompletterande pensionssystem i en annan medlemsstat.
Medlemsstaterna skall vidta åtgärder så att arbetsgivare, förvaltare eller andra, som har ansvar för förvaltningen av de kompletterande pensionssystemen, när försäkringstagarna flyttar till en annan medlemsstat förser dem med adekvat information i fråga om deras pensionsrättigheter och om de valmöjligheter som finns att tillgå för dem enligt systemet. Denna information skall minst motsvara den information som ges de försäkringstagare för vilka avgifter inte längre betalas men som bor kvar i samma medlemsstat.
Artikel 8
Medlemsstaterna skall i sin nationella lagstiftning införa de bestämmelser som behövs för att alla, som anser sig förfördelade på grund av underlåtenhet att tillämpa bestämmelserna i detta direktiv, skall kunna föra talan vid domstol, efter att i förekommande fall ha vänt sig till andra behöriga myndigheter.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
3. På grundval av de upplysningar som medlemsstaterna lämnar skall kommissionen inom sex år efter detta direktivs ikraftträdande överlämna en rapport som till Europaparlamentet, rådet och Ekonomiska och sociala kommittén.
RÅDETS DIREKTIV 98/57/EG av den 20 juli 1998 om bekämpning av Ralstonia solanacearum (Smith) Yabuuchi m.fl.
med beaktande av kommissionens förslag (1),
av följande skäl: Skadegöraren Ralstonia solanacearum (Smith) Yabuuchi m.fl. var tidigare känd som Pseudomonas solanacearum (Smith) Smith. Ralstonia solanacearum (Smith) Yabuuchi m.fl. kommer förmodligen att bli det allmänt godtagna namnet på skadegöraren. I detta direktiv bör hänsyn tas till denna vetenskapliga utveckling.
Skyddsåtgärder mot införsel av skadegörare till en medlemsstats territorium skulle endast ha begränsad effekt om inte sådana skadegörare samtidigt och metodiskt bekämpades inom hela gemenskapen och hindrades från att sprida sig.
För att säkerställa detta måste vissa åtgärder vidtas inom gemenskapen. Medlemsstaterna måste dessutom kunna vidta ytterligare eller strängare åtgärder, där detta är nödvändigt förutsatt att dessa inte hindrar handeln med potatis eller tomater inom gemenskapen än de som anges i rådets direktiv 77/93/EEG av den 21 december 1976 om skyddsåtgärder mot att skadegörare på växter eller växtprodukter förs in till medlemsstaterna (4). Sådana åtgärder måste anmälas till de andra medlemsstaterna och till kommissionen.
Den nuvarande kunskapen om de biologiska och epidemiologiska egenskaperna hos Ralstonia solanacearum (Smith) Yabuuchi m.fl. under europeiska förhållanden är ofullständig, och det förutses att en översyn av de föreslagna åtgärderna kommer att bli nödvändig om ett antal säsonger. Förbättringar av testprocedurerna förväntas också mot bakgrund av ytterligare forskning, särskilt kring testmetodernas sensibilitet och noggrannhet, för att optimala testmetoder skall kunna väljas ut och standardiseras.
Artikel 1
b) förhindra dess förekomst och spridning, och
1. Medlemsstaterna skall varje år genomföra systematiska officiella undersökningar för att kontrollera förekomst av skadegöraren på det förtecknade växtmaterialet med ursprung i deras territorium. För att identifiera andra möjliga smittkällor som hotar produktionen av det förtecknade växtmaterialet skall medlemsstaterna göra en riskbedömning och, om ingen risk för spridning av skadegöraren har konstaterats under den bedömningen skall de, i produktionsområdena för det förtecknade växtmaterialet, genomföra riktade officiella undersökningar för att kontrollera förekomst av skadegöraren på andra växter än det förtecknade växtmaterialet, även på vilda värdväxter av familjen Solanaceae samt på ytvatten som används för bevattning eller duschning av det förtecknade växtmaterialet och på flytande avfall som släpps ut från anläggningar för industriell bearbetning eller förpackning där det förtecknade växtmaterialet hanteras och som används för bevattning och duschning av det förtecknade växtmaterialet. Omfattningen av dessa riktade undersökningar skall bestämmas med beaktande av den konstaterade risken. Medlemsstaterna kan också utföra officiella undersökningar för att kontrollera förekomst av skadegöraren på annat material, t.ex. odlingssubstrat, jord och fast avfall från anläggningar för industriell bearbetning eller förpackning.
b) på värdväxter som inte återfinns i det förtecknade växtmaterialet och på vatten, inklusive flytande avfall, i enlighet med lämpliga metoder, och stickprov skall, när så är lämpligt, tas och genomgå officiella eller officiellt övervakade laboratorietest, och
3. Resultaten av och detaljerna i fråga om de officiella undersökningar som fastställs i punkt 1 skall varje år anmälas till de andra medlemsstaterna och till kommissionen i enlighet med bestämmelserna i punkt 2 i avsnitt II i bilaga I. Dessa anmälningar skall göras senast den 1 juni, med undantag av anmälningar om utsädespotatis som skall ges in före den 1 september. Detaljerna och resultaten ifråga om grödor skall avse föregående års produktion. Innehållet i dessa anmälningar kan överlämnas till kommittén.
5. Följande bestämmelser får antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
Artikel 3
1. Vid varje fall av misstänkt förekomst av skadegöraren skall de ansvariga officiella organen i den berörda medlemsstaten eller de berörda medlemsstaterna säkerställa att officiella eller officiellt övervakade laboratorietest genomförs på det förtecknade växtmaterialet enligt den lämpliga metod som anges i bilaga II och enligt de villkor som anges i punkt 1 i bilaga III, eller, i andra fall, någon annan officiellt godkänt metod, för att bekräfta eller vederlägga den misstänkta förekomsten. Om misstanken bekräftas skall de krav som fastställs i punkt 2 i bilaga III gälla.
a) förbjuda flyttning av plantor och knölar från alla grödor, partier eller sändningar från vilka stickproven har tagits, förutom då det sker under deras övervakning och förutsatt att det har konstaterats att det inte finns någon identifierbar risk för att skadegöraren skall spridas,
3. I fall av misstänkt förekomst av skadegöraren skall, om det finns risk för angrepp på det förtecknade växtmaterialet eller ytvattnet från eller till en annan medlemsstat, den medlemsstat där misstanken har rapporterats omedelbart till den eller de andra berörda medlemsstaterna, beroende på den konstaterade risken, anmäla den nämnda misstänkta förekomsten, och de nämnda medlemsstaterna skall då samarbeta på lämpligt sätt. Den eller de medlemsstater som fått anmälan skall vidta försiktighetsåtgärder enligt punkt 2 c och i förekommande fall vidta ytterligare åtgärder enligt punkterna 1 och 2.
Artikel 5
i) Genomföra en utredning för att, i enlighet med bestämmelserna i bilaga IV, fastställa angreppets omfattning och dess primärkälla eller -källor, med ytterligare test i enlighet med artikel 4.1 på åtminstone alla lager av utsädespotatis ur kloner som är närbesläktade.
iv) Avgränsa ett område på grundval av förklaringen om angreppet enligt punkt ii, fastställa omfattningen av det troliga angreppet enligt punkt iii och skadegörarens möjliga spridning, i enlighet med bestämmelserna i punkt 2 i i bilaga V.
ii) Förklara de av skadegörarens värdväxter som provet har tagits från för angripna.
i) Genomföra en utredning som omfattar en officiell undersökning vid lämpliga tidpunkter på prov av ytvattnet och, om sådana finns, på vilda värdväxter av familjen Solanaceae för att fastställa angreppets omfattning.
2. Medlemsstaterna skall, i enlighet med bestämmelserna i punkt 3 i bilaga V, omedelbart till de andra medlemsstaterna och till kommissionen anmäla varje angrepp som fastställs enligt punkterna 1 a ii och 1 c ii och uppgifterna om avgränsning av områden enligt punkt 1 a iv och, där så är tillämpligt, enligt punkt 1 c iii. Innehållet i denna anmälan enligt detta stycke får överlämnas till kommittén.
Artikel 6
3. Medlemsstaterna skall föreskriva att alla maskiner, fordon, fartyg, lager, eller delar av dessa, och alla andra föremål, inklusive förpackningsmaterial, som har förklarats angripna enligt artikel 5.1 a ii eller förklarats troligen angripna enligt artikel 5.1 a iii och 5.1 c iii, antingen skall förstöras eller saneras med lämpliga metoder som fastställs i punkt 3 i bilaga VI. Efter saneringen skall inga sådana föremål längre betraktas som angripna.
1. Medlemsstaterna skall föreskriva att utsädespotatis skall uppfylla kraven i direktiv 77/93/EEG och att de i direkt led skall härstamma ur potatismaterial som erhållits enligt ett officiellt godkänt program och som har konstaterats vara fritt från skadegöraren vid officiella eller officiellt övervakade tester då den lämpliga metod, som anges i bilaga II, har använts.
i) genom tester av tidigare generationer inklusive det ursprungliga klonurvalet och systematiska tester av det ursprungliga klonurvalet av utsädespotatisen, eller
2. Följande bestämmelser får antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
Artikel 8
Utan att det påverkar tillämpningen av bestämmelserna i direktiv 77/93/EEG får bestämmelserna bevilja undantag från de åtgärder som avses i artiklarna 6 och 8 i det här direktivet i enlighet med bestämmelserna i direktiv 95/44/EG i experimentellt eller vetenskapligt syfte och för växtförädling (5).
Ändringar i bilagorna till detta direktiv mot bakgrund av nya vetenskapliga eller tekniska rön skall antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG. När det gäller de metoder som anges i bilaga II och åtgärderna i punkt 4.1 och 4.2 i bilaga VI till detta direktiv, skall kommissionen förbereda en rapport där metoderna och åtgärderna granskas mot bakgrund av gjorda erfarenheter som vunnits, och rapporten skall överlämnas till kommittén före den 1 januari 2002.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning till detta direktiv när de offentliggörs. Närmare föreskrifter för hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
RÅDETS DIREKTIV 98/93/EG av den 14 december 1998 om ändring av direktiv 68/414/EEG om en skyldighet för medlemsstaterna i EEG att inneha minimilager av råolja och/eller petroleumprodukter
med beaktande av kommissionens förslag (1),
av följande skäl: (1) Den 20 december 1968 antog rådet direktiv 68/414/EEG om en skyldighet för medlemsstaterna i EEG att inneha minimilager av råolja och/eller petroleumprodukter (4).
(4) Det är viktigt att öka försörjningssäkerheten för olja.
(7) I enlighet med subsidiaritetsprincipen och proportionalitetsprincipen fastställd i artikel 3b i fördraget går det lättare att på gemenskapsnivå uppnå målet att upprätthålla en hög nivå av försörjningssäkerhet för olja i gemenskapen genom säkra system, som är öppna för insyn och som bygger på solidaritet mellan medlemsstaterna, och som samtidigt uppfyller bestämmelserna om den inre marknaden och om konkurrens. Detta direktiv sträcker sig inte utöver vad som behövs för att uppnå detta mål.
(10) Lagerhållningssystemen bör bygga på öppenhet för insyn för att säkerställa att den börda som lagerhållningsskyldigheten innebär fördelas rättvist och utan någon diskriminering. Medlemsstaterna kan göra information om kostnaden för att hålla oljelager tillgänglig för berörda parter.
(13) Det är lämpligt att tillämpa tillvägagångssätt som gemenskapen och medlemsstaterna redan följer inom ramen för sina internationella skyldigheter och avtal. På grund av förändringar i oljeförbrukningsmönstret har flygbränsle för internationell luftfart blivit ett viktigt inslag i denna förbrukning.
(16) För att säkerställa att den inre marknaden fungerar smidigt är det önskvärt att främja användningen av avtal mellan medlemsstater när det gäller minimilagerhållning för att främja användningen av lageranläggningar i andra medlemsstater. Beslut att ingå sådana avtal skall fattas av de berörda medlemsstaterna.
(19) Det är lämpligt att med jämna mellanrum informera rådet om läget beträffande beredskapslagren i gemenskapen.
Direktiv 68/414/EEG ändras på följande sätt:
3. Nuvarande artikel 3 skall betecknas artikel 2 och skall kompletteras med följande stycke:
Medlemsstaterna skall till kommissionen överlämna ett statistiskt sammandrag över de lager som finns i slutet av varje månad, upprättat enligt artiklarna 5 och 6 och med närmare angivande av antalet dagar med genomsnittlig förbrukning under det föregående kalenderåret som dessa lager representerar. Detta sammandrag skall överlämnas senast den tjugofemte dagen i den andra månaden efter den månad som sammandraget avser.
"Artikel 5
- fördelade i förhållande till de kvantiteter av varje produktkategori som erhållits under föregående kalenderår från den berörda statens raffinaderier, eller
Blandningsprodukter får, när de är avsedda för bearbetning till de färdiga produkter som anges i artikel 2, tjäna som ersättning för de produkter för vilka de är avsedda." 7. Artikel 6 skall ändras enligt följande:
"2. För genomförandet av detta direktiv får lager, enligt avtal mellan regeringar, upprättas inom en medlemsstats territorium för företag eller organ/enheter som är etablerade i en annan medlemsstat. Beslut om att hålla en del av sina lager utanför sitt nationella territorium skall fattas av den berörda medlemsstatens regering.
Utkast till de avtal som nämns i första stycket skall överlämnas till kommissionen, som får lämna sina kommentarer till de berörda regeringarna. När avtalen väl har ingåtts skall de anmälas till kommissionen, som skall underrätta de övriga medlemsstaterna om dem.
- De skall fastställa villkor och tillvägagångssätt för lagerhållning som är inriktade på att trygga kontrollen av lagren och deras tillgänglighet.
- De skall, om en part kan säga upp avtalet, föreskriva att sådan uppsägning inte skall gälla i händelse av en försörjningskris och att kommissionen under alla förhållanden skall erhålla förhandsinformation om uppsägning sker.
- Minsta avtalsperiod skall vara 90 dagar.
- Det företag, organ/enhet som håller lagren för det företag, organ/enhet som har rätt till dem, skall vara underkastad lagstiftningen i den medlemsstat på vars territorium lagren befinner sig, när det gäller den medlemsstatens lagliga befogenheter att kontrollera och verifiera förekomsten av lagren." c) Punkt 3 andra stycket skall ersättas med följande:
Medlemsstaterna skall anta alla bestämmelser som är nödvändiga och vidta alla åtgärder som är nödvändiga för att säkerställa kontrollen och övervakningen av lagren. De skall inrätta system för verifiering av lagren i enlighet med bestämmelserna i detta direktiv."
Medlemsstaterna skall bestämma vilka straff som skall gälla för överträdelser av de nationella bestämmelser som antas i enlighet med detta direktiv och vidta alla åtgärder som är nödvändiga för att säkerställa genomförandet av dessa bestämmelser. Straffen skall vara effektiva, proportionerliga och avskräckande."
Artikel 3
Artikel 4
Kommissionen skall regelbundet till rådet överlämna en rapport om läget beträffande lagren i gemenskapen, inbegripet, när så är lämpligt, om behovet av en harmonisering för att säkerställa en effektiv kontroll och övervakning av lagren. Den första rapporten skall överlämnas till rådet under det andra året efter det datum som fastställs i artikel 3.1.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
I enlighet med förordning (EEG) nr 2377/90 måste gränsvärden för högsta tillåtna restmängder successivt fastställas för samtliga farmakologiskt verksamma substanser som används inom gemenskapen i veterinärmedicinska läkemedel som är avsedda att ges till livsmedelsproducerande djur.
För kontroll av resthalter bör enligt tillämplig gemenskapslagstiftning gränsvärden vanligtvis fastställas för målvävnaderna lever eller njure. I den internationella handeln avlägsnas dock ofta lever och njure från slaktkroppen, och gränsvärden bör därför alltid fastställas även för muskel- eller fettvävnader.
Lini oleum, folsyra, betain och cefazolin skall införas i bilaga II till förordning (EEG) nr 2377/90.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
Bilaga I, II och III till förordning (EEG) nr 2377/90 skall ändras i enlighet med bilagan till den här förordningen.
KOMMISSIONENS FÖRORDNING (EG) nr 179/98 av den 23 januari 1998 om ändring av rådets förordning (EG) nr 3051/95 om säkerhetsorganisation för roll-on/roll-off-passagerarfartyg (ro-ro-fartyg)
med beaktande av rådets förordning (EG) nr 3051/95 av den 8 december 1995 om säkerhetsorganisation för roll-on/roll-off-passagerarfartyg (ro-ro-fartyg) (1), särskilt artikel 9 i denna, och
Det är nödvändigt att ta hänsyn till utvecklingen på det internationella planet genom att införa närmare bestämmelser om utfärdandet av interimistiska dokument och certifikat, formulär för ISM-dokument och ISM-certifikat samt vissa standarder avseende ISM-certifieringsarrangemang.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som inrättats enligt artikel 12 i rådets direktiv 93/75/EEG (2), senast ändrat genom kommissionens direktiv 97/34/EG (3).
KOMMISSIONENS FÖRORDNING (EG) nr 496/98 av den 27 februari 1998 om klassificering av vissa varor i Kombinerade nomenklaturen
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 2509/97 (2), särskilt artikel 9 i denna, och med beaktande av följande:
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från sektionen för tulltaxe- och statistiknomenklatur inom tullkodexkommittén.
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Genom kommissionens förordning (EEG) nr 3077/78 (3), senast ändrad genom förordning (EG) nr 2132/95 (4), godkänns intyg för humle som importeras från vissa tredje länder såsom likvärdiga med gemenskapsintygen samt upprättas en förteckning över de förvaltningar i dessa länder som har befogenhet att utfärda likvärdiga intyg, liksom en förteckning över de produkter som omfattas. Till följd av de uppgifter som Polen har lämnat in är det nödvändigt att ändra bilagan till förordning (EEG) nr 3077/78.
Artikel 1
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Enligt artikel 5.1 fjärde strecksatsen i kommissionens förordning (EEG) nr 3719/88 av den 16 november 1988 om gemensamma tillämpningsföreskrifter för systemet med import- och exportlicenser och förutfastställelselicenser för jordbruksprodukter (5), senast ändrad genom förordning (EG) nr 1404/97 (6), krävs ingen licens för export vid en säkerhet på högst 5 ecu. Det låga säkerhetsbeloppet för export utan bidrag innebär att mycket skulle kunna exporteras utan licens, vilket skulle försvaga kontrollen av kvantiteterna i fråga. För att undvika den risken bör särskilda villkor gälla i nämnda fall.
Artikel 1
2. Artikel 2 skall ändras på följande sätt:
a) 10 ecu per 100 kg netto för licenser med förutfastställelse av bidraget,
"4. Genom undantag från artikel 5.1 fjärde strecksatsen i förordning (EEG) nr 3719/88 skall ingen licens krävas vid export av en kvantitet på 50 kg eller mindre."
"1. Ansökningar om exportlicenser med förutfastställelse av bidraget skall inlämnas hos den behöriga myndigheten från och med tisdag till och med torsdag varje vecka. Ansökningar som inlämnas en måndag eller fredag skall behandlas som om de vore inlämnade närmast följande tisdag."
3. Den sista meningen i punkt 3 skall ersättas med följande:
"I de fall den enhetliga procentsatsen för godkännande på under 80 % endast gäller de licenser som är bidragsberättigande, får operatören begära att en licens som inte berättigar till bidrag skall utfärdas inom samma tidsfrist för den kvantitet som inte har godkänts."
4. Artikel 5 skall ändras på följande sätt:
"a) de ansökningar om exportlicenser med förutfastställelse av bidraget, vilka har lämnats in från och med tisdag till och med torsdag i enlighet med artikel 3.1."
"Det meddelande om ansökningar som avses i punkt 1 a och, vad gäller tillämpningen av artikel 3.5 de upplysningar som avses i punkt 1 b, skall innehålla följande:"
"Dessa upplysningar skall anges separat om licenser för livsmedelshjälp utfärdas."
5. I bilagan skall delarna B och D ersättas med de som anges i bilagan till denna förordning.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EG) nr 3072/95 av den 22 december 1995 om den gemensamma organisationen av marknaden för ris (3), ändrad genom förordning (EG) nr 192/98 (4), särskilt artikel 7 i denna, och
För att den särskilda säkerheten skall kunna frisläppas för framför allt förestrad och företrad stärkelse är det lämpligt att fastställa de huvudsakliga krav som måste vara uppfyllda. De särskilda bestämmelser som gäller för dessa produkter bör även fortsättningsvis kompletteras med vissa åtgärder inriktade på effektiviteten i kontroller och på sanktioner i fall då villkoren för bearbetning och användning inte iakttas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Bidraget per ton stärkelse av majs, vete, korn, havre, potatis, ris eller brutet ris skall beräknas framför allt på grundval av skillnaden mellan
multiplicerad med koefficienten 1,60.
2) I artikel 6 skall punkterna 3 och 4 ersättas med följande:
4. Den bidragssats som är tillämplig och anges i licensen skall vara den som gäller den dag då ansökan inkommer.
"Det primära kravet, enligt artikel 20 i förordning (EEG) nr 2220/85, är att produkten skall användas eller exporteras i enlighet med de respektive bestämmelserna i artikel 10.1 a och 10.1 b i denna förordning. Användningen eller exporten skall ske inom tolv månader efter det att licensens giltighet har löpt ut. En förlängning av detta slutdatum med som mest sex månader får övervägas på grundval av en välgrundad begäran som lagts fram för den behöriga myndigheten."
5) Artikel 12 skall ersättas med följande: "Artikel 12
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Till följd av de tre nya medlemsstaternas anslutning räknas den tidsfrist på sex månader som föreskrivs i artikel 17 i förordning (EEG) nr 2081/92 från deras anslutningsdag. Vissa av de beteckningar som meddelats av medlemsstaterna överensstämmer med artiklarna 2 och 4 i nämna förordning och bör därför registreras.
Artikel 1
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De jordbruksrelaterade komponenterna i dessa substrat bör i princip komma från jordbruksföretag där en ekologisk produktionsmetod används.
Det bör dock övervägas ytterligare förbättringar av bestämmelserna i denna förordning. Detta gäller särskilt bestämmelserna om villkoren för användning, inbegripet villkoren för högsta tillåtna procentandel gödsel som inte kommer från jordbruksföretag där en ekologisk produktionsmetod används samt mycelets egenskaper och ursprung. Det förberedande arbetet bör inledas i tillräckligt god tid så att det kan avslutas innan övergångsperioden går ut.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
- produkter som anges i punkt 5.1 a i bilagan och som inte kommer från jordbruksföretag där en ekologisk produktionsmetod används, men som uppfyller de krav som anges i del A första till fjärde strecksatsen i bilaga II till förordning (EEG) nr 2092/91, och/eller
I dessa fall skall märkningen och annonseringen innehålla uppgiften "Svamp som odlats på substrat från extensivt jordbruk som är tillåtet i ekologiskt jordbruk under en övergångsperiod". Ordet "ekologiskt" får inte i denna uppgift, för övrigt på etiketten eller i annonseringen vara mer framträdande än något annat ord i uppgiften.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Med beaktande av rådets förordning (EG, EKSG, Euratom) nr 2458/98 av den 12 november 1998 om ändring av förordning (EEG, Euratom, EKSG) nr 259/68 om fastställande av tjänsteföreskrifter för tjänstemännen i Europeiska gemenskaperna och anställningsvillkor för övriga anställda i dessa gemenskaper samt andra förordningar som skall tillämpas på dessa tjänstemän och anställda vad avser fastställande av löner, pensioner och andra ekonomiska ersättningar i euro (1), bör förordningarna nr 7/66/Euratom och nr 122/66/EEG (2) ändras.
I förordningarna nr 7/66/Euratom, nr 122/66/EEG skall "belgiska franc" ersättas med "euro" och beloppen i belgiska franc ersättas med motsvarande belopp i euroenheter till den av rådet fastställda omräkningskursen.
KOMMISSIONENS FÖRORDNING (EG) nr 2521/98 av den 24 november 1998 om ändring av förordning (EG) nr 577/97 om vissa tillämpningsföreskrifter för rådets förordning (EG) nr 2991/94 om regler för bredbara fetter och rådets förordning (EEG) nr 1898/87 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter
med beaktande av rådets förordning (EG) nr 2991/94 av den 5 december 1994 om regler för bredbara fetter (1), särskilt artikel 8 i denna,
Granskningen av de uppgifter som har lämnats har visat att de toleranser som föreskrivs för kontrollen av fetthalten är alltför snäva. Det har visat sig vara befogat att fördubbla toleranserna för genomsnittet av de prov som tagits samt för de enskilda proven. Under dessa omständigheter kan inte kravet på att resultatet av varje prov skall ligga inom de gränser som fastställs i bilagan till förordning (EG) nr 2991/94 bibehållas. Det bör föreskrivas att de genomsnittliga fetthalter som fastställs skall motsvara dessa gränser.
a) Punkterna 1.b och c skall ersättas med följande:
b) Punkt 2 skall ersättas med följande:
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande (2),
(1) Artikel 19.2, jämförd med artikel 43.1, i stadgan, punkt 8 i protokollet nr 11 om vissa bestämmelser angående Förenade konungariket Storbritannien och Nordirland och punkt 2 i protokollet nr 12 om vissa bestämmelser angående Danmark, skall inte medföra att en icke deltagande medlemsstat får några rättigheter eller skyldigheter.
(4) Enligt artikel 19.1 i stadgan får ECB-rådet fastställa regler för att beräkna och fastställa de minimireserver som krävs.
(7) De sanktioner som föreskrivs vid åsidosättande av skyldigheterna enligt den här förordningen påverkar inte ECBS:s möjligheter att fastställa lämpliga bestämmelser för genomförande och påföljder i förhållande till sina motparter, inbegripet möjligheten att helt eller delvis utestänga ett institut från penningpolitiska transaktioner vid allvarligt åsidosättande av kraven på minimireserver.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
4) reservkvot: den andel i procent av basen för minimireserverna som ECB får fastställa i enlighet med artikel 19.1 i stadgan,
Rätt att undanta institut
Bas för minimireserver
ii) institutets skyldigheter som härrör från poster utanför balansräkningen; i basen skall dock inte ingå
2. För skyldigheter i form av omsättningsbara skuldförbindelser kan ECB som alternativ till bestämmelsen i punkt 1 iii ovan föreskriva att ett instituts skyldigheter gentemot ett annat institut helt eller delvis skall undantas från basen för det fordringsägande institutets minimireserver.
Reservkvoter
Artikel 5
Artikel 6
2. ECB skall ha rätt att med avseende på korrekthet och kvalitet kontrollera den information som instituten tillhandahåller för att visa att de uppfyller kraven på minimireserver. ECB skall underrätta instituten om sitt beslut att verifiera eller inhämta uppgifter.
b) granska institutens räkenskaper och register,
Om ett institut förhindrar inhämtandet och/eller kontrollen av information skall den deltagande medlemsstat i vilken de relevanta lokalerna är belägna ge det bistånd som krävs, däribland säkerställa tillträde till institutets lokaler så att de ovannämnda rättigheterna kan utövas.
Sanktioner vid åsidosättande av kraven
b) Ett åläggande av det berörda institutet att göra en räntelös insättning i ECB eller de nationella centralbankerna till ett belopp av högst tre gånger det belopp varmed institutets reserver understiger kravet på minimireserver. Insättningens löptid skall inte överstiga den period under vilken institutet underlåter att hålla minimireserverna.
Artikel 8
VERKSTÄLLANDE KOMMITTÉNS BESLUT
(SCH/Com-ex (98) 57)
med beaktande av artikel 9 i samma konvention, och av följande skäl:
Enligt kapitel V punkt 1.4 i de gemensamma konsulära anvisningarna "Prövning av övriga för ansökan nödvändiga verifikationer" skall ett enhetligt formulär användas som bevis för att bostad finns.
Följande delar av dokumentet skall således vara enhetliga:
Det enhetliga formuläret skall användas under 1999 i de stater som tillämpar Schengenkonventionen där detta slags bevis föreskrivs i den nationella lagstiftningen.
3. Det enhetliga formulär som skall användas av de avtalsslutande parterna i Schengenavtalet för inbjudningar, åtagandeförklaringar och bevis för att bostad finns skall utarbetas centralt enligt anvisningarna i bilaga A (teknisk beskrivning av säkerhetsdetaljerna) och bilagorna A1 och A2 (modellformulär). De obligatoriska enhetliga uppgifterna i det enhetliga formuläret anges i bilaga B.
6. Dokumentets säkerhetsmässiga utformning skall kontrolleras regelbundet (eventuellt vartannat år). Säkerhetsdetaljerna skall anpassas vartannat år oberoende av de ändringar av allmän karaktär som visar sig nödvändiga om formuläret förfalskas eller om åtgärder för att skydda de tekniska säkerhetsdetaljerna har blivit kända.
KOMMISSIONENS BESLUT av den 25 januari 1999 om förfarandet för bestyrkande av överensstämmelse av byggprodukter enligt artikel 20.2 i rådets direktiv 89/106/EEG beträffande värmeisoleringsprodukter [delgivet med nr K(1999) 115] (Text av betydelse för EES) (1999/91/EG)
med beaktande av rådets direktiv 89/106/EEG av den 21 december 1988 om tillnärmning av medlemsstaternas lagar och andra författningar om byggprodukter (1), ändrat genom direktiv 93/68/EEG (2), särskilt artikel 13.4 i detta, och av följande skäl:
De två förfaranden som avses i artikel 13.3 beskrivs i detalj i bilaga III till direktiv 89/106/EEG. Det är därför nödvändigt att klart ange de metoder genom vilka de två förfarandena skall genomföras, i enlighet med bilaga III, för varje produkt eller produktgrupp, eftersom bilaga III anger att vissa system i första hand skall användas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Förfarandet för bestyrkande av överensstämmelse enligt bilaga III skall anges i uppdragen för harmoniserade standarder.
KOMMISSIONENS DIREKTIV 1999/68/EG
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
1. I kommissionens direktiv 93/78/EEG(2) fastställs genomförandebestämmelser för listor över sorter av prydnadsväxter som förs av leverantörer i enlighet med rådets direktiv 91/682/EEG(3).
4. Ett system för sortbeskrivning finns redan på gemenskapsnivå inom ramen för gemenskapens växtförädlarrätt.
7. Direktiv 93/78/EEG bör upphöra att gälla.
Artikel 1
1. De listor som förs av leverantörer skall innehålla följande:
iii) Sortbeskrivning, åtminstone på grundval av de egenskaper och dessas yttringar såsom de beskrivs i enlighet med bestämmelserna för de ansökningar som skall fyllas i för gemenskapens växtförädlarrätt där denna är tillämplig.
Artikel 3
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv den 31 december 1999. De skall genast underrätta kommissionen om detta.
Artikel 5
om minimikrav för förbättring av säkerhet och hälsa för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär (femtonde särdirektivet enligt artikel 16.1 i direktiv 89/391/EEG)
med beaktande av kommissionens förslag(1), som överlämnats efter samråd med Rådgivande kommittén för arbetarskyddsfrågor och Kommissionen för säkerhet och hälsa för gruvindustrin och andra utvinningsindustrier,
av följande skäl:
3. Målsättningen att förbättra arbetstagarnas säkerhet, arbetshygieniska förhållanden och hälsa på arbetsplatsen får inte underordnas rent ekonomiska överväganden.
6. Detta direktiv bidrar konkret till att förverkliga den inre marknadens sociala dimension.
9. För att fastställa en sammanhängande strategi för explosionsskydd krävs att organisatoriska åtgärder kompletterar de tekniska åtgärderna på arbetsplatsen. I direktiv 89/391/EEG krävs att arbetsgivaren skall ha tillgång till en bedömning av riskerna för arbetstagarnas hälsa och säkerhet på arbetsplatsen. I detta direktiv preciseras detta krav genom att det här föreskrivs att arbetsgivaren skall utarbeta ett explosionsskyddsdokument eller ett antal dokument som uppfyller de minimikrav som fastställs i detta direktiv och som skall hållas aktuellt/a. Detta/dessa explosionsskyddsdokument inbegriper fastställande av farorna, en bedömning av riskerna och fastställande av de särskilda åtgärder som skall vidtas för att säkra arbetstagares hälsa och säkerhet, när de är utsatta för fara orsakad av explosiv atmosfär i enlighet med artikel 9 i direktiv 89/391/EEG. Explosionsskyddsdokument kan vara en del av den riskbedömning i fråga om hälsa och säkerhet i arbetet som krävs enligt artikel 9 i direktiv 89/391/EEG.
12. Samordning bör ske när arbetstagare från flera företag befinner sig på samma arbetsplats.
15. I direktiv 94/9/EG, delas den utrustning och de säkerhetssystem som omfattas in i utrustningsgrupper och -kategorier. I detta direktiv föreskrivs att arbetsgivaren klassificerar områden där explosiv atmosfär kan uppstå i zoner och beslutar vilka grupper och kategorier av utrustning och säkerhetssystem, som skall användas i varje zon.
ALLMÄNNA BESTÄMMELSER
1. I detta direktiv, som är det femtonde särdirektivet i den mening som avses i artikel 16.1 i direktiv 89/391/EEG, fastställs minimikrav för säkerhet och hälsa för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär enligt definitionen i artikel 2.
b) användning av anordningar för förbränning av gasformiga bränslen enligt direktiv 90/396/EEG(7).
e) användning av land-, sjö- och lufttransportmedel på vilka tillämpliga bestämmelser i internationella avtal (till exempel ADNR, ADR, ICAO, IMO, RID) och de gemenskapsdirektiv som ger verkan åt dessa avtal tillämpas. Transportmedel som är avsedda att användas i potentiellt explosiv atmosfär skall inte vara undantagna.
Definition
ARBETSGIVARENS SKYLDIGHETER
I syfte att i enlighet med artikel 6.2 i direktiv 89/391/EEG förhindra och skydda mot explosioner skall arbetsgivaren med hänsyn till verksamhetens art vidta de tekniska och/eller organisatoriska åtgärder som är lämpliga, i prioriterad ordning, och i enlighet med de grundläggande principerna nedan, för att
- begränsa de skadliga effekterna av en explosion, för att säkerställa arbetstagarnas hälsa och säkerhet.
Bedömning av explosionsrisker
- sannolikheten för att tändkällor, inklusive elektrostatiska laddningar, förekommer och att dessa aktiveras och får effekt,
Explosionsriskerna skall bedömas som en helhet.
Allmänna skyldigheter
- lämplig övervakning under arbetstagares närvaro säkerställs i enlighet med riskbedömningen genom användning av lämpliga tekniska medel i en arbetsmiljö där explosiv atmosfär kan uppstå i sådana mängder att arbetstagares säkerhet och hälsa äventyras.
Om arbetstagare från flera företag befinner sig på samma arbetsplats skall varje arbetsgivare ansvara för alla frågor som ligger under hans kontroll.
Områden där explosiv atmosfär kan uppstå
3. Områden där explosiv atmosfär kan uppstå i sådana mängder att arbetstagarnas säkerhet och hälsa äventyras skall vid behov märkas med skyltar vid deras ingångar i enlighet med bilaga III.
Vid uppfyllandet av de skyldigheter som anges i artikel 4 skall arbetsgivaren säkerställa att ett dokument, nedan kallat explosionsskyddsdokumentet, utarbetas och hålls aktuellt.
- att lämpliga åtgärder kommer att vidtas för att uppnå syftet med det här direktivet,
- att arbetsplatsen och arbetsutrustning, inbegripet varningsanordningar, utformas, används och underhålls med vederbörlig hänsyn till säkerhet,
Arbetsgivaren får kombinera befintliga explosionsriskbedömningar, dokument eller andra jämförliga rapporter som upprättas enligt andra gemenskapsrättsakter.
1. Arbetsutrustning, som skall användas i områden där explosiv atmosfär kan uppstå och som redan används eller tillhandahålls i företaget eller i verksamheten för första gången före den 30 juni 2003, skall från och med detta datum uppfylla minimikraven i bilaga II del A, om inga andra gemenskapsdirektiv är tillämpliga eller endast delvis är tillämpliga.
4. Arbetsplatser med områden där explosiv atmosfär kan uppstå som redan tagits i bruk före den 30 juni 2003 skall senast tre år efter den tidpunkten uppfylla minimikraven i detta direktiv.
ÖVRIGA BESTÄMMELSER
Rent tekniska ändringar i bilagorna som föranleds av
skall antas enligt det förfarande som fastställs i artikel 17 i direktiv 89/391/EEG.
Kommissionen skall i en handbok för god praxis av icke bindande natur utarbeta praktiska riktlinjer. Handboken skall behandla de ämnen som anges i artiklarna 3, 4, 5, 6, 7 och 8, bilaga I och bilaga II del A.
Artikel 12
Artikel 13
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 14
om anpassning till den tekniska utvecklingen av Europaparlamentets och rådets direktiv 96/79/EG om skydd av förare och passagerare i motorfordon vid frontalkollision
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
3. De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från den kommitté för anpassning till teknisk utveckling som inrättats i enlighet med direktiv 70/156/EEG.
Bilaga II till direktiv 96/79/EG skall ändras i enlighet till bilagan till detta direktiv.
- vägra EG-typgodkännande för en ny fordonstyp, eller
2. Från och med den 1 april 2001 får medlemsstaterna inte längre bevilja EG-typgodkännande för en fordonstyp i enlighet med artikel 4 i direktiv 70/156/EEG om den inte uppfyller kraven i direktiv 96/79/EG, i dess lydelse efter ändringar genom det här direktivet.
När medlemsstaterna antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
INTERINSTITUTIONELLT AVTAL
med hänvisning till Europaparlamentets resolution av den 7 oktober 1998 om oberoende, roll och ställning för enheten för samordning av bedrägeribekämpning (Uclaf)(1),
och av följande skäl: (1) Europaparlamentets och rådets förordning (EG) nr 1073/1999(3) och rådets förordning (Euratom) nr 1074/1999(4) om utredningar som utförs av Europeiska byrån för bedrägeribekämpning innehåller bestämmelser om att byrån skall inleda och utföra administrativa utredningar inom de institutioner, organ och byråer som inrättats genom EG-fördraget och Euratomfördraget eller på grundval av dessa fördrag.
(4) Alla institutioner, organ och byråer bör i kraft av sin administrativa självständighet ge byrån i uppdrag att inom dessa utföra administrativa utredningar för att efterforska sådana omständigheter av allvarlig art som har samband med tjänsteutövningen och som skulle kunna utgöra sådana brister när det gäller att uppfylla de skyldigheter som åligger tjänstemän och anställda i gemenskaperna som avses i artiklarna 11, 12 andra och tredje styckena, 13, 14, 16 och 17 första stycket i tjänsteföreskrifterna för tjänstemän och anställningsvillkoren för övriga anställda i Europeiska gemenskaperna (nedan kallade "Tjänsteföreskrifterna"), brister som kan skada dessa gemenskapers intressen och som kan leda till disciplinära åtgärder och, i förekommande fall, straffrättsliga åtgärder, eller ett allvarligt fel i tjänsten enligt artikel 22 i tjänsteföreskrifterna eller en bristande uppfyllelse av motsvarande skyldigheter som åvilar ledamöter, chefer eller medlemmar av personalen vid gemenskapens institutioner, organ eller byråer, som inte omfattas av tjänsteföreskrifterna.
(7) De praktiska villkoren bör fastställas för hur institutionernas och organens ledamöter, byråernas chefer och tjänstemännen och de anställda inom dessa skall samarbeta för att de interna utredningarna skall kunna utföras väl, i avvaktan på att tjänsteföreskrifterna ändras,
INGÅTT FÖLJANDE AVTAL:
- efterforska sådana omständigheter av allvarlig art som har samband med tjänsteutövningen och som skulle kunna utgöra brister när det gäller att uppfylla de skyldigheter som åligger tjänstemän och anställda i gemenskaperna, brister som skulle kunna leda till disciplinära åtgärder och, i förekommande fall, straffrättsliga åtgärder, eller en bristande uppfyllelse av motsvarande skyldigheter, som åvilar ledamöter, chefer eller medlemmar av personalen, som inte omfattas av tjänsteföreskrifterna.
2. Institutionerna åtar sig att inrätta en sådan ordning och att göra den omedelbart tillämplig genom att anta ett internt beslut enligt den modell som bifogas detta avtal och att inte avvika från modellbeslutet annat än om särskilda förhållanden inom den egna institutionen gör detta nödvändigt av tekniska skäl.
Detta avtal får bara ändras efter uttryckligt medgivande från de undertecknande institutionerna.
RÅDETS FÖRORDNING (EG) nr 150/1999 av den 19 januari 1999 om ändring av förordning (EEG) nr 2262/84 om särskilda bestämmelser för olivolja
med beaktande av kommissionens förslag (1),
Det har fattats beslut om en treårig övergångsperiod från och med regleringsåret 1998/1999 med hänvisning till reformen av den gemensamma organisationen av marknaden för olivolja. De arbetsuppgifter som vanligtvis åläggs organen måste genomföras under övergångsperioden och under det första regleringsåret efter denna period. Det är därför lämpligt att föreskriva att gemenskapen delar organens kostnader för denna period för att se till att de fungerar effektivt och kontinuerligt inom ramen för det administrativa självstyre som föreskrivs i förordning (EEG) nr 2262/84.
I artikel 1.5 i förordning (EEG) nr 2262/84 skall de två sista styckena ersättas med följande:
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EEG) nr 1898/87 av den 2 juli 1987 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter (2), senast ändrad genom förordning (EG) nr 222/98 (3), särskilt artikel 4.2 i denna, och
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl: I artikel 2.2 a första strecksatsen i kommissionens förordning (EG) nr 785/95 av den 6 april 1995 om tillämpningsföreskrifter för rådets förordning (EG) nr 603/95 (3), senast ändrad genom förordning (EG) nr 1794/97 (4), föreskrivs att dehydratisering av färskt foder skall ske med hjälp av torkar som håller en temperatur på minst 93 °C i början av processen.
På de flesta företag äger bearbetning av foder rum vid hög temperatur. Det är därför lämpligt att föreskriva att de anläggningar som fortfarande håller en temperatur på 93 °C i början av processen inom rimlig tid justeras för att vara anpassade till torkning av foder vid hög temperatur.
I artikel 15 b i ovannämnda förordning (EG) nr 785/95 föreskrivs att medlemsstaterna skall meddela kommissionen de arealer och kvantiteter som berörs av kontrakt och leveransdeklarationer. Erfarenheten har visat att denna rapportering är en källa till motsägelsefulla och otillfredsställande uppgifter. Den bör därför avskaffas.
Artikel 1
Artikel 2
Artikel 3
av den 7 april 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Det är följaktligen nödvändigt att omarbeta nämnda förordning och låta bilaga I till förordning nr 920/89 utgå. För att förbättra överskådligheten på världsmarknaden bör därför de normer för morötter beaktas som rekommenderats av den arbetsgrupp för standardisering av lättfördärvliga livsmedel samt för kvalitetsförbättring som inrättats vid Förenta nationernas ekonomiska kommission för Europa (ECE/FN).
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för färsk frukt och färska grönsaker.
Handelsnormerna för morötter som omfattas av KN-nummer 0706 10 00 anges i bilagan.
- uppvisa en viss bristande färskhet och saftspändhet, och
Förordning (EEG) nr 920/89 ändras på följande sätt:
Artikel 3
av den 26 maj 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1095/96 av den 18 juni 1996 om genomförande av medgivandena i lista CXL som fastställs sedan förhandlingarna enligt GATT artikel XXIV.6 avslutats(5), särskilt artikel 1.1 i denna, och av följande skäl:
(3) Erfarenheten visar att begränsningen av importen kan ge upphov till ansökningar om importlicens i spekulativt syfte. För att de planerade åtgärderna skall fungera som avsett bör huvuddelen av de tillgängliga kvantiteterna förbehållas s.k. traditionella importörer av tjurar, kor och kvigor av vissa alp- och bergraser. I vissa fall finns det en risk för att administrativa felaktigheter som begåtts av den nationella behöriga myndigheten begränsar importörernas tillträde till denna del av kovten. Bestämmelser bör fastställas för att korrigera eventuella felaktigheter.
(6) För att undvika spekulationer bör s.k. traditionella importörer som inte längre var verksamma inom nötköttssektorn den 1 juni före importåret i fråga inte vara berättigade till kvoten.
(9) I artikel 82 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(10), senast ändrad genom förordning (EG) nr 955/1999(11), fastställs att varor som övergår till fri omsättning till en nedsatt tullsats med hänvisning till deras särskilda slutanvändning skall stå under tullens övervakning. En kontroll skall utföras för att säkerställa att de importerade djuren inte slaktas under en viss period. En säkerhet bör ställas för att garantera att dessa djur inte slaktas, vilken skall täcka skillnaden mellan tullarna enligt den gemensamma tulltaxan (GTT) och de nedsatta tullar som gäller den dag då djuren i fråga övergår till fri omsättning.
(12) För tydlighetens skull bör bestämmelserna i artiklarna 2.1 a och 8 c i förordning (EG) nr 1143/98 rättas till.
Artikel 1
2. Vid tillämpningen av denna förordning skall de djur som avses i punkt 1 inte anses vara slaktdjur om de inte slaktas inom fyra månader från det att deklarationen om övergång till fri omsättning har godkänts.
- För tjurar: Stamtavla.
1. De två kvoter som avses i artikel 1.1 skall delas i två delar om 80 %, dvs. 4000 djur, respektive 20 %, dvs. 1000 djur.
b) Den andra delen av kvoten om 20 % förbehålls sökande som kan styrka att de under de tolv månader som föregick importåret i fråga har importerat minst 15 levande nötkreatur som omfattas av KN-nummer 0102 från tredje land.
3. På grundval av ansökningarna om importtillstånd skall fördelningen av den andra delen ske i proportion till de kvantiteter som de importörer som nämns i punkt 1 b har ansökt om.
- får inte avse mer än 50 djur.
Medlemsstaterna får godta kopior av dessa dokument, som vederbörligen bestyrkts av den utfärdande myndigheten, om den sökande till den behöriga myndighetens tillfredsställelse kan visa att det varit omöjligt för honom att skaffa fram originaldokumentet.
2. Ett företag som uppstått genom en sammanslagning av företag som vart och ett enligt artikel 2.2 var berättigat att delta, skall ha samma rättigheter som de ursprungliga företaget.
2. Endast en ansökan per kvot får lämnas in av en och samme aktör och den får avse endast en av delarna av en enskild tullkvot.
4. Efter kontroll av dokumenten skall medlemsstaterna senast den tionde arbetsdagen efter det att perioden för inlämnande av ansökningar löpt ut för varje löpnummer anmäla följande till kommissionen:
5. Samtliga sådana anmälningar, även anmälningar om att inga ansökningar tagits emot, skall göras via telefax, och utformas enligt förlagorna i bilagorna II och III i de fall då ansökningar har lämnats in.
2. Om de kvantiteter för vilka ansökningar enligt artikel 4.4 andra strecksatsen har lämnats in överstiger de disponibla kvantiteterna, skall kommissionen minska kvantiteterna i ansökningarna med en enhetlig procentsats.
1. För att de tilldelade kvantiteterna skall få importeras, krävs det att en eller flera importlicenser uppvisas.
4. Licenserna skall vara giltiga i 90 dagar från och med utfärdandedagen enligt artikel 21.1 i förordning (EEG) nr 3719/88. Licenserna får dock endast utfärdas från och med den 1 juli varje importår och skall upphöra att gälla senast den 30 juni.
7. Genom undantag från artikel 9.1 i förordning (EEG) nr 3719/88 får importlicenser, som utfärdats i enlighet med denna förordning, inte överlåtas och de kan endast ge tillgång till tullkvoter om de är utfärdade i samma namn som de deklarationer om övergång till fri omsättning som åtföljer dem.
1. Kontrollen av att de importerade djuren inte slaktas under en period på fyra månader från dagen för övergång till fri omsättning skall ske i överensstämmelse med bestämmelserna i artikel 82 i förordning (EEG) nr 2913/92.
a) inte har slaktats före utgången av perioden på fyra månader från dagen för deras övergång till fri omsättning,
a) I fält 8, uppgift om ursprungslandet. Licensen innebär skyldighet att importera från det angivna landet.
- Bergrassen (Verordening (EG) nr. 1081/1999), invoerjaar: ...
2. I detta syfte skall medlemsstaterna senast den 22 mars under importåret för varje löpnummer till kommissionen anmäla de kvantiteter för vilka det inte har ansökts om importlicens.
Oavsett om en ansökan avser en kvantitet som överstiger denna kvantitet, skall endast den kvantiteten beaktas.
6. Samtliga ansökningar om importtillstånd skall vara de behöriga myndigheterna till handa senast fem arbetsdagar efter dagen för ikraftträdandet för det kommissionsbeslut som avses i punkt 3.
Artikel 10
Förordning (EG) nr 1143/98 ändras på följande sätt:
3) Artikel 8 c skall ersättas med följande: "c) I fält 20, en av följande uppgifter:
Artikel 12
av den 28 maj 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(2) Mot bakgrund av de tekniska arrangemang som överenskommits mellan de ryska myndigheterna och kommissionen, efter det att förordningen trädde i kraft, bör de allmänna tillämpningsföreskrifterna ändras på ett antal punkter, särskilt när det gäller bestämmelserna för hur mottagarlandet övertar produkterna och kommissionens förfarande för kontroll av hur leveranserna genomförs.
(5) Det är lämpligt att föreskriva omedelbar tillämpning av de ändringar som följer av de tekniska arrangemang som överenskommits med de ryska myndigheterna beträffande bestämmelserna för produktövertag och beträffande vissa bestämmelser för kontroll i samband med produktuttag och för frisläppande av säkerheter till förmån för aktörerna.
Artikel 1
8) I artikel 5.1 g skall punkt 4 utgå.
Varorna kan lastas så snart interventionsorganet erhållit bevis för att det har ställts en leveranssäkerhet i enlighet med punkt 4."
17) I artikel 9.1 skall andra stycket ersättas med följande: "För de leveranser som avser produktion av helt slipat ris eller anskaffande av griskött på gemenskapsmarknaden skall det uttagsintyg som utfärdas i enlighet med bilaga V och som undertecknas av det organ som ansvarar för utfärdandet av detsamma utgöra bevis för att produkten uppfyller de krav som fastställts för leveransen."
a) i de fall då artikel 2.1 b tillämpas, åtföljas av
- intyg om överensstämmelse vid bestämmelseorten i enlighet med artikel 9.7,
3. Vid leverans enligt artikel 2.1 a eller b skall leveranskostnaderna betalas för den kvantitet som anges i övertagandeintyget som skall utfärdas av det kontrollorgan som kommissionen utser och som skall viseras av de företrädare för mottagarlandet som anges i förordningen om öppnande av ett anbudsförfarande. Övertagandeintyget skall utfärdas i enlighet med bilaga I.
6. Om övertagandet på bestämmelseorten fördröjs på grund av omständigheter som inte kan påverkas av kontraktsinnehavaren, skall mottagarlandet ersätta anbudsgivaren för dennes extrakostnader på grundval av bestyrkande handlingar.
3. I de fall då det för export av en produkt krävs att exportlicensansökan uppvisas skall denna åtföljas av ett bevis för att sökanden är innehavare av ett kontrakt avseende leveranser enligt förordning (EG) nr 2802/98. Beviset skall utgöras av en kopia av det meddelande om tilldelning av leveranskontrakt som avses i artikel 6.3.
28) Bilaga B till den här förordningen skall införas som bilaga VII.
KOMMISSIONENS FÖRORDNING (EG) nr 1245/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
(1) Enligt direktiv 70/524/EEG får nya fodertillsatser och nya användningsområden för fodertillsatser tillåtas mot bakgrund av den vetenskapliga och tekniska utvecklingen.
(4) Nya fodertillsatser och nya användningsområden för fodertillsatser får tillåtas tillfälligt under förutsättning att de halter som tillåts i foder inte medför fara för miljön eller människors eller djurs hälsa och inte är till skada för konsumenterna genom att djurproduktens egenskaper förändras, att tillsatsens närvaro i foder kan kontrolleras och att närvaron av fodertillsatsen enligt tillgängliga forskningsresultat sannolikt har en gynnsam effekt på foderegenskaperna eller på djuruppfödningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
om finansiering av den gemensamma jordbrukspolitiken
med beaktande av kommissionens förslag(1),
med beaktande av revisionsrättens yttrande(4), och
3. Fondens utvecklingssektion bör finansiera utgifter för vissa åtgärder för landsbygdsutveckling i regioner som utvecklas långsammare samt för gemenskapens initiativ för landsbygdsutveckling.
6. I samband med granskning och godkännande av räkenskaperna kan kommissionen inom skälig tid besluta om de totala utgifter som skall införas i garantisektionen i räkenskaperna, endast om den får tillfredsställande garantier för att de nationella kontrollerna är tillräckliga och ger insyn i verksamheten, och att utbetalningsställena försäkrar sig om att de utbetalningar som de gör är lagliga och riktiga. Bestämmelser bör därför antas för ackreditering av utbetalningsställena från medlemsstaternas sida. För att säkerställa konsekvens i den standard som krävs för ackreditering i medlemsstaterna skall kommissionen dra upp riktlinjer avseende de kriterier som skall tillämpas. Det bör därför föreskrivas att enbart utbetalningar som görs av de utbetalningsställen som är ackrediterade av medlemsstaterna får verkställas. För alt säkerställa insyn i de nationella kontrollsystemen, särskilt såvitt avser förfarandet för godkännande, bemyndigande och utbetalning, bär i förekommande fall antalet myndigheter och organ som anförtros detta ansvar begränsas med hänsyn till varje medlemsstats konstitutionella bestämmelser.
9. Det är lämpligt att föreskriva två olika slag av beslut, ett som avser granskning och godkännande av räkenskaperna för fondens garantisektion, och ett som lägger fast vilka slutsatser, inbegripet finansiella rättelser, som kan dras av resultaten av granskningen huruvida utgifterna överensstämmer med gemenskapsbestämmelserna.
12. Gemenskapens utgifter måste noga övervakas. Utöver den övervakning som medlemsstaterna utför på eget initiativ och som förblir av största vikt, bör bestämmelser fastställas så att kommissionens tjänstemän kan genomföra kontroller och ha rätt att begära hjälp från medlemsstaterna.
15. För att förenkla den finansiella förvaltningen är det önskvärt att närma fondens finansieringsperiod till budgetåret såsom det anges i artikel 272.1 i fördraget. För att detta skall kunna göras måste det finnas en klar bild av vilka medel som finns tillgängliga vid utgången av budgetåret i fråga. Det bör därför föreskrivas att kommissionen får nödvändig befogenhet att anpassa fondens finansieringsperiod om tillräckliga budgetmedel finns tillgängliga.
Den skall bestå av följande två sektioner:
2. Garantisektionen skall finansiera
c) åtgärder för landsbygdsutveckling utanför mål 1-program med undantag av gemenskapsinitiativet för landsbygdsutveckling,
3. Utveckingssektionen skall finansieras sådana åtgärder för landsbygdsutveckling som inte omfattas av punkt 2 c.
1. Bidrag vid export till tredje land, beviljade i enlighet med gemenskapsbestämmelserna inom ramen för den gemensamma organisationen av jordbruksmarknaderna skall finansieras enligt artikel 1.2 a.
Artikel 3
3. Informationsåtgärder och utvärderingsåtgärder som vidtas enligt gemenskapsbestämmelser skall finansieras enligt artikel 1.2 e.
1. Varje medlemsstat skall underrätta kommissionen om följande:
2. Utbetalningsställena skall vara medlemsstaternas myndigheter och organ som, såvitt avser de betalningar som skall göras inom deras områden skall ge tillräckliga garantier för att
c) nödvändiga handlingar ges in inom den tid och i den form som föreskrivs i gemenskapsbestämmelserna.
5. Varje medlemsstat skall, med beaktande av landets konstitutionella bestämmelser och institutionella struktur, begränsa antalet ackrediterade utbetalningsställen till minsta möjliga antal för att de utgifter som avses i artiklarna 2 och 3 skall kunna betalas under tillfredsställande förvaltnings- och redovisningsförhållanden.
b) Förvaltnings- och redovisningsförhållanden samt interna kontrollförhållanden under vilka betalningar skall göras i samband med genomförandet av gemenskapsbestämmelserna inom ramen för den gemensamma jordbrukspolitiken.
7. Om ett eller flera av villkoren för ackrediteringen inte har uppfyllts eller inte längre uppfylls av ett godkänt utbetalningsställe skall ackrediteringen återkallas, såvida inte utbetalningsstället genomför nödvändiga anpassningar inom den tid som bestäms utifrån hur allvarligt problemet är. Den berörda medlemsstaten skall underrätta kommissionen om detta.
1. De ekonomiska resurser som krävs för att täcka de utgifter som avses i artiklarna 2 och 3 skall göras tillgängliga för medlemsstaterna av kommissionen genom förskott på utgifter som verkställts under en referensperiod.
3. Tillämpningsföreskrifterna för denna artikel skall antas i enlighet med förfarandet i artikel 13.
a) En redovisning av utgifterna och en bedömning av finansieringsbehoven.
Artikel 7
Utgifterna för oktober skall hänföras till oktober om de verkställs mellan den 1 och den 15 oktober och till november om de verkställs mellan den 16 och den 31 oktober. Förskottsbetalningar skall göras till medlemsstaten senast den tredje arbetsdagen i den andra månaden efter den månad då utgifterna verkställs.
Beslutet att granska och godkänna räkenskaperna skall omfatta den överlämnade redovisningens fullständighet, exakthet och sanningsenlighet. Beslutet skall inte påverkar antagandet av ett senare beslut i enlighet med punkt 4.
Om ingen överenskommelse nås får medlemsstaten begära att ett förfarande inleds i syfte att medla mellan deras respektive ståndpunkter inom en tid av fyra månader; resultaten härav skall anges i en rapport, som skall överlämnas till och granskas av kommissionen innan ett beslut om att vägra finansiering fattas.
a) De utgifter som avses i artikel 2 och som verkställts före de tjugofyra månader som föregick kommissionens skriftliga meddelande till den berörda medlemsstaten om resultaten av kontrollerna.
a) av oegentligheter enligt artikel 8.2,
Artikel 8
b) förhindra och ingripa mot oegentligheter,
2. Om en fullständigt indrivning inte kan åstadkommas skall de ekonomiska följderna av oegentligheter eller försumlighet bäras av gemenskapen, med undantag för följderna av sådana oegentligheter eller sådan försumlighet som kan tillskrivas medlemsstaternas myndigheter eller andra organ.
Artikel 9
2. Utan att det påverkar den kontroll som medlemsstaterna utför i enlighet med nationella bestämmelser i lagar och andra författningar och utan att det påverkar tillämpningen av bestämmelserna i artikel 248 i fördraget eller sådana kontroller som företas med stöd av artikel 279 c i fördraget skall företrädare som kommissionen utsett att genomföra kontroller på plats ha tillgång till alla böcker och andra handlingar, inbegripet uppgifter som upprättas eller lagras i elektronisk form, avseende utgifter som finansieras av fonden.
b) om de erforderliga underlagen finns och om dessa överensstämmer med de transaktioner som finansieras av fonden,
På begäran av kommissionen och med medlemsstatens samtycke skall kontroller eller utredningar beträffande de transaktioner som avses i denna förordning utföras av den medlemsstatens behöriga myndigheter. Tjänstemän från kommissionen får också delta.
Artikel 10
Kommittén för Europeiska utvecklings- och garantifonden för jordbruket (nedan kallad fondkommittén) skall bistå kommissionen med förvaltningen av fonden i enlighet med bestämmelserna i artiklarna 12-15.
Artikel 13
3. a) Kommissionens beslut skall ha omedelbar verkan.
- Rådet får inom den tidsfrist som anges i föregående strecksats fatta ett annat beslut med kvalificerad majoritet.
a) i samtliga fall där det är föreskrivet att den skall höras,
2. Fondkommittén får undersöka alla andra frågor som dess ordförande, antingen på eget initiativ eller på begäran av en företrädare för en medlemsstat, har hänskjutit till den.
Ordföranden skall sammankalla fondkommittén.
Artikel 16
Artikel 17
De åtgärder som krävs för att underlätta övergången från bestämmelserna i förordning (EEG) nr 729/70 till bestämmelserna i den här förordningen skall antas enligt förfarandet i artikel 13.
Artikel 20
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
1. Enligt bestämmelserna i direktiv 70/524/EEG får nya fodertillsatser och nya användningsområden för fodertillsatser godkännas om detta verkar rimligt mot bakgrund av den vetenskapliga och tekniska utvecklingen.
4. Bestämmelserna i rådets direktiv 89/391/EEG av den 12 juni 1989(5) om åtgärder för att främja förbättringar av arbetstagarnas säkerhet och hälsa i arbetet och andra enskilda direktiv, särskilt rådets direktiv 90/679/EEG av den 26 november 1990(6) om skydd för arbetstagare mot risker vid exponering för biologiska agenser i arbetet, senast ändrat genom direktiv 97/65/EG(7), kan till fullo tillämpas när det gäller arbetstagare som handlar fodertillsatser.
7. De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga foderkommittén.
De preparat av typen enzymer som förtecknas i bilaga I till denna förordning får godkännas som fodertillsatser i enlighet med direktiv 70/524/EEG på de villkor som anges i nämnda bilaga.
Artikel 3
av den 9 november 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
1. För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
4. Det är lämpligt att bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning fortfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3), senast ändrad genom rådets och Europaparlamentets förordning (EG) nr 955/1999(4), under en period av tre månader.
Artikel 1
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställas i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
KOMMISSIONENS FÖRORDNING (EG) nr 2562/1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
1. På grund av den risk som dåliga plagiat av zootekniska tillsatser inom gemenskapen utgör för människors och djurs hälsa, skall enligt direktiv 70/524/EEG, ändrat genom rådets direktiv 96/51/EG(3), godkännandet av vissa grupper av tillsatser knytas till den som är ansvarig för avyttringen.
4. För de tillsatser som förtecknas i bilagorna till den här förordningen har den som är ansvarig för den dokumentation utifrån vilken det tidigare godkännandet meddelades eller dennes efterträdare lämnat in nya ansökningar om godkännande. Ansökningarna för dessa tillsatser åtföljdes av erforderlig monografi och identitetsbeskrivning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EEG) nr 2921/90 om beviljande av stöd för framställningen av kasein och kaseinater av skummjölk
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), särskilt artikel 15 i denna, och
2. Förvaltningskommittén för mjölk och mjölkprodukter har inte avgivit något yttrande inom den tid som dess ordförande har bestämt.
Artikel 1 i förordning (EEG) nr 2921/90 skall ändras på följande sätt:
c) kasein: den, i vatten olösliga, tvättade och torkade produkt som erhålls från råkasein eller skummjölk genom utfällning medelst syrning med bakteriekultur eller tillsats av syra, löpe eller andra mjölkkoagulerande enzymer, utan hänsyn till eventuell föregående jonbytes- eller koncentreringsbehandling,
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
om allmänna principer för ersättning till uppgiftslämnare och infiltratörer
Arbetsgruppen för narkotikafrågor åtog sig detta ämne under det tyska ordförandeskapet och den har granskat rättsläget och rättspraxis i var och en a
om ändring av kommissionens beslut 93/436/EEG om särskilda villkor för import av fiskeriprodukter med ursprung i Chile
(2000/61/EG)
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktionen och marknadsföringen av fiskeriprodukter(1), senast ändrat genom rådets direktiv 97/79/EG(2), särskilt artikel 11 i detta, och
4. De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Bilaga A till beslut 93/436/EEG skall ersättas med bilagan till det här beslutet.
Kommissionens beslut
[delgivet med nr K(2000) 656]
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av kommissionens förordning (EEG) nr 3600/92 av den 11 december 1992 om närmare bestämmelser för genomförandet av den första etappen i det arbetsprogram som avses i artikel 8.2 i rådets direktiv 91/414/EEG om utsläppande av växtskyddsprodukter på marknaden(3), senast ändrad genom förordning (EG) nr 1199/97(4), särskilt artikel 7.3a led b i denna, och
(2) Monolinuron är ett av de 90 verksamma ämnen som omfattas av den första etappen av det arbetsprogram som fastställs i artikel 8.2 i rådets direktiv 91/414/EEG.
(5) Det framgår av de utvärderingar som gjorts att de uppgifter som lämnats inte visar att växtskyddsmedel som innehåller det verksamma ämnet i fråga uppfyller kraven enligt artikel 5.1 a, 5.1 b i direktiv 91/414/EEG.
(8) Ett tidsbegränsat anstånd skall fastställas i enlighet med artikel 4.6 i direktiv 91/414/EEG under vilken tid kvarvarande lager får omhändertas, lagras, släppas ut på marknaden och användas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
2. inga tillstånd för växtskyddsmedel som innehåller monolinuron beviljas eller förnyas enligt undantaget i artikel 8.2 i direktiv 91/414/EEG från och med dagen för anmälan av detta beslut.
Artikel 4
av den 25 juli 2000
(Text av betydelse för EES)
med beaktande av rådets direktiv 90/539/EEG av den 15 oktober 1990 om djurhälsovillkor för handel inom, gemenskapen med och för import från tredje land av fjäderfä och kläckningsägg(1), senast ändrat genom rådets direktiv 1999/90/EG(2), särskilt artikel 23.1, artikel 24, artikel 26.2 samt artiklarna 27a och 34 i detta,
(1) I kommissionens beslut 96/482/EG(5), senast ändrat genom beslut 1999/549/EG(6), fastställs djurhälsovillkor och veterinärintyg för import från tredje land av fjäderfä och kläckägg med undantag av strutsfåglar och ägg från strutsfåglar, inbegripet djurhälsoåtgärder som skall vidtas efter sådan import.
(4) Det är nödvändigt att den behöriga myndigheten i den avsändande medlemsstaten via Animo-systemet informerar den behöriga myndigheten på de dagsgamla kycklingarnas slutliga destinationsort om de djurhälsokrav avseende isoleringstid som skall tillämpas i dessa fall.
Artikel 1
Följande skall läggas till i artikel 3.1 i beslut 96/482/EG:"Om dagsgamla kycklingar inte föds upp i den medlemsstat till vilken kläckäggen importerats skall de direkt transporteras till och förvaras på den anläggning som avses i punkt 9.2 i förlaga 2 till hälsointyg i bilaga IV till rådets direktiv 90/539/EEG under åtminstone tre veckor från kläckningsdagen."
Artikel 4
av den 26 juli 2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) Enligt direktiv 95/46/EG skall bedömningen av skyddsnivån ske på grundval av alla de förhållanden som har samband med en överföring eller en grupp överföringar av uppgifter och vissa omständigheter skall särskilt beaktas. Arbetsgruppen för skydd av enskilda med avseende på behandling av personuppgifter som inrättats genom det direktivet(2) har utfärdat riktlinjer för hur sådana beddömningar skall göras(3).
(6) Områden och/eller databehandling som inte lyder under någon av de myndigheter i Förenta staterna som anges i bilaga VII till detta beslut bör inte omfattas av beslutet.
(9) Systemet med safe harbor sådant det utformats enligt principerna och FoS kan behöva ses över i ljuset av erfarenheter från utveckling på integritetsskyddets område under förhållanden då tekniken ständigt gör det lättare att överföra och behandla personuppgifter och i ljuset av rapporter om genomförande av berörda tillsynsmyndigheter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) En översikt över genomförandet av safe harbor, bilaga III.
d) En skrivelse från Förenta staternas transportministerium, bilaga VI.
b) denna organisation omfattas av de lagstadgade befogenheter som tillkommer någon av de myndigheter i Förenta staterna som anges i bilaga VII till detta beslut och som är bemyndigade att handlägga klagomål och ge upprättelse vid användning av illojala och bedrägliga metoder och att utverka skadestånd åt enskilda, oberoende av deras bosättningsland eller nationalitet, om principerna inte följs i överensstämmelse med FoS.
Detta beslut gäller endast frågan om den skyddsnivå är adekvat som enligt principerna och FoS erbjuds i Förenta staterna, i förhållande till de krav som ställs i artikel 25.1 i direktiv 95/46/EG, och det påverkar inte tillämpningen av andra bestämmelser i det direktivet som gäller behandling av personuppgifter inom medlemsstaterna, särskilt artikel 4 i direktivet.
a) den myndighet i Förenta staterna som avses i bilaga VII till detta beslut eller en sådan oberoende instans för handläggning av klagomål som avses under a i avsnittet om kontroll av efterlevnaden i bilaga I till detta beslut, har funnit att organisationen agerar i strid med principerna tillämpade i överensstämmelse med FoS, eller
2. Medlemsstaterna skall utan dröjsmål underrätta kommissionen om åtgärder som vidtagits med stöd av punkt 1.
Artikel 4
Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att följa detta beslut senast nittio dagar efter det att beslutet har delgivits medlemsstaterna.
Kommissionens beslut
[delgivet med nr K(2000) 2285]
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I direktiv 91/414/EEG (nedan kallat direktivet) föreskrivs att en gemenskapsförteckning skall upprättas över verksamma ämnen som får användas i växtskyddsmedel.
(4) Företaget BASF AG lämnade den 28 februari 2000 in en akt med dokumentation för det verksamma ämnet BAS500F (pyraclostrobin) till de tyska myndigheterna.
(7) Akterna för RH-7281 (zoxamid), B-41; E-187 (milbemectin), BAS500F (pyraclostrobin) och AEF130360 (foramsulfuron) remitterades till Ständiga kommittén för växtskydd den 31 maj 2000.
(10) Ett sådant beslut hindrar inte att ytterligare faktauppgifter och upplysningar kan komma att begäras in från de ansökande företagen för att klargöra vissa punkter i den dokumentation som lagts fram. Då den rapporterande medlemsstaten begär in sådana upplysningar som är nödvändiga för att klargöra innehållet i dokumentationen skall detta inte påverka tidsfristen för inlämnande av den rapport som avses i skäl 12.
(13) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för växtskydd.
Med hänsyn till de föreslagna användningsområdena uppfyller följande akter med dokumentation i princip de krav beträffande uppgifter och upplysningar som anges i bilaga II och, vad beträffar minst ett växtskyddsmedel som innehåller det verksamma ämnet i fråga, i bilaga III till direktivet:
3. Den dokumentation som lämnats in av BASF AG till kommissionen och medlemsstaterna beträffande införandet av BAS500F (pyraclostrobin) som ett verksamt ämne i bilaga I till direktiv 91/414/EEG, och som överlämnades till Ständiga kommittén för växtskydd den 31 maj 2000.
av den 20 mars 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 95 i detta,
i enlighet med det förfarande som anges i artikel 251 i fördraget(2) och
(2) Skillnader mellan medlemsstaternas lagar och andra författningar om märkning av livsmedel kan hämma den fria rörligheten av dessa varor och kan leda till ojämlika konkurrensvillkor.
(5) Specialregler som tillämpas vertikalt endast på vissa livsmedel bör fastställas inom ramen för de bestämmelser som behandlar dessa varor.
(8) Detaljerad märkning för att ange produktens exakta art och beskaffenhet gör det möjligt för konsumenten att göra sitt val med full sakkännedom och är det lämpligaste eftersom det medför minsta möjliga hinder för den fria handeln.
(11) Medlemsstaterna bör vidare, om det saknas specialregler inom gemenskapen, behålla rätten att fastställa vissa nationella bestämmelser som komplement till de allmänna bestämmelserna i detta direktiv, dock bör dessa bestämmelser vara underkastade en gemenskapsprocedur.
(14) Reglerna för märkning bör också förbjuda användning av information som skulle kunna vilseleda köparen eller som tillskriver livsmedel hälsobringande egenskaper; detta förbud bör för att vara verksamt gälla också presentation av och reklam för livsmedel.
(17) För att förenkla och påskynda förfarandet bör kommissionen anförtros uppgiften att besluta om verkställighetsåtgärder av teknisk natur.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) märkning: varje ord, uppgift, varumärke, märkesnamn, illustration eller symbol i samband med livsmedel som anbringas på förpackning, dokument, meddelande, etikett, ring eller hylsa som medföljer eller avser sådant livsmedel,
1. Märkningen och dess närmare utformning får inte
ii) genom att tillskriva livsmedlet verkningar eller egenskaper som det inte har,
2. Rådet skall på det sätt som anges i artikel 95 i fördraget, upprätta en icke uttömmande förteckning över sådana påståenden som avses i punkt 1 och vilkas användning i alla händelser måste förbjudas eller begränsas.
b) reklam.
1. Det namn under vilket varan säljs.
4. Nettokvantitet i fråga om färdigförpackade livsmedel.
7. Förpackarens eller tillverkarens namn eller firma samt adress eller uppgift om säljare som är etablerad inom gemenskapen.
8. Uppgift om den plats där livsmedlet är producerat eller varifrån det kommer i fall då underlåtenhet att lämna sådana uppgifter kan vilseleda konsumenten i fråga om livsmedlets rätta ursprung eller härkomst.
2. Utan hinder av punkt 1 får medlemsstaterna behålla nationella bestämmelser som föreskriver att tillverkaren eller förpackaren skall anges, såvitt avser deras nationella livsmedelsproduktion.
1. Gemenskapsbestämmelser som gäller endast för vissa livsmedel och inte livsmedel i allmänhet får i särskilda fall avvika från de krav som fastställs i artikel 3.1 punkterna 2 och 5, under förutsättning att detta inte leder till att köparen blir bristfälligt informerad.
1. Det namn under vilket ett livsmedel säljs skall vara det namn som förbehållits livsmedlet i gemenskapens bestämmelser för livsmedlet.
b) Det skall också vara tillåtet att i den medlemsstat där livsmedlet saluförs använda det namn under vilken produkten tillverkas och saluförs i den medlemsstat där tillverkningen sker.
2. Inget varumärke, märkesnamn eller fantasinamn får användas i stället för det namn under vilket varan säljs.
- på spanska:
"bestrålet/..." eller "strålekonserveret" eller "behandlet med ioniserende stråling" eller "konserveret med ioniserende stråling"
- på engelska:
"traité par rayonnements ionisants" eller "traité par ionisation."
- på nederländska:
"irradiado" eller "tratado por irradiação" eller "tratado por radiação ionizante".
- på svenska:
1. Ingredienser skall anges i enlighet med denna artikel och bilagorna I, II och III.
- kolsyrat vatten, om det framgår av försäljningsnammet att vattnet har kolsyrats,
- smör,
c) varor som består av en enda ingrediens
3. I fråga om drycker som innehåller mer än 1,2 volymprocent alkohol skall rådet på förslag av kommissionen före den 22 december 1982, bestämma reglerna för hur ingredienser skall anges.
c) Som ingredienser anses inte
- vilkas förekomst i ett visst livsmedel uteslutande beror på att de ingått i en eller flera ingredienser i det aktuella livsmedlet, förutsatt att tillsatserna inte har någon teknisk funktion i den färdiga varan,
d) Enligt der förfarande som fastställs i artikel 20.2 kan det i vissa fall avgöras huruvida villkoren i c ii och iii är uppfyllda.
- Tillsatt vatten och flyktiga ämnen skall anges i storleksordning efter vikt i den färdiga varan; den mängd vatten som tillsatts som ingrediens i ett livsmedel skall beräknas genom att den färdiga varans totala mängd minskas med den totala mängden av övriga använda ingredienser. Denna mängd behöver inte beaktas om den inte överstiger 5 % av den färdiga varans vikt.
- Ingredienserna i frukt eller grönsaksblandningar, i vilka ingen särskild frukt eller grönsak påtagligt dominerar med hänsyn till vikt får anges i annan ordning, förutsatt att denna ingrediensförteckning åtföljs av uttrycket "i varierande proportion" eller liknande uttryck.
Undantag:
Beteckningen "stärkelse" i bilaga I måste dock alltid kompletteras med en angivelse av vilken specifik växt den framställts ur, då denna ingrediens kan innehålla gluten.
Beteckningen "modifierad stärkelse" i bilaga II måste dock alltid kompletteras med en angivelse av vilken specifik växt den framställs ur, då denna ingrediens kan innehålla gluten.
7. Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser, får fastställa att det namn, som ett visst livsmedel säljs under, skall åtföljas av uppgift om en eller flera särskilda ingredienser.
8. I det fall som avses i punkt 4 b får en sammansatt ingrediens uttryckt i total vikt ingå i ingrediensförteckningen under sin egen beteckning, om denna fastställts enligt lag eller sedvana, förutsatt att den omedelbart följs av en uppräkning av de ingredienser som ingår i den sammansatta ingrediensen.
b) Om den sammansatta ingrediensen är ett livsmedel för vilket någon ingrediensförteckning inte krävs enligt gemenskapsregler.
b) om detta utgör en lag som normalt inte konsumeras.
2. Den angivelse som avses i punkt 1 skall vara obligatorisk,
c) om den berörda ingrediensen eller kategorin av ingredienser är nödvändig för att känneteckna livsmedlet och särskilja det från produkter som det skulle kunna förväxlas med på grund av sitt namn och utseende, eller
a) på en ingrediens eller kategori av ingredienser
- som används i små mängder i aromgivande syfte, eller
c) i de fall som avses i artikel 6.5 fjärde och femte strecksatserna,
5. Den angivelse som avses i punkt 1 skall antingen ingå i det namn under vilket livsmedlet säljs eller anges omedelbart därintill eller också anges i ingrediensförteckningen i anslutning till ingrediensen eller kategorin av ingredienser i fråga.
1. Nettoinnehållet i färdigförpackade livsmedel skall anges
varvid liter, centiliter, milliliter, kilogram eller gram skall användas allt efter omständigheterna.
2. a) Om gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser innehåller föreskrifter om att ett innehåll skall anges på ett visst sätt (t.ex. nominell kvantitet, minimikvantitet, genomsnittskvantitet) skall denna kvantitet anses som nettoinnehåll enligt detta direktiv.
Det förfarande som fastställs i artikel 19 skall tillämpas på varje sådan nationell bestämmelse.
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24 skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt denna punkt.
4. Om ett livsmedel i fast form ligger i en lag, skall även livsmedlets avrunna vikt anges i märkningen.
Metoder för att kontrollera avrunnen vikt skall bestämmas i enlighet med det förfarande som fastställs i artikel 20.2.
b) vars nettoinnehåll är mindre än 5 g eller 5 ml; dock skall denna bestämmelse inte gälla för kryddor och örter.
6. De gemenskapsbestämmelser som avses i punkterna 1 andra stycket, 2 b, 2 d och 5 andra stycket skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
Det skall anges i enlighet med bestämelserna i punkterna 2-5.
- "Bäst före utgången av... " i övriga fall.
- en hänvisning till var på märkningen datumet finns angivet.
Dock är det i fråga om livsmedel
- med längre hållbarhetstid än 18 månader tillräckligt att ange året.
- Färsk frukt och färska grönsaker, inklusive potatis, som inte skalats, delats i bitar eller behandlats på liknande sätt. Detta undantag skall inte tillämpas på groddar och liknande produkter såsom skott av baljväxter.
- Läskedrycker, fruktjuice, fruktnektar och alkoholhaltiga drycker i separata kärl på mer än fem liter och avsedda för storkök.
- Koksalt.
Artikel 10
Orden skall följas av
Dessa uppgifter skall följas av en beskrivning av de förvaringsanvisningar som man måste rätta sig efter.
Artikel 11
Det förfarande som fastställs i artikel 19 skall tillämpas på sådana nationella bestämmelser.
De bestämmelser som gäller angivande av alkoholhalten uttryckt i volym skall i fråga om varor som faller under tariffrubrikerna nr 22.04 och 22.05 fastställas i särskilda gemenskapsbestämmelser som gäller för dessa varor.
1. a) I fråga om färdigpackade livsmedel skall de uppgifter som anges i artikel 3 och artikel 4.2 finnas på förpackningen eller på en etikett som är fästad vid denna.
c) I de fall som avses i b skall de uppgifter som avses i artikel 3.1.1, 3.1.5 och 3.1.7 och, i tilllämpliga fall, de som avses i artikel 10 också finas på den yttre förpackning, i vilken livsmedlen presenteras när de saluförs.
3. De uppgifter som räknas upp i artikel 3.1.1, 3.1.4, 3.1.5 och 3.1.10 skall förekomma i samma synfält.
I detta fall skall punkt 3 inte gälla.
Artikel 14
Artikel 15
1. Medlemsstaterna skall säkerställa att det inom deras territorier är förbjudet att saluföra livsmedel för vilka uppgifterna enligt artikel 3 och artikel 4.2 inte ges på ett språk som med lätthet förstås av konsumenten, såvida inte konsumenten faktiskt informeras genom andra åtgärder som fastställs i enlighet med det förfarande som anges i artikel 20.2 beträffande en eller flera uppgifter i märkningen.
Artikel 17
1. Medlemsstater får inte förbjuda handel med livsmedel som följer reglerna i detta direktiv genom att tillämpa nationella icke harmoniserade bestämmelser för märkning och presentation av vissa livsmedel eller av livsmedel i allmänhet.
- förebygga oredlighet, såvida inte sådana bestämmelser kan befaras hindra tillämpningen av de definitioner och regler som fastställs genom detta direktiv,
När det hänvisas till denna artikel skall följande förfarande användas, om en medlemsstat skull bedöma det som nödvändigt att anta ny lagstiftning:
Om så skulle vara fallet, skall kommissionen före utgången av denna period inleda det förfarande som fastställs i artikel 20.2 för att avgöra huruvida de planerade åtgärdena kan genomföras, om det är nödvändigt med lämpliga ändringar.
2. När det hänvisas till denna punkt, skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i beslutet.
Artikel 21
Detta direktiv skall inte inverka på sådana gemenskapsbestämmelser om märkning och presentation av vissa livsmedel som redan antagits den 22 december 1978.
Detta direktiv skall inte gälla varor avsedda för export utanför gemenskapen.
Artikel 25
1. Direktiv 79/112/EEG i dess lydelse enligt direktiven i bilaga IV del A skall upphöra att gälla utan att det påverkar medlemsstaternas förpliktelsre vad gäller de tidsfrister för genomförande som anges i bilaga IV del B.
Kommissionens direktiv 2000/63/EG
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(2) I kommissionens direktiv 96/77/EG av den 2 december 1996 om särskilda renhetskriterier för andra livsmedelstillsatser än färgämnen och sötningsmedel(5), ändrat genom direktiv 98/86/EG(6), fastställs renhetskriterier för ett antal livsmedelstillsatser. Detta direktiv bör nu kompletteras med renhetskriterier för de återstående livsmedelstillsatserna i direktiv 95/2/EG.
(5) Om livsmedelstillsatser bereds genom produktionsmetoder eller från utgångsmaterial som avsevärt skiljer sig från dem som utvärderats av Vetenskapliga livsmedelskommittén, eller från dem som anges i detta direktiv, bör Vetenskapliga livsmedelskommittén göra en säkerhetsutvärdering av dessa tillsatser, med särskild tonvikt på renhetskriterierna.
Artikel 1
2) Bilaga II till detta direktiv skall läggas till i bilagan.
2) När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Europaparlamentets och rådets direktiv 2000/69/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) I enlighet med artikel 4.5 i rådets direktiv 96/62/EG av den 27 september 1996 om utvärdering och säkerställande av luftkvaliteten(6) skall rådet anta de bestämmelser som avses i punkt 1 samt i punkterna 3 och 4 i den artikeln.
(6) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(7).
(9) Bensen är ett för människor genotoxiskt carcinogen, och det är inte möjligt att fastställa något tröskelvärde under vilket det inte föreligger någon hälsorisk.
(12) Standardiserade och tillförlitliga mätmetoder och gemensamma kriterier för placeringen av mätstationer är av stor betydelse för bedömningen av luftkvaliteten om man vill uppnå jämförbara uppgifter över hela gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Syftet med detta direktiv är att
c) inhämta tillförlitliga uppgifter om koncentrationer av bensen och koloxid i luften, och säkerställa att dessa uppgifter görs tillgängliga för allmänheten,
Definitioner
a) övre utvärderingströskel: den nivå som avses i bilaga III under vilken en kombination av mätningar och modelleringsmetoder kan användas för att utvärdera luftkvaliteten, i enlighet med artikel 6.3 i direktiv 96/62/EG,
Artikel 3
Den toleransmarginal som anges i bilaga I skall tillämpas i enlighet med artikel 8 i direktiv 96/62/EG.
- tillhandahåller erforderlig motivering för en sådan förlängning,
Det gränsvärde för bensen som tillåts under den tidsbegränsade förlängningen får emellertid inte överskrida 10 μg/m3.
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att koncentrationen av koloxid i luften, som utvärderats i enlighet med artikel 5, inte överskrider gränsvärdet som anges i bilaga II med hänsyn till de datum som där anges.
Utvärdering av koncentrationer
2. Kriterierna för att bestämma var provtagningsplatserna för mätning av bensen- och koloxid i luften skall placeras är de som anges i bilaga IV. Minsta antalet provtagningsplatser för fasta mätningar av koncentrationer av de berörda föroreningarna fastställs i bilaga V, och de skall installeras i alla zoner eller tätbebyggelser där mätningar krävs om fasta mätningar är den enda källan för uppgifter om koncentrationer i dessa.
5. Referensmetoderna för analys och provtagning av bensen och koloxid anges i avsnitten I och II i bilaga VII. I avsnitt III i bilaga VII kommer referensmetoder för luftkvalitetsmodellering att anges när sådana tekniker finns tillgängliga.
Artikel 6
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 7
Informationen om koncentrationerna av bensen i luften skall, i form av ett genomsnittsvärde för de tolv senaste månaderna, uppdateras minst var tredje månad och, där det är praktiskt genomförbart, en gång i månaden. Information om koncentrationerna av koloxid i luften skall, i form av ett högsta genomsnittsvärde för åtta timmar i följd, uppdateras minst en gång per dag och där det är praktiskt genomförbart en gång per timme.
3. Information till allmänheten och organisationer i enlighet med punkterna 1 och 2 skall vara tydlig, begriplig och lättillgänglig.
1. Senast den 31 december 2004 skall kommissionen till Europaparlamentet och rådet överlämna en rapport som är grundad på de erfarenheter som gjorts vid tillämpningen av detta direktiv, och särskilt på resultaten av den senaste vetenskapliga forskningen om effekterna på människors hälsa, varvid särskild hänsyn skall tas till känsliga befolkningsgrupper, och på ekosystemen av exponering för bensen och koloxid, samt på den tekniska utvecklingen, inbegripet framsteg i fråga om mätmetoder och andra sätt att utvärdera bensen- och koloxidkoncentrationer i luften.
b) Möjligheterna till ytterligare minskningar av förorenande utsläpp från alla relevanta källor, med beaktande av teknisk genomförbarhet och kostnadseffektivitet.
e) De erfarenheter som gjorts i medlemsstaterna vid tillämpningen av detta direktiv, i synnerhet de förhållanden, enligt föreskrifterna i bilaga IV, under vilka mätningarna utförts.
Påföljder
Genomförande
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Kommissionens förordning (EG) nr 645/2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets direktiv 90/642/EEG av den 27 november 1990 om fastställande av gränsvärden för bekämpningsmedelsrester i och på produkter av vegetabiliskt ursprung inklusive frukt och grönsaker(3), senast ändrat genom direktiv 1999/71/EG, särskilt artikel 4 i detta, och
(2) Erfarenheterna från utformning och tillämpning av kommissionens rekommendationer har visat att flerårig planering, med möjlighet till årliga justeringar, torde vara det effektivaste sättet att upprätta Europeiska gemenskapens samordnade kontrollprogram.
(5) Kommissionen bör bidra ekonomiskt till åtgärder som stärker andra aspekter av samarbetet beträffande kontroll av bekämpningsmedelsrester på gemenskapsnivå. Särskilt bör sådan verksamhet stödjas som på sikt främjar utvecklingen av ett system på gemenskapsnivå som gör det möjligt att på grundval av data från kontrollprogrammen beräkna det dagliga intaget av bekämpningsmedelsrester via kosten.
(8) Både i direktiv 90/642/EEG i dess ändrade form och i direktiv 86/362/EEG i dess ändrade form ges förutsättningar för att det skall kunna vidtas åtgärder på gemenskapsnivå vid rapporterade överträdelser och att de tillämpningsföreskrifter skall antas som krävs för att kontrollen skall fungera väl.
(11) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för växtskydd.
1. Kommissionens rekommendationer enligt bestämmelserna i artikel 7.2 b i direktiv 86/362/EEG och artikel 4.2 b i direktiv 90/642/EEG får omfatta perioder på mellan ett och fem år.
Kommissionen skall underlätta tillämpningen av bestämmelserna i artikel 7.2 och 7.3 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG på följande sätt:
a) regelbundet anordnade kvalifikationsprövningar, i princip vartannat år, av alla laboratorier som utför analyser, i syfte att säkerställa kvalitet, noggrannhet och jämförbarhet av de uppgifter som medlemsstaterna lämnar till kommissionen och övriga medlemsstater årligen och som insamlas och sammanställs av kommissionen för offentliggörande i enlighet med artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG,
d) till organisation av andra åtgärder på gemenskapsnivå, definierade av kommissionen och Ständiga kommittén för växtskydd, som krävs för en korrekt tillämpning av artikel 7.2 och 7.3 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG.
2. I det kommissionsbeslut som avses i punkt 1 skall särskilt anges
- en sammanfattande beskrivning av åtgärden,
Medlemsstaterna skall säkerställa att de analysresultat som årligen översänds till kommissionen och till övriga medlemsstater i enlighet med bestämmelserna i artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG har erhållits från laboratorier som
Medlemsstaterna skall dessutom säkerställa att endast laboratorier som har deltagit i en tidigare eller skall delta i nästa omgång av gemenskapens relevanta kvalifikationsprövningar enligt artikel 2.2 a i denna förordning deltar i gemenskapens samordnade program.
2. Tjänstemännen skall besöka de nationella myndigheterna i varje medlemsstat, som skall samarbeta med kommissionens utsedda tjänstemän och ge dem all nödvändig assistans i deras arbete. Besöksprogrammen skall organiseras och genomföras i samarbete med den berörda medlemsstaten. De nationella myndigheterna skall under alla omständigheter fortsätta att ansvara för att kontrollåtgärderna genomförs.
5. Kommissionen skall regelbundet genom skriftliga rapporter inom Ständiga kommittén för växtskydd underrätta alla medlemsstater om resultatet av kontrollbesöken i varje medlemsstat. Kommissionen skall underrätta Europaparlamentet. Kommissionen skall också regelbundet offentliggöra rapporterna.
Denna förordning träder i kraft den 1 april 2000.
av den 27 mars 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
(2) Mot bakgrund av uppdragen för den rådgivande kommittén för fiske och vattenbruk (nedan kallad den rådgivande kommittén), vilken förnyades genom kommissionens beslut 1999/478/EG(1), kan målen dialog och öppenhet främjas genom nya åtgärder, som syftar dels till att bättre organisera den rådgivande kommitténs möten, dels till att sprida information till de berörda grupperna om insatser och resultat.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- de europeiska branschorganisationernas möten för att förbereda mötena i den rådgivande kommittén,
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om komplettering av bilagan till kommissionens förordning (EG) nr 1107/96 om registrering av geografiska beteckningar och ursprungsbeteckningar enligt förfarandet i artikel 17 i förordning (EEG) nr 2081/92
med beaktande av kommissionens förslag,
(1) För vissa beteckningar som medlemsstaterna har meddelat i enlighet med artikel 17 i förordning (EEG) nr 2081/92 har det begärts kompletterande uppgifter för att säkerställa att dessa beteckningar uppfyller kraven i artiklarna 2 och 4 i nämnda förordning. Efter granskning av dessa kompletterande uppgifter har det visat sig att dessa beteckningar stämmer överens med nämnda artiklar. De bör därför registreras och läggas till i bilagan till kommissionens förordning (EG) nr 1107/96(2).
Artikel 1
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
om närmare bestämmelser för genomförandet av rådets förordning (EG) nr 1260/1999 avseende stödberättigande utgifter i samband med insatser som medfinansieras av strukturfonderna
med beaktande av rådets förordning (EG) nr 1260/1999 av den 21 juni 1999 om allmänna bestämmelser för strukturfonderna(1), särskilt artikel 30.3 och artikel 53.2 i denna,
(1) I artikel 1.3 i rådets förordning (EG) nr 1257/1999 av den 17 maj 1999 om stöd från Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) till utveckling av landsbygden och om ändring och upphävande av vissa förordningar(2) anges att åtgärder för utveckling av landsbygden som är integrerade med åtgärder som främjar utvecklingen och den strukturella anpassningen i regioner vars utveckling släpar efter (mål 1) eller som åtföljer åtgärder till stöd för ekonomisk och social omställning i områden med strukturella svårigheter (mål 2) i de berörda områdena, skall beakta strukturfondernas särskilda syften med gemenskapens stöd i enlighet med villkoren i förordning (EG) nr 1260/1999. I artikel 2 i förordning (EG) nr 1257/1999 anges vilka typer av åtgärder som kan komma i fråga för stöd till utveckling av landsbygden.
(4) I artikel 2 i rådets förordning (EG) nr 1263/1999 av den 21 juni 1999 om Fonden för fiskets utveckling(5) anges vilken typ av åtgärder som kan genomföras med finansiellt stöd från FFU. I rådets förordning (EG) nr 2792/1999(6) fastställs närmare föreskrifter och villkor för strukturåtgärderna inom fiskerisektorn.
(7) Artiklarna 87 och 88 i fördraget är tillämpliga på verksamhet som medfinansieras av strukturfonderna. Ett kommissionsbeslut om att godkänna en stödform innebär inte någon förhandsbedömning av statsstödsreglerna och befriar inte medlemsstaten från sina skyldigheter enligt dessa artiklar.
Artikel 1
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EG) nr 2037/2000 om ämnen som bryter ned ozonskiktet vad gäller dosaerosoler och läkemedelspumpar
med beaktande av Ekonomiska och sociala kommitténs yttrande(1),
av följande skäl:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"f) dosaerosoler som innehåller klorfluorkarboner och doseringsmekanismer som innehåller klorfluorkarboner för hermetiskt tillslutna apparater avsedda att implanteras i människokroppen för att avge uppmätta läkemedelsdoser, vilka enligt artikel 4.1 kan erhålla ett tillfälligt undantag enligt det förfarande som avses i artikel 18.2."
Rådets förordning (EG) nr 2578/2000
med beaktande av rådets förordning (EEG) nr 3759/92 av den 17 december 1992 om den gemensamma organisationen av marknaden för fiskeri- och vattenbruksprodukter(1), särskilt artikel 2.3 i denna,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 3 skall
- Havsruda (Spondyliosoma cantharus) och"
- Stor kammussla (Pecten maximus)
3. Artikel 7.1 skall ersättas med följande text:
Artikel 2
av den 16 november 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 26, 95 och 133 i detta,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) Varje översyn av kodexen bör, utan att det införs några hinder för den internationella handeln, utgöra ett tillfälle att inrätta instrument och förfaranden som gör det möjligt att förebygga bedrägeri, med tanke på att förebyggande av bedrägeri är ett av de bästa sätten att skydda skattebetalarnas pengar enligt rådets slutsatser av den 19 maj 1998.
(5) Det bör föreskrivas att en tulldeklaration som har upprättats med databehandlingsteknik inte behöver åtföljas av vissa dokument.
(8) Det kan vara lämpligt att i vissa frizoner tillåta att tullformaliteter fullgörs och myndigheternas tullkontroller utförs i enlighet med tullagerförfarandet.
(11) Det är, när det gäller förmånsbehandling, nödvändigt att definiera vad som avses med begreppen misstag som begåtts av tullmyndigheter och god tro hos gäldenären. Gäldenären bör inte bära ansvaret för att systemet fungerar dåligt på grund av ett misstag som har begåtts av myndigheter i tredje land. Sådana myndigheters utfärdande av ett oriktigt ursprungsintyg bör emellertid inte anses som ett misstag om ursprungsintyget har utfärdats på grundval av en ansökan som innehåller oriktiga uppgifter. Oriktigheten i de uppgifter som exportören lämnat i sin ansökan bör bedömas på grundval av alla de faktiska förhållanden som ansökningen innehåller. En gäldenär kan åberopa god tro när han kan visa att han handlat med tillbörlig aktsamhet, utom då ett yttrande om att det finns välgrundade tvivel har offentliggjorts i Europeiska gemenskapernas officiella tidning.
(14) De åtgärder som krävs för att genomföra förordning (EEG) nr 2913/92 bör fastställas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(6).
Artikel 1
"24. kommittéförfarande: det förfarande som avses dels i artiklarna 247 och 247a, dels i artiklarna 248 och 248a."
"2. För tulldeklarationer som upprättas med hjälp av databehandlingsteknik får tullmyndigheterna tillåta att de åtföljande dokument som avses i artikel 62.2 inte bifogas deklarationen. I detta fall skall dokumenten hållas tillgängliga för tullmyndigheterna."
5. I artikel 117 c skall följande mening läggas till:"De fall där de ekonomiska villkoren skall anses vara uppfyllda får fastställas enligt kommittéförfarandet."
1. Restitutionssystemet får användas för alla varor. Det får dock inte användas i de fall där, vid tidpunkten för mottagandet av deklarationen om övergång till fri omsättning
- importvarorna omfattas av krav på att import- eller exportintyg skall uppvisas enligt den gemensamma jordbrukspolitiken, eller
3. Undantag från bestämmelserna i punkterna 1 och 2 får fastställas enligt kommittéförfarandet."
De fall i vilka förfarandet för bearbetning under tullkontroll får användas och de särskilda villkoren för användningen skall fastställas enligt kommittéförfarandet."
"Artikel 142
10. I artikel 153 skall följande stycke läggas till:"Utan hinder av artikel 151 får det enligt kommittéförfarandet fastställas i vilka fall och på vilka särskilda villkor som det vid övergång till fri omsättning av varor efter passiv förädling kan medges att kostnaden för förädlingsprocessen används som grund för taxeringen vid tillämpningen av Europeiska gemenskapernas tulltaxa."
12. I artikel 168 skall punkt 1 ersättas med följande:
"Artikel 168a
2. De frizoner som avses i artiklarna 37, 38 och 205 omfattar inte frizoner enligt punkt 1."
När det i tullagstiftningen föreskrivs en gynnsam behandling i tullhänseende för varor med anledning av deras beskaffenhet eller deras användning för särskilda ändamål, eller fullständig eller partiell befrielse från import- eller exporttullar med stöd av artiklarna 21, 82, 145 eller 184-187, skall den gynnsamma behandlingen eller befrielsen även tillämpas då en tullskuld har uppkommit i enlighet med artiklarna 202-205, 210 eller 211, om den berörda partens uppträdande inte låter förmoda bedrägligt förfarande eller påtaglig försummelse och om denne kan styrka att de övriga villkoren för tillämpning av den gynnsamma behandlingen eller befrielsen är uppfyllda."
16. I artikel 220.2 skall punkt b ersättas med följande:
Utfärdande av ett felaktigt ursprungsintyg skall emellertid inte anses utgöra ett misstag när det grundar sig på felaktiga uppgifter från exportören, utom t.ex. i sådana fall då det är uppenbart att de utfärdande myndigheterna var eller borde ha varit medvetna om att varorna inte uppfyllde villkoren för förmånsbehandling.
17. I artikel 221 skall punkt 3 ersättas med följande punkter:
18. I artikel 222 skall punkt 2 ersättas med följande:
- när varor tas i beslag för att därefter förverkas i enlighet med artikel 233c andra strecksatsen eller artikel 233d, eller
"Artikel 247
1. Kommissionen skall biträdas av en tullkodexkommitté (nedan kallad kommittén).
3. Kommittén skall själv anta sin arbetsordning.
Artikel 248a
Den tid som avses i artikel 4.3 i beslut 1999/468/EG skall vara tre månader.
Kommittén får behandla alla de frågor om tullagstiftningen som tas upp av ordföranden, antingen på dennes initiativ eller på begäran av företrädaren för en medlemsstat."
Kommissionens förordning (EG) nr 2785/2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) I artikel 4.1a a i kommissionens förordning (EG) nr 296/96 av den 16 februari 1996 om de uppgifter som medlemsstaterna skall sända in för månatlig bokföring av de utgifter som finansieras genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) samt fastställande av vissa tillämpningsföreskrifter för rådets förordning (EG) nr 1259/1999(5), senast ändrad genom förordning (EG) nr 2761/1999(6), föreskrivs att förskotten för utgifter, bokförda under EUGFJ:s garantisektion, skall upprättas och utbetalas i euro till deltagande medlemsstater. Förskotten som skall utbetalas i början av januari 2001 avser utgifter som verkställts under perioden 16.10.2000-30.11.2000. I Greklands fall bör dessa förskott för sista gången utbetalas i nationell valuta.
Artikel 1
2. I artikel 4.1a c skall följande läggas till:"För utgifter som Grekland verkställt under perioden 16.10.2000-30.11.2000 skall förskotten utbetalas i nationell valutaenhet eller i nationell valuta."
Kommissionens förordning (EG) nr 2858/2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för bearbetade produkter av frukt och grönsaker.
Förordning (EG) nr 2125/95 ändras på följande sätt:
av den 19 december 2000
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Vissa översättningsskillnader mellan den tyska texten och de övriga språkversionerna bör utjämnas när det gäller gränsöverskridande handel med obearbetad gödsel. Med tanke på möjliga sjukdomsrisker är det också lämpligt att införa bättre kontroll av sådana förflyttningar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"1. a) Handel med obearbetad gödsel av andra arter än fjäderfä och hästdjur skall vara förbjuden, med undantag för gödsel som:
är avsedd att spridas under kontroll av behöriga myndigheter på mark som utgör en del av eller tillhör samma anläggning som, vare sig åtskild eller ej, ligger på båda sidor om gränsen mellan medlemstater och inom ett avstånd på cirka 20 km. För att en anläggning skall kunna godkännas måste dess ägare föra register över sådana förflyttningar över gränser. Den behöriga myndigheten skall föra register över sådana godkända anläggningar."
Artikel 3
av den 24 januari 2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av rådets direktiv 88/407/EEG av den 14 juni 1988 om djurhälsokrav som är tillämpliga vid handel inom gemenskapen med och import av djupfryst sperma från tamdjur av nötkreatur(3), senast ändrat genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 5.2 i detta,
med beaktande av rådets direktiv 90/429/EEG av de 26 juni 1990 om djurhälsokrav som är tillämpliga vid handel inom gemenskapen med och import av sperma från tamdjur av svin(6), senast ändrat genom beslut 1999/608/EG(7), särskilt artikel 5.3 i detta,
(1) Det är tillåtet att bedriva handel inom gemenskapen med nötkreatur, svin, får, getter och hästdjur från sådana uppsamlingscentraler som godkänts av de behöriga myndigheterna i de medlemsstater där de är belägna.
(4) Varje enskild medlemsstat bör till kommissionen och övriga medlemsstater sända förteckningar över de uppsamlingscentraler, seminstationer och embryosamlingsgrupper i det egna landet som medlemsstaten har godkänt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Förteckningarna skall vara utformande enligt mallarna i bilaga II.
Detta beslut riktar sig till medlemsstaterna.
om ändring av avfallsförteckningen i beslut 2000/532/EG
(2001/118/EG)
med beaktande av rådets direktiv 75/442/EEG av den 15 juli 1975 om avfall(1), senast ändrat genom kommissionens beslut 96/350/EG(2), särskilt artikel 1 a i detta,
(1) Kommissionens beslut 2000/532/EG(5) av den 3 maj 2000 om ersättning av beslut 94/3/EG om en förteckning över avfall i enlighet med artikel 1 a i rådets direktiv 75/442/EEG om avfall, och rådets beslut 94/904/EG om upprättande av en förteckning över farligt avfall i enlighet med artikel 1.4 i rådets direktiv 91/689/EEG om farligt avfall bör ändras mot bakgrund av de anmälningar som inkommit från medlemsstaterna i enlighet med artikel 1.4 andra strecksatsen i direktiv 91/689/EEG.
Artikel 1
"Artikel 2
- ett eller flera ämnen som klassificeras(7) som mycket giftiga vid en total koncentration >= 0,1 %,
- ett eller flera frätande ämnen som klassificeras som R35 vid en total koncentration >= 1 %,
- ett eller flera irriterande ämnen som klassificeras som R36, R37 eller R38 vid en total koncentration >= 20 %,
- ett ämne som är skadligt för fortplantningen (kategori 1 eller 2) och som klassificeras som R60 eller R61 vid en koncentration >= 0,5 %,
- ett mutagent ämne (kategori 3) som klassificeras som R40 vid en koncentration >= 1 %."
Det här beslutet skall tillämpas från och med den 1 januari 2002.
Kommissionens beslut
[delgivet med nr K(2001) 426]
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) Ändringarna gäller undersökning och identifiering av virus som orsakar viral hemorragisk septikemi (VHS) och smittsam hematopoetisk nekros (IHN) samt anpassning till ändringarna av direktiv 91/67/EEG.
(6) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Provtagningsplaner och diagnostiska metoder för påvisande och bekräftelse av viral hemorragisk septikemi (VHS) och infektiös hematopoetisk nekros (IHN) fastställs i bilagan.
Artikel 3
av den 23 juli 2001
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT
med beaktande av kommissionens förslag, och
(2) Förteckningen kan kompletteras eller ändras med hänsyn till hur hälsosituationen utvecklas i gemenskapen.
(5) Bluetongue är en insektsburen virussjukdom hos får, getter, nötkreatur och andra idisslare.
(8) Vissa områden inom gemenskapen måste, på grund av klimatförhållanden, betraktas som högriskområden för bluetongue.
(11) För att det finansiella stödet från gemenskapen skall kunna ges, måste de relevanta bestämmelser följas som anges i beslut 90/424/EEG och, när det gäller infektiös laxanemi, i rådets direktiv 93/53/EEG av den 24 juni 1993 om gemenskapens minimiåtgärder för bekämpning av vissa fisksjukdomar(2).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Bluetongue i högriskområden eller områden där sjukdomen är endemisk(6)".
Rådets beslut
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(3) För tydlighetens skull bör det uttryckligen anges att uteslutande fett- och oljeblandningar från oljeavskiljare som endast innehåller ätliga oljor och fetter får betraktas som icke-farliga.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
om uppdatering av beslut 2000/112/EG om fördelning av beredskapslager av antigener mellan antigenbanker
(2001/660/EG)
med beaktande av rådets beslut 90/424/EEG av den 26 juni 1990 om utgifter inom veterinärområdet(1), senast ändrat genom beslut 2001/12/EG(2), särskilt artikel 14 i detta,
(1) I enlighet med beslut 91/666/EEG ingår inköp av antigener som ett led i gemenskapens åtgärder för att upprätta beredskapslager av vacciner mot mul- och klövsjuka.
(4) Genom kommissionens beslut 97/348/EG(7), senast ändrat genom beslut 2000/112/EG, fastställs bestämmelser för inköp av mul- och klövsjukevirusantigen A22-Iraq, C1 och ASIA1.
(7) Efter skriftliga uppgifter från leverantören om tilldelning och fördelning till de godkända anläggningarna av antigen som inköpts enligt beslut 2000/569/EG är det också lämpligt att uppdatera bilagan till beslut 2000/112/EG med närmare uppgifter om antigenreservernas fördelning mellan de antigenbanker som upprättats inom ramen för gemenskapens åtgärder för att skapa beredskapslager av vacciner mot mul- och klövsjuka och att ändra kommissionens beslut 93/590/EG och 97/348/EG.
Artikel 1
Detta beslut riktar sig till medlemsstaterna.
om bekämpning av bedrägeri och förfalskning som rör andra betalningsmedel än kontanter
med beaktande av Fördraget om Europeiska unionen, särskilt artikel 34.2 b i detta,
av följande skäl:
(3) Rådet anser att vissa former av bedrägeri som rör andra betalningsmedel än kontanter är så allvarliga och utvecklas på ett sådant sätt att det krävs övergripande lösningar. Rekommendation nr 18 i handlingsplanen för bekämpande av den organiserade brottsligheten(3), godkänd av Europeiska rådet i Amsterdam den 16-17 juni 1997, samt punkt 46 i rådets och kommissionens handlingsplan för att på bästa sätt genomföra bestämmelserna i Amsterdamfördraget om upprättande av ett område med frihet, säkerhet och rättvisa(4), godkänd av Europeiska rådet i Wien den 11-12 december 1998, innebär att åtgärder måste vidtas på detta område.
(6) Kommissionen överlämnade till rådet den 1 juli 1998 meddelandet "En ram för åtgärder för att bekämpa bedrägeri och förfalskning som rör andra betalningsmedel än kontanter", i vilket det förespråkas en EU-politik som omfattar både förebyggande och repressiva aspekter av problemet.
(9) Det är nödvändigt att dessa typer av beteenden anses vara straffbara gärningar i samtliga medlemsstater och att effektiva, proportionella och avskräckande påföljder införs för fysiska och juridiska personer som har begått eller är ansvariga för sådana brott.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
I detta rambeslut avses med
Artikel 2
a) Stöld eller annat olovligt tillgrepp av ett betalningsinstrument.
d) Bedräglig användning av ett betalningsinstrument som stulits eller olovligen tillgripits eller som är helt eller delvis förfalskat.
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att följande handlingar är straffbara när de är uppsåtliga:
Artikel 4
Bedräglig tillverkning, mottagande, anskaffande, försäljning eller överlämnande till annan person eller innehav av
Artikel 5
Artikel 6
Artikel 7
- befogenhet att företräda den juridiska personen, eller
samt för medhjälp eller anstiftan till ett sådant brott.
Artikel 8
a) fråntagande av rätt till offentliga förmåner eller stöd,
d) rättsligt beslut om avveckling av verksamheten.
Behörighet
b) av en av dess medborgare, dock med förbehåll för att den medlemsstatens lagstiftning kan kräva att gärningen är straffbar även i det land där den begicks, eller
- punkt 1 b,
Artikel 10
b) Varje medlemsstat skall, när en av dess medborgare anklagas för att i en annan medlemsstat ha begått ett brott som innefattar de handlingar som beskrivs i artiklarna 2, 3, 4 och 5 och om den inte utlämnar denna person till den andra medlemsstaten enbart på grund av dennes nationalitet, lägga fram fallet för sina behöriga myndigheter i syfte att om så är lämpligt väcka åtal. För att möjliggöra att åtal väcks skall akter, information och bevisföremål som rör brottet överlämnas enligt förfarandena i artikel 6.2 i Europeiska utlämningskonventionen av den 13 december 1957. Den ansökande medlemsstaten skall informeras om det åtal som väcks och om dess resultat.
Samarbete mellan medlemsstaterna
Artikel 12
2. Varje medlemsstat skall meddela rådets generalsekretariat eller kommissionen vilket eller vilka organ som utgör kontaktpunkt enligt punkt 1. Generalsekretariatet skall meddela övriga medlemsstater vilka dessa kontaktpunkter är.
Detta rambeslut skall tillämpas i Gibraltar.
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta rambeslut senast den 2 juni 2003.
Ikraftträdande
av den 21 januari 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 47.2 i detta,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) Med hänsyn till utvecklingen på marknaden bör fondföretagens investeringsmöjligheter utökas till att omfatta andra, tillräckligt likvida, finansiella instrument än överlåtbara värdepapper. Finansiella instrument som kan ingå som tillgångar i ett fondföretags värdepappersportfölj anges i detta direktiv. Att investera så att en portfölj återspeglar ett visst index är en förvaltningsteknik.
(5) Det är lämpligt att säkerställa att begreppet "reglerad marknad" i detta direktiv stämmer överens med det i direktiv 93/22/EEG av den 10 maj 1993 om investeringstjänster inom värdepappersområdet(5).
(8) För att beakta marknadsutvecklingen och mot bakgrund av genomförandet av den ekonomiska och monetära unionen, bör fondföretag tillåtas att investera i inlåning. För att säkerställa en tillräcklig likviditet för sådana investeringar skall dessa tillgodohavanden kunna betalas ut på begäran eller kunna dras tillbaka. Om tillgodohavandena finns i ett kreditinstitut med säte i en icke-medlemsstat, bör detta institut omfattas av tillsynsregler likvärdiga med dem som gäller inom gemenskapslagstiftningen.
(11) Fondföretag bör uttryckligen tillåtas att investera i finansiella derivatinstrument, såväl inom ramen för sin allmänna investeringspolicy som i syfte att säkra tillgångar, för att uppnå ett finansiellt mål eller den riskprofil som angetts i prospektet. För att säkerställa att investerarna skyddas är det nödvändigt att begränsa den maximala riskexponeringen i förhållande till finansiella derivatinstrument så att den inte överskrider det totala nettovärdet av fondföretagets portfölj. För att säkerställa ständig medvetenhet om riskerna och åtagandena vid derivattransaktioner och kontrollera att investeringsgränserna hålls, måste dessa risker och åtaganden fortlöpande mätas och övervakas. Slutligen, för att skapa ett skydd för investerarna genom tillhandahållande av information, bör fondföretagen beskriva sina strategier, metoder och sina investeringsgränser för derivattransaktioner.
(14) Vissa portföljförvaltningsmetoder för företag för kollektiva investeringar som främst investerar i aktier och/eller skuldebrev bygger på efterbildningen av aktieindex och/eller index för skuldebrev. Fondföretag bör tillåtas att efterbilda välkända och erkända aktieindex och/eller index för skuldförbindelser. Det kan därför vara nödvändigt att införa flexiblare riskspridningsregler för sådana fondföretag som investerar i aktier och/eller skuldförbindelser för detta ändamål.
(17) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(6).
Artikel 1
2. I artikel 1 skall följande punkter införas: "8. I detta direktiv avses med 'överlåtbara värdepapper':
- försäljningsbara värdepapper av annat slag som ger rätt att förvärva sådana överlåtbara värdepapper genom teckning eller utbyte,
3. Artikel 19.1 a skall ersättas med följande: "a) överlåtbara värdepapper och penningmarknadsinstrument som får omsättas eller omsätts på en sådan reglerad marknad som avses i artikel 1.13 i direktivet om investeringstjänster och/eller"
- Orden "och/eller" skall läggas till i slutet av punkt d.
- skyddsnivån för andelsägare i det andra företaget för kollektiva investeringar motsvarar det skydd som ett fondföretags andelsägare har, särskilt genom att reglerna för separation av tillgångarna, in- och utlåning och försäljning av överlåtbara värdepapper och penningmarknadsinstrument som företaget inte innehar uppfyller villkoren i detta direktiv, och
f) inlåning i kreditinstitut, antingen som avistakonton eller som konton med högst 12 månaders uppsägningstid, under förutsättning att kreditinstitutet har sitt säte i en medlemsstat eller, om kreditinstitutet har sitt säte i tredje land, förutsatt att det omfattas av tillsynsregler som av behöriga myndigheter med ansvar för fondföretag anses motsvara dem som fastställs i gemenskapslagstiftningen, och/eller
- motparterna vid affärer med OTC-derivat är institutioner som omfattas av tillsyn och tillhör de kategorier som godkänts av de behöriga myndigheterna med ansvar för fondföretaget, och
- emitterats eller garanterats av en central, regional eller lokal myndighet, av en medlemsstats centralbank, av Europeiska centralbanken, av Europeiska unionen eller Europeiska investeringsbanken, av en icke-medlemsstat eller, i fråga om förbundsstater, av en av de stater som utgör förbundsstaten eller av en internationell offentlig organisation som en eller flera medlemsstater tillhör, eller
- emitterats av andra organ som tillhör de kategorier som godkänts av de behöriga myndigheterna med ansvar för fondföretaget förutsatt att investeringar i sådana instrument omfattas av ett investerarskydd som är likvärdigt med det som fastställs i första, andra eller tredje strecksatsen och att emittenten är ett bolag vars kapital och reserver uppgår till minst 10 miljoner euro och som lägger fram och offentliggör sin årsredovisning i enlighet med direktiv 78/660/EEG(7), är en enhet som inom en grupp företag som omfattar ett eller flera börsnoterade företag ägnar sig åt gruppens finansiering eller är en enhet som ägnar sig åt att finansiera värdepapperisering som omfattas av kreditförstärkning från en bank."
8. Artikel 20 skall utgå.
2. Medlemsstaterna får ge fondföretag tillstånd att använda sig av sådan teknik och sådana instrument som hänför sig till överlåtbara värdepapper och penningmarknadsinstrument på de villkor och inom de gränser medlemsstaterna föreskriver, förutsatt att sådan teknik och sådana instrument används i syfte att åstadkomma en effektiv förvaltning av värdepappersportföljen. Om denna verksamhet gäller användning av derivatinstrument skall dessa villkor och gränser överensstämma med bestämmelserna i detta direktiv.
Exponeringen skall beräknas med hänsyn till det aktuella värdet av de underliggande tillgångarna, motpartsrisken, kommande marknadsrörelser och den tid som finns tillgänglig för att lösa in positionerna. Detta skall även gälla följande stycken.
4. Senast den 13 februari 2004 skall medlemsstaterna till kommissionen överlämna fullständig information om, och eventuella förändringar i, reglerna för de metoder som används för att beräkna riskexponering enligt punkt 3, inklusive riskexponeringen för en motpart vid transaktioner med OTC-derivat. Kommissionen skall vidarebefordra denna information till övriga medlemsstater. Sådan information kommer att vara föremål för överväganden inom kontaktkommittén i enlighet med förfarandet i artikel 53.4."
Riskexponeringen mot ett fondföretags motpart vid en transaktion med OTC-derivat får inte överstiga:
2. Medlemsstaterna får höja den 5-procentsgräns som anges i första meningen i punkt 1 till högst 10 %. I den mån fondföretaget investerar mer än 5 % av fondtillgångarna i överlåtbara värdepapper och penningmarknadsinstrument med samma utgivare, får det sammanlagda innehavet av sådana investeringar inte överstiga 40 % av fondtillgångarna. Begränsningen gäller inte inlåning hos och transaktioner med OTC-derivat med finansiella institut som står under tillsyn.
- inlåning hos, och/eller
Medlemsstaterna skall till kommissionen överlämna en förteckning över de ovan nämnda kategorier av obligationer och över de kategorier av emittenter, vilka enligt gällande lag och enligt sådana tillsynsregler som avses i första stycket, beviljas tillstånd att emittera sådana obligationer som uppfyller kriterierna ovan. Till förteckningen skall fogas uppgifter om vad slags garantier som erbjudits. Kommissionen skall till övriga medlemsstater genast vidarebefordra denna information jämte de kommentarer som bedömts erforderliga samt göra informationen tillgänglig för allmänheten. Sådana underrättelser kan göras till föremål för överväganden i kontaktkommittén i enlighet med förfarandet i artikel 53.4.
Bolag som ingår i samma grupp för sammanställd redovisning enligt definitionen i direktiv 83/349/EEG(8) eller i enlighet med erkända internationella redovisningsregler räknas som ett organ vid beräkningen av gränserna i denna artikel.
1. Utan att det påverkar tillämpningen av de gränser som fastställs i artikel 25 får medlemsstaterna på följande villkor höja de gränser som anges i artikel 22 till högst 20 % för investeringar i aktier och/eller skuldförbindelser emitterade av samma organ, då fondföretagets investeringspolicy enligt fondbestämmelserna eller enligt bolagsordningen syftar till att efterbilda sammansättningen av ett visst aktieindex eller index för skuldförbindelser som är erkänt av de behöriga myndigheterna:
- Det skall offentliggöras på lämpligt vis.
13. Artikel 24 skall ersättas med följande: "Artikel 24
Medlemsstaterna får, när ett fondföretag har förvärvat andelar i fondföretag och/eller andra företag för kollektiva investeringar, medge att värdet av dessa företags tillgångar inte behöver rymmas inom de gränser som anges i artikel 22.
14. Följande artikel skall införas: "Artikel 24a
3. Om nettovärdet av ett fondföretags tillgångar tenderar att ha hög volatilitet på grund av portföljens sammansättning och förvaltningsmetoderna måste detta anges på framträdande plats i prospektet och i förekommande fall i allt övrigt reklammaterial.
1. Tredje strecksatsen skall ersättas med följande: "- 25 % av andelarna i ett enskilt fondföretag och/eller annat företag för kollektiva investeringar enligt artikel 1.2 första och andra strecksatsen,"
17. I artikel 25.3 a, b och c skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
Medlemsstaterna får, med beaktande av principen om riskspridning, tillåta nyligen auktoriserade fondföretag att under en tid av högst sex månader från auktorisationsdagen avvika från artiklarna 22, 22a, 23 och 24."
1. Utöver de funktioner som finns angivna i artikel 53.1 kan kontaktkommittén också sammanträda som en föreskrivande kommitté i enlighet med artikel 5 i beslut 1999/468/EG(9) för att bistå kommissionen med tekniska ändringar i detta direktiv på följande områden:
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 2
b) en översyn av direktivets tillämpningsområde vad gäller olika produkttyper (till exempel institutionella fonder, fastighetsfonder, matarfonder och hedgefonder); översynen bör särskilt inriktas på storleken på marknaden för sådana fonder, eventuell reglering av sådana fonder i medlemsstaterna och bedömning av behovet av ytterligare harmonisering av dessa fonder,
e) en analys av konkurrenssituationen mellan fonder som förvaltas av förvaltningsföretag respektive investeringsföretag som sköter förvaltningen själva.
Artikel 3
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 5
av den 12 januari 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
efter samråd med Rådgivande kommittén för statligt stöd, och
(2) Genom förordning (EG) nr 994/98 bemyndigas också kommissionen att i enlighet med artikel 87 i fördraget förklara att stöd som är förenliga med den av kommissionen för varje medlemsstat godkända regionalstödskartan är förenliga med den gemensamma marknaden och undantagna från anmälningsskyldigheten enligt artikel 88.3 i fördraget.
(5) Små och medelstora företag spelar en avgörande roll för att skapa arbetstillfällen och medverkar allmänt till social stabilitet och en dynamisk ekonomi. Brister i marknadens sätt att fungera kan emellertid hämma deras utveckling. De har ofta svårigheter att få tillgång till kapital och krediter till följd av obenägenheten att ta risker på vissa finansiella marknader och de begränsade garantier som dessa företag kan erbjuda. De små och medelstora företagens begränsade resurser kan också inskränka deras möjligheter att få tillgång till information, särskilt om ny teknik och nya marknader. Mot bakgrund av dessa överväganden bör det stöd som genom denna förordning undantas från anmälningsskyldigheten syfta till att underlätta utvecklingen av verksamheten i de små och medelstora företagen, under förutsättning att stödet inte påverkar handeln i negativ riktning i en omfattning som strider mot det gemensamma intresset.
(8) För att vid tillämpningen av denna förordning eliminera olikheter som kan medföra snedvridningar av konkurrensen och för att underlätta samordningen mellan olika initiativ inom gemenskapen och på nationell nivå som rör små och medelstora företag samt av hänsyn till administrativ klarhet och rättssäkerhet, bör definitionen av små och medelstora företag i denna förordning vara densamma som fastställs i kommissionens rekommendation 96/280/EG av den 3 april 1996 om definitionen av små och medelstora företag(5). Den definitionen används också i gemenskapens riktlinjer för statligt stöd till små och medelstora företag(6).
(11) Med hänsyn till skillnaderna mellan små företag och medelstora företag bör olika stödtak fastställas för små företag respektive medelstora företag.
(14) Genom denna förordning bör stöd till små och medelstora företag undantas från anmälningsskyldigheten oberoende av var företagen är belägna. Investeringar och skapande av arbetstillfällen kan bidra till den ekonomiska utvecklingen i gemenskapens mindre gynnade regioner. Små och medelstora företag i dessa regioner har strukturella nackdelar på grund av sin lokalisering och svårigheter på grund av sin begränsade storlek. De bör därför beviljas högre stödtak.
(17) Med hänsyn till behovet att uppnå balans mellan minsta möjliga snedvridning av konkurrensen inom den understödda sektorn och denna förordnings mål bör enskilda stöd som överskrider ett fastställt maximibelopp inte medges undantag enligt denna förordning, oavsett om de omfattas av en stödordning som har beviljats undantag enligt denna förordning eller inte.
(20) I syfte att säkerställa insyn och effektiv kontroll i enlighet med artikel 3 i förordning (EG) nr 994/98 är det lämpligt att utarbeta ett standardformulär som medlemsstaterna bör använda för att förse kommissionen med sammanfattande information för offentliggörande i Europeiska gemenskapernas officiella tidning, varje gång en stödordning genomförs eller ett enskilt stöd som inte täcks av någon sådan stödordning beviljas enligt denna förordning. Av samma skäl är det lämpligt att fastställa regler för de register som medlemsstaterna bör föra över stöd som har beviljats undantag enligt denna förordning. Beträffande den årliga rapport som medlemsstaterna är skyldiga att överlämna till kommissionen, är det lämpligt att kommissionen fastställer de närmare kraven på rapportens utformning, inbegripet information i elektronisk form, då den teknik som krävs för detta är allmänt tillgänglig.
Artikel 1
2. Denna förordning får inte tillämpas på
c) stöd som förutsätter att inhemska produkter används på bekostnad av importerade produkter.
I denna förordning används följande beteckningar med de betydelser som här anges:
c) investering i materiella tillgångar: investering i materiella anläggningstillgångar som hänför sig till skapandet av en ny anläggning, utvidgning av en existerande anläggning, eller igångsättande av en verksamhet som innebär en grundläggande förändring av en existerande anläggningsprodukt eller produktionsprocess (genom rationalisering, omställning eller modernisering). En investering i anläggningstillgångar som genomförs i form av övertagande av en anläggning som har lagts ned eller som skulle ha lagts ned om den inte hade förvärvats skall också betraktas som en materiell investering.
f) stödnivå netto: stödbeloppet efter avdrag för skatt i procent av projektets stödberättigande kostnader.
Förutsättningar för undantag
a) varje stöd som skulle kunna beviljas inom ramen för stödordningen uppfyller samtliga villkor i denna förordning,
Artikel 4
2. Stödnivån brutto får inte överskrida
3. Om investeringen äger rum i områden som är berättigade till regionalstöd får stödnivån inte överstiga det tak för regionalt investeringsstöd som fastställts i den karta som kommissionen har godkänt för varje medlemsstat med mer än
De högre regionala stödtaken skall endast gälla om stödet beviljas på villkor att investeringen bibehålls i den stödmottagande regionen under minst fem år och att stödmottagarens bidrag till finansieringen av investeringen uppgår till minst 25 %.
6. Om stödet beräknas på grundval av skapade arbetstillfällen skall stödbeloppet uttryckas i procent av lönekostnaderna för den sysselsättning som skapats under en tvåårsperiod enligt följande villkor:
c) Den skapade sysselsättningen måste bibehållas under en period av minst fem år.
Stöd till små och medelstora företag som uppfyller följande villkor skall vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget:
Artikel 6
a) de totala stödberättigande kostnaderna för hela projektet är minst 25 miljoner euro, och
b) det totala stödbeloppet brutto är minst 15 miljoner euro.
Stöd får beviljas undantag enligt denna förordning endast om medlemsstaten innan arbetet på det berörda projektet inleds
Artikel 8
2. Stöd som undantas genom denna förordning får inte kumuleras med något annat statligt stöd i den mening som avses i artikel 87.1 i fördraget eller med annan gemenskapsfinansiering, i förhållande till samma stödberättigande kostnader, om en sådan kumulering skulle leda till en högre stödnivå än den som fastställs i denna förordning.
1. Vid genomförandet av en stödordning eller vid beviljandet av ett enskilt stöd som inte omfattas av någon stödordning, skall medlemsstaterna, om stödordningen eller stödet är undantaget enligt denna förordning, till kommissionen inom tjugo arbetsdagar överlämna en sammanfattning av uppgifterna om stödordningen eller det enskilda stödet enligt det formulär som anges i bilaga II för offentliggörande i Europeiska gemenskapernas officiella tidning.
Artikel 10
Kommissionens förordning (EG) nr 283/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Följaktligen bör förordning (EG) nr 2734/2000 ändras.
(6) Följaktligen bör förordning (EG) nr 562/2000 ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"1. Trots vad som sägs i artikel 4.2 g i förordning (EG) nr 562/2000 skall den maximala vikten för de slaktkroppar som avses i ovannämnda bestämmelse vara 430 kg. Dock
Artikel 2
"d) De har försetts med etiketter i enlighet med det system som införs genom Europaparlamentets och rådets förordning (EG) nr 1760/2000(7), samt för avtal som sluts från och med den 12 februari 2001 även de uppgifter som anges i artikel 13.5 i den förordningen."
Artikel 3
av den 18 april 2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) Vid fastställandet av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung är det nödvändigt att ange de djurarter i vilka restmängder kan förekomma, vilka mängder som kan förekomma i var och en av de relevanta vävnaderna från det behandlade djuret (målvävnad) samt vilket slag av restmängd som är relevant vid övervakningen av restmängder (restmarkör).
(6) Tiamylal och Tiopentalnatrium skall införas i bilaga II till förordning (EEG) nr 2377/90.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 14 maj 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I artikel 24 i förordning (EG) nr 104/2000, som upphävde rådets förordning (EEG) nr 3759/92(2) med verkan från och med den 1 januari 2001, föreskrivs att ett schablonmässigt stöd på vissa villkor skall beviljas producentorganisationer som återtar produkter som förtecknas i bilaga IV till den förordningen.
(4) Det bör fastställas bestämmelser som producentorganisationerna skall följa när det gäller schablonmässigt stöd.
(7) För att säkerställa produkternas kvalitet och underlätta deras avsättning på marknaden bör det fastställas vilka minimikrav för beredningen som skall vara tillgodosedda och vilka villkor som skall gälla för lagring och återförande till marknaden av de bearbetade produkterna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
KAPITEL II
Villkoren i artiklarna 1-4 och artikel 7 i förordning (EG) nr 2509/2000 skall i tillämpliga delar gälla för beviljande av schablonersättning.
För alla producentorganisationer som medlemsstaten har erkänt skall det fastställas ett schablonvärde vid fiskeårets början på grundval av de genomsnittliga inkomster som i samband med dessa avsättningar uppnåtts och konstaterats i de berörda medlemsstaterna under sex månader innan detta schablonvärde fastställs. Värdet skall emellertid ändras om väsentliga och bestående inkomstvariationer konstateras på medlemsstatens marknad.
Artikel 5
3. Följande skall betraktas som tekniska kostnader:
c) Kostnader för material vid direktförpackning.
4. De ekonomiska kostnaderna skall utgöras av ett schablonbelopp på 10 euro per ton för 2001. Därefter skall schablonbeloppet justeras årligen enligt den räntesats som årligen fastställs i enlighet med artikel 5 i rådets förordning (EEG) nr 1883/78(11).
Bestämmelserna i artikel 3.1 och 3.2 samt artikel 4 i förordning (EG) nr 2814/2000 skall i tillämpliga delar gälla för beviljande av schablonbidrag.
KAPITEL IV
1. Ansökningar om utbetalning av schablonmässigt stöd skall av producentorganisationerna överlämnas till de behöriga myndigheterna i medlemsstaten inom fyra månader från det aktuella fiskeårets slut. Ansökningarna skall minst innehålla de uppgifter som anges i bilagan.
4. De nationella myndigheterna skall betala ut det schablonmässiga stödet senast åtta månader efter fiskeårets slut. Varje medlemsstat skall underrätta övriga medlemsstater och kommissionen om namn på och adress till det organ som utsetts att betala ut det schablonmässiga stödet.
2. Producentorganisationerna skall se till att stödmottagarna för lagerbokföring i enlighet med den förlaga som finns i bilagan.
Medlemsstaterna skall underrätta kommissionen om de åtgärder som vidtagits för tillämpningen av den här förordningen så snart de antagits, och i vart fall senast den 1 juli 2001. De skall senast den 1 juli 2001 underrätta kommissionen om redan gällande åtgärder på det område som omfattas av artikel 9.1.
Artikel 12
om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati
med beaktande av kommissionens förslag(1),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) Sedan 1990 har gemenskapen beslutat om en rad åtgärder för att skydda människor och djur mot BSE-risken. Dessa åtgärder grundar sig på skyddsbestämmelserna i direktiven om kontrollåtgärder på veterinärområdet. Med hänsyn till omfattningen av den hälsorisk som människor och djur utsätts för genom vissa typer av TSE är det lämpligt att anta särskilda bestämmelser om förebyggande, kontroll och utrotning av dessa.
(5) Dessa bestämmelser bör gälla produktion och avyttring av levande djur och animaliska produkter. De behöver däremot inte gälla kosmetiska eller medicinska produkter, medicintekniska produkter, deras utgångsmaterial eller mellanprodukter, för vilka andra särskilda bestämmelser gäller, särskilt avseende förbud mot användning av vissa typer av riskmaterial. De bör inte heller gälla animaliska produkter som inte innebär någon hälsorisk för människor och djur eftersom de är avsedda att användas till annat än livsmedel, foder eller gödningsmedel. Det är däremot nödvändigt att säkerställa att animaliska produkter som inte omfattas av denna förordning hålls åtskilda från dem som omfattas av förordningen, om de inte uppfyller minst samma hälsovillkor som de sistnämnda.
(8) Medlemsstaterna bör införa utbildningsprogram för dem som har till uppgift att förebygga och bekämpa TSE, liksom för veterinärer, jordbrukare och personer som har hand om transport, avyttring och slakt av livsmedelsproducerande djur.
(11) Åtgärder bör vidtas för att förhindra att TSE överförs till människor och djur genom förbud mot att utfodra vissa kategorier djur med vissa kategorier djurprotein, samt genom förbud mot att använda vissa material från idisslare i livsmedel. Dessa förbud bör stå i proportion till de risker det handlar om.
(14) Medlemsstaterna bör upprätta beredskapsplaner i vilka de nationella åtgärder som skall vidtas vid ett utbrott av BSE anges. Beredskapsplanerna bör godkännas av kommissionen. Bestämmelser bör införas för att kunna utsträcka denna bestämmelse till att gälla andra typer av TSE än BSE.
(17) För att säkerställa att reglerna om förebyggande, kontroll och utrotning av TSE respekteras är det lämpligt att ta prover för laboratorietester på grundval av ett på förhand fastställt protokoll som kan ge en fullständig epidemiologisk bild av läget när det gäller TSE. För att garantera att testförfarandena och testresultaten är enhetliga bör referenslaboratorier inrättas, nationellt och på gemenskapsnivå; därtill måste det införas tillförlitliga vetenskapliga metoder, bland annat specifika snabbtest för TSE. Man bör i möjligaste mån använda snabbtest.
(20) Det bör föreskrivas att denna förordning skall ses över när nya vetenskapliga uppgifter blir tillgängliga.
(23) I syfte att genomföra denna förordning bör förfaranden fastställas för ett nära och effektivt samarbete mellan kommissionen och medlemsstaterna inom Ständiga veterinärkommittén, Ständiga foderkommittén och Ständiga livsmedelskommittén.
KAPITEL I
Tillämpningsområde
a) kosmetiska, medicinska eller medicintekniska produkter, eller utgångsmaterial och mellanprodukter till dessa,
d) levande djur som används vid eller är avsedda för forskning.
För att undvika korskontaminering eller substitution av levande djur eller animaliska produkter som avses i artikel 1.1, med de animaliska produkter som avses i artikel 1.2 a-1.2 c eller de levande djur som avses i artikel 1.2 d, skall de hållas permanent åtskilda, såvida inte dessa levande djur eller dessa animaliska produkter har framställts under åtminstone likvärdiga hälsoskyddsvillkor när det gäller TSE.
Definitioner
b) avyttring: all verksamhet som har till syfte att sälja levande djur eller animaliska produkter som omfattas av denna förordning, till tredje man inom gemenskapen, eller varje annan form av överlåtelse mot eller utan betalning till en sådan tredje man, eller lagring i syfte att senare tillhandahålla en sådan tredje man produkterna.
e) behörig myndighet: den centrala myndighet i en medlemsstat som har till uppgift att se till att kraven i denna förordning efterlevs, eller varje annan myndighet till vilken den centrala myndigheten har delegerat nämnda uppgift, särskilt för foderkontroll. Denna definition skall också, i förekommande fall, omfatta motsvarande myndighet i tredje land.
h) djur som misstänks vara smittade med TSE: levande, slaktade eller döda djur som uppvisar eller har uppvisat neurologiska eller beteendemässiga störningar eller ett gradvis försämrat allmäntillstånd som har samband med en störning i centrala nervsystemet och för vilka ingen alternativ diagnos kan fastställas på grundval av information som inhämtats på grundval av en klinisk undersökning, svar på behandling, obduktion eller laboratorieanalys före eller efter djurets död. Alla nötkreatur som har gett positivt resultat i ett snabbtest för bovin spongiform encefalopati (BSE) skall också misstänkas vara smittade med BSE.
k) gödningsmedel: varje ämne som innehåller animaliska produkter som används på mark för att främja tillväxten. Det får innehålla rötningsrester från biogasproduktion eller kompostering.
2. De särskilda definitionerna i bilaga I skall också gälla.
Skyddsåtgärder
KAPITEL II
Klassificering
2. Ett beslut om att fatta ett avgörande om varje ansökan för att klassificera den medlemsstat eller det tredje land eller den region i medlemsstaten eller det tredje landet som har lämnat in ansökan såsom hörande till någon av kategorierna i kapitel C i bilaga II, skall fattas med beaktande av de kriterier och potentiella riskfaktorer som anges i punkt 1, i enlighet med det förfarande som avses i artikel 24.2.
3. Om kommissionen finner att den information som en medlemsstat eller ett tredje land har lämnat i enlighet med kapitlen A och B i bilaga II är otillräcklig eller oklar, kan den i enlighet med det förfarande som avses i artikel 24.2 fastställa BSE-status för den berörda medlemsstaten eller det berörda tredje landet på grundval av en fullständig riskanalys.
Detta screeningförfarande kan även utnyttjas av de medlemsstater eller tredje länder som vill att kommissionen - enligt det förfarande som avses i artikel 24.2 - skall godkänna den klassificering som de gjort på denna grund.
5. Medlemsstaterna skall utan dröjsmål till kommissionen anmäla alla epidemiologiska bevis eller annan information som skulle kunna leda till förändringar i deras BSE-status, särskilt resultaten av de övervakningsprogram som föreskrivs i artikel 6.
7. Ett beslut får antas i enlighet med det förfarande som avses i artikel 24.2 om att ändra BSE(klassificeringen för en medlemsstat eller ett tredje land eller någon av deras regioner i enlighet med resultaten av de kontroller som föreskrivs i artikel 21.
FÖREBYGGANDE AV TSE
1. Varje medlemsstat skall genomföra ett årligt övervakningsprogram för BSE och scrapie i enlighet med kapitel A i bilaga III. Ett screeningförfarande med hjälp av snabbtest skall ingå i detta program.
3. Alla officiella undersökningar och laboratorieprov skall registreras enligt kapitel B.1 bilaga III.
Förbud avseende foder
3. Punkterna 1 och 2 skall tillämpas utan att det påverkar tillämpningen av punkt 2 i bilaga IV.
5. Tillämpningsföreskrifterna för denna artikel, inbegripet reglerna om förebyggande av korskontaminering och om de metoder för provtagning och provanalys som krävs för att kontrollera att denna artikel efterlevs, skall antas enligt det förfarande som avses i artikel 24.2.
1. Det specificerade riskmaterialet skall avlägsnas och destrueras i enlighet med punkterna 2, 3, 4 och 8 i bilaga V.
De medlemsstater som godkänner detta alternativa test skall underrätta de övriga medlemsstaterna och kommissionen om detta.
5. Trots vad som sägs i punkterna 1-4 kan ett beslut antas i enlighet med det förfarande som avses i artikel 24.2 om den dag då bestämmelserna i artikel 7.1 skall börja gälla eller i förekommande fall i tredje land om den dag förbudet skall träda i kraft mot användning av proteiner som härrör från däggdjur i foder för idisslare i samtliga länder eller regioner som placerats i kategori 3 eller 4, i syfte att begränsa tillämpningen av denna artikel till djur som har fötts före denna dag i dessa länder eller regioner.
Artikel 9
2. Skallben och kotpelare från nötkreatur, får och getter från länder eller regioner som är placerade i kategori 2, 3, 4 eller 5 får inte användas för framställning av mekaniskt urbenat kött.
Artikel 10
2. För att de utbildningsprogram som avses i punkt 1 skall kunna genomföras effektivt får gemenskapen bevilja ekonomiskt stöd. Beloppet för ett sådant stöd skall bestämmas enligt det förfarande som avses i artikel 24.2.
Artikel 11
Medlemsstaterna skall regelbundet underrätta övriga medlemsstater och kommissionen om anmälda fall av TSE.
Åtgärder vid misstänkta fall
Om man misstänker BSE hos ett får eller en get på en anläggning i en medlemsstat på grundval av objektiva faktorer såsom resultaten av ett test som på ett praktiskt sätt kan göra åtskillnad mellan olika typer av TSE, skall alla övriga får och getter på anläggningen vara föremål för officiella restriktioner vad avser förflyttning i avvaktan på att resultaten av undersökningen blir tillgängliga.
2. Om den behöriga myndigheten beslutar att det inte kan uteslutas att ett djur har smittats av TSE, skall djuret - om det fortfarande är vid liv - avlivas; dess hjärna, liksom alla övriga vävnader som den behöriga myndigheten bestämmer, skall avlägsnas och skickas till ett officiellt godkänt laboratorium, det nationella referenslaboratoriet enligt artikel 19.1 eller gemenskapens referenslaboratorium enligt artikel 19.2, för att undersökas där enligt de testmetoder som anges i artikel 20.
Artikel 13
a) Samtliga delar av det smittade djurets kropp skall destrueras fullständigt i enlighet med bilaga V, med undantag för det material som skall bevaras för registren i enlighet med kapitel B.III.2 i bilaga III.
En medlemsstat får, trots bestämmelserna i detta stycke, tillämpa andra åtgärder som erbjuder motsvarande skyddsnivå, om dessa åtgärder har godkänts enligt det förfarande som avses i artikel 24.2.
3. De medlemsstater som har genomfört ett alternativt system som erbjuder likvärdiga garantier enligt artikel 12.1 femte stycket får, enligt det förfarande som avses i artikel 24.2 och med avvikelse från kraven i punkterna 1 b och 1 c, undantas från skyldigheten att tillämpa det officiella förbudet mot förflyttning av djuren och från kravet på att avliva och destruera djuren.
6. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
1. Medlemsstaterna skall - i enlighet med de allmänna kriterierna i gemenskapens bestämmelser för kontroll av djursjukdomar - utarbeta riktlinjer som specificerar vilka nationella åtgärder som skall genomföras och ange behörighet och ansvar om TSE-fall bekräftas.
AVYTTRING OCH EXPORT
1. Avyttring eller i förekommande fall export av nötkreatur, får eller getter och deras sperma, embryon och ägg skall omfattas av de villkor som anges i bilaga VIII eller, vid import, de villkor som anges i bilaga IX. De levande djuren och deras embryon och ägg skall åtföljas av de relevanta hälsointyg som föreskrivs i gemenskapslagstiftningen i enlighet med artikel 17 eller, vid import, i enlighet med artikel 18.
Artikel 16
a) Animaliska produkter som omfattas av bestämmelserna i artikel 15, särskilt sperma, embryon och ägg.
iii) Värmebehandlad konsumtionsmjölk enligt definitionen i direktiv 92/46/EEG.
vi) Gelatin i den mening som avses i direktiv 92/118/EEG som härrör från hudar och skinn enligt punkt v.
3. Animaliska produkter som innehåller material från nötkreatur med ursprung i en medlemsstat, en region i en medlemsstat eller ett tredje land som placerats i kategori 5 får inte avyttras utom i de fall då de härrör från
Animaliska produkter får inte skickas från en medlemsstat eller en region i en medlemsstat som placerats i kategori 5, från en annan medlemsstat eller importeras från ett tredje land som placerats i kategori 5. Detta förbud gäller inte sådana animaliska produkter som avses i kapitel C i bilaga VIII och som uppfyller kraven i kapitel C i bilaga VIII. De skall åtföljas av ett hälsointyg som utfärdats av en officiell veterinär som intygar att de framställts i enlighet med denna förordning.
6. För import till gemenskapen skall animaliska produkter uppfylla kraven i kapitlen A, C, F och G i bilaga IX.
Enligt det förfarande som avses i artikel 24.2 skall de hälsointyg som avses i bilaga F till direktiv 64/432/EEG och i modellerna II och III i bilaga E till rådets direktiv 91/68/EEG, samt de lämpliga hälsointyg som föreskrivs i gemenskapslagstiftningen om handel med sperma, ägg och embryon från nötkreatur, får eller getter vid behov kompletteras med en uppgift om kategori med angivande av den klassificering av medlemsstaten eller ursprungsregionen som gjorts enligt artikel 5.
Lämpliga hälsointyg för import som föreskrivs i gemenskapslagstiftningen skall, enligt det förfarande som avses i artikel 24.2, kompletteras med de särskilda kraven i bilaga IX när det gäller tredje länder som klassificerats i en kategori i enlighet med artikel 5, så snart detta beslut om klassificering har antagits.
Artikel 19
2. Gemenskapens referenslaboratorium, dess behörighet och uppgifter fastställs i kapitel B i bilaga X.
1. Provtagning och laboratorieundersökningar för att fastställa förekomst av TSE skall genomföras enligt de metoder och protokoll som anges i kapitel C i bilaga X.
Gemenskapskontroller
2. Gemenskapskontrollerna vad avser tredje land skall ske i enlighet med artiklarna 20 och 21 i direktiv 97/78/EG.
Artikel 22
2. Resultaten av en avgörande statistisk undersökning, som under övergångsperioden utförs i enlighet med bestämmelserna i artikel 5.3, skall utnyttjas för att bekräfta eller vederlägga slutsatserna från den riskanalys som avses i artikel 5.1, varvid de klassificeringskriterier som fastställts av Internationella byrån för epizootiska sjukdomar skall beaktas.
Artikel 23
Enligt det förfarandet skall övergångsbestämmelser antas för en period på högst två år för att möjliggöra en övergång från nuvarande ordning till den ordning som fastställs i denna förordning.
1. Kommissionen skall biträdas av Ständiga veterinärkommittén. I frågor som uteslutande rör foder skall kommissionen dock biträdas av Ständiga foderkommittén, och i frågor som uteslutande rör livsmedel skall kommissionen biträdas av Ständiga livsmedelskommittén.
3. Varje kommitté skall själva anta sin arbetsordning.
De relevanta vetenskapliga kommittéerna skall höras i alla frågor som omfattas av tillämpningsområdet för denna förordning och som kan ha konsekvenser för folkhälsan.
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om tillämpningsföreskrifter för rådets förordning (EG) nr 1493/1999 om framtagning av uppgifter för produktinformation och marknadsuppföljning inom vinsektorn och om ändring av förordning (EG) nr 1623/2000
med beaktande av rådets förordning (EG) nr 1493/1999 av 17 maj 1999 om den gemensamma organisationen av marknaden för vin(1), senast ändrad genom förordning (EG) nr 2826/2000(2), särskilt artiklarna 23, 33 och 73 i denna, och
(2) I samma artikel föreskrivs att medlemsstaterna även får kräva att försäljare av druvor varje år skall deklarera vilka mängder som saluförts från den senaste skörden.
(5) Medlemsstaterna får själva närmare besluta om på vilket sätt företagen skall lämna de uppgifter som skall ingå i deklarationen, men för att underlätta tillämpningen av denna förordning bör det föreskrivas att uppgifterna skall lämnas i tabellform. Det är också nödvändigt att fastställa tidsfrister inom vilka medlemsstaterna skall sammanställa och överlämna de insamlade uppgifterna till kommissionen, samt att ange på vilket sätt de skall överlämnas.
(8) Påföljdssystemet bör tillåta en tillräcklig grad av proportionalitet för de av vinproducenternas deklarationer som vid kontroll har visats vara ofullständiga eller oriktiga. Påföljden bör anpassas efter de rättelser som görs i en deklaration.
(11) Vissa uppgifter om vinmarknaden är nödvändiga för marknadsuppföljningen. Utöver uppgifter från sammanställningar av de olika deklarationerna måste även tillgängliga mängden, deras användning samt vinpriser uppges. Därför bör det föreskrivas att medlemsstaterna skall samla in uppgifterna och överlämna dem till kommissionen senast vissa angivna datum.
(14) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för vin.
Denna förordning gäller tillämpningsföreskrifter för förordning (EG) nr 1493/1999, främst när det gäller framtagning av uppgifter som ökar produktkunskapen och som kan användas för marknadsuppföljning inom vinsektorn.
I förekommande fall får medlemsstaterna tillåta att en deklaration lämnas per jordbruksföretag.
b) Skördare vars jordbruksföretag omfattar mindre än 10 ar vinodlingsareal och som varken har sålt eller kommer att sälja någon del av sin produktion i någon form.
ii) den mängd druvor som levereras,
3. Med undantag från punkt 1 första stycket, och utan att detta påverkar de skyldigheter som följer av artikel 4, får medlemsstaterna undanta följande personer från skyldigheten att lämna skördedeklarationer:
Artikel 3
2. Medlemsstaterna får föreskriva att fysiska eller juridiska personer eller sammanslutningar av sådana personer, inbegripet vinkooperativ, som före de tidpunkter som anges i artikel 11.1 har behandlat eller salufört produkter i tidigare produktionsled än vin under innevarande vinår, till de behöriga myndigheterna skall lämna in behandlings- eller saluföringsdeklarationer som minst skall innehålla uppgifterna enligt tabell C.
5. Beträffande fysiska eller juridiska personer eller sammanslutningar av sådana personer, som överlåter vinprodukter i produktionsleden före vin, skall medlemsstaterna vidta nödvändiga åtgärder för att se till att producenter som skall lämna deklarationer har tillgång till de uppgifter som skall ingå.
I dessa fall skall de behöriga myndigheter som har utsetts av medlemsstaten själva fylla i de deklarationer som avses i denna artikel med uppgifter om arealen som bygger på uppgifterna i vinodlingsregistret.
Medlemsstater med en årlig vinproduktion av högst 25000 hektoliter får emellertid utöver detaljister undanta även andra handelsidkare som innehar små lager från skyldigheten att lämna de deklarationer som avses i första stycket, förutsatt att de behöriga myndigheterna kan ge kommissionen en statistisk uppskattning av dessa lagers storlek i medlemsstaten.
3. Den deklaration som avses i punkt 1 skall innehålla minst de uppgifter som framgår av tabell D i bilagan.
Formulären behöver inte innehålla någon uttrycklig hänvisning till areal om medlemsstaten med säkerhet kan bestämma denna med hjälp av andra uppgifter som lämnas i deklarationen eller i vinodlingsregistret, särskilt produktionsarealen och jordbruksföretagets totala skörd.
De skall underrätta kommissionen om dessa åtgärder och översända de formulär som utarbetas enligt första stycket.
- fått alla de uppgifter som skall anges i deklarationerna enligt kapitlen I och II från andra administrativa handlingar får undanta aktörerna i fråga från skyldigheten att lämna in en eller flera av deklarationerna.
- fått alla de uppgifter som skall anges i deklarationerna enligt kapitel III från andra administrativa handlingar får undanta aktörerna i fråga från skyldigheten att lämna in deklarationerna.
När det gäller den deklaration som avses i artikel 4 skall emellertid endast sådant vin betraktas som "annat vin" enligt första stycket som enbart skall användas för framställning av vinsprit med skyddad ursprungsbeteckning eller sådan obligatorisk destillation som avses i artikel 28 i förordning (EG) nr 1493/1999.
Medlemsstaterna får dock föreskriva att mängderna skall uttryckas i deciton i stället för i hektoliter i de deklarationer som avses i artikel 2.
Artikel 10
1. De deklarationer som avses i artiklarna 2 och 4 skall lämnas senast den 10 december. Medlemsstaterna får emellertid fastställa ett eller flera tidigare datum. De får dessutom fastställa ett visst datum vid vilket de kvantiteter som innehas skall tas med i deklarationen.
Personer som skall lämna in skörde-, produktions-, saluförings- och/eller behandlings- eller lagerdeklarationer och som inte har lämnat in dessa vid de tidpunkter som anges i artikel 11 skall, utom i fall av force majeure, inte omfattas av de åtgärder som föreskrivs i artiklarna 24, 29, 30, 34 och 35 i förordning (EG) nr 1493/1999 för innevarande och närmast därpå följande vinår.
1. Personer som skall lämna in skörde-, produktions-, saluförings-, behandlings- eller lagerdeklarationer och som lämnar in deklarationer som de behöriga myndigheterna i medlemsstaterna finner ofullständiga eller oriktiga får endast omfattas av de åtgärder som avses i artiklarna 24, 29, 30, 34 och 35 i förordning (EG) nr 1493/1999 om de uppgifter som saknas eller som är oriktiga inte är avgörande för ett korrekt genomförande av åtgärderna i fråga.
- samma procentsats som det konstaterade felet om felet medför att den deklarerade volymen justeras med 5 % eller mindre,
Om den oriktighet som fastställts i deklarationen kan hänföras till uppgifter från andra aktörer eller anslutna vilkas namn finns med i de föreskrivna handlingarna och inte kan kontrolleras i förväg av deklaranten skall stödet endast minskas med procentsatsen för justeringen.
Dessa priser skall inte betalas om felet medför att den deklarerade volymen justeras med mer än 20 %, vare sig för vinåret i fråga eller för det därpå följande vinåret.
Artikel 14
b) En sammanställning på nationell nivå av de lagerdeklarationer som avses i artikel 6 i denna förordning.
e) En provisorisk försörjningsbalans för senast föregående vinår och en slutlig försörjningsbalans för det näst senaste vinåret.
2. För varje produktionsområde skall medlemsstaterna välja plats för prisnoteringen.
Artikel 16
b) senast den 30 november, en sammanställning av lagerdeklarationerna enligt artikel 14 b,
e) senast den 15 februari, en sammanställning av produktionsdeklarationerna enligt artikel 14 a, eller en preliminär sammanställning. I det senare fallet skall det slutliga resultatet meddelas senast den 15 april.
- Definitionen av de fastställda produktionsområdena.
- Bestämmelserna för prisnotering.
Medlemsstaterna skall underrätta kommissionen om alla nya omständigheter av betydelse som i nämnvärd grad kan påverka den bedömning av tillgängliga mängder och deras användning som görs på grundval av den slutgiltiga informationen från tidigare år.
Artikel 19
Artikel 74.4 i förordning (EG) nr 1623/2000 skall ersättas med följande: "4. Interventionsorganet skall från producenten återvinna ett belopp som motsvarar en del eller hela det stöd som betalats ut till destillatören i de fall producenten inte uppfyller kraven i gemenskapens bestämmelser för destillationen i fråga, och orsaken är något av följande:
b) Producenten har lämnat in en deklaration enligt punkt a ovan som medlemsstatens behöriga myndigheter anser vara ofullständig eller felaktig, och de uppgifter som saknas eller är felaktiga anses vara av väsentlig betydelse för tillämpningen av den berörda åtgärden.
Hela det stöd som har betalats ut till destillatören skall återvinnas."
Kommissionens förordning (EEG) nr 2396/84(8) och (EG) nr 1294/96(9) upphör att gälla.
Kommissionens förordning (EG) nr 1322/2001
(Text av betydelse för EES)
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), senast ändrad genom kommissionens förordning (EG) nr 807/2001(2), särskilt artikel 6, 7 och 8 i denna, och
(2) Gränsvärden bör fastställas först efter det att Kommittén för veterinärmedicinska läkemedel har granskat all relevant information beträffande säkerheten med restmängder av ämnet i fråga för den som konsumerar livsmedel med animaliskt ursprung samt restmängdernas påverkan på den industriella bearbetningen av livsmedel.
(5) För veterinärmedicinska läkemedel som är avsedda för äggläggande fåglar, mjölkdjur eller honungsbin, måste gränsvärden även fastställas för ägg, mjölk eller honung.
(8) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
Bilaga I och III till förordning (EEG) nr 2377/90 skall ändras i enlighet med bilagan till den här förordningen.
Kommissionens förordning (EG) nr 1637/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) ICES har utvidgat sin förteckning över de arter vilkas fångst i nordöstra Atlanten skall inläggas i ICES:s databas och där medlemsstaterna när det gäller dessa ytterligare arter således skall uppmuntras att lämna tillgänglig fångststatistik.
(6) De åtgärder, som föreskrivs i denna förordning står i överensstämmelse med yttrandet från Ständiga kommittén för jordbruksstatistik inrättad genom rådets förordning 72/279/EEG(2).
Bilaga I till förordning (EEG) nr 3880/91 skall ersättas med bilaga I till denna förordning.
Artikel 3
av den 16 augusti 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I artikel 58 i kommissionens förordning (EG) nr 1623/2000 av den 25 juli 2000 om tillämpningsföreskrifter för rådets förordning (EG) nr 1493/1999 om den gemensamma organisationen av marknaden för vin, vad beträffar marknadsmekanismerna(3), senast ändrad genom förordning (EG) nr 1282/2001(4), föreskrivs vinproducenters skyldigheter vid levererans av resterande kvantiteter till destillerier. Erfarenheten visar att tidsfristen bör senareläggas.
(4) Förvaltningskommittén för vin har inte avgivit något yttrande inom den tid som dess ordförande har bestämt.
Förordning (EG) nr 1623/2000 ändras på följande sätt:
a) Punkterna 1 och 2 skall ersättas med följande: "1. För bordsvin och vin som lämpar sig för framställning av bordsvin skall destillationen enligt artikel 29 i förordning (EG) nr 1493/1999 börja från och med den 16 oktober varje vinår.
3. Artikel 86 första stycket skall ersättas med följande: "Kommissionen skall enligt förfarandet i artikel 75 i förordning (EG) nr 1493/1999 kvartalsvis inleda flera anbudsinfordringar som var och en skall omfatta minst 50000 hektoliter vinalkohol, och kvartalsvis tillsammans högst 600000 hektoliter hundraprocentig alkohol, för export till vissa tredje länder för slutlig användning endast inom bränslesektorn."
b) per dag efter den överskridna exporttidsfristen till 0,33 % av återstående belopp, efter avdrag av de tidigare 15 %."
6. Artikel 98 skall ändras på följande sätt:
a) får anbudsgivare eller godkända företag enligt artikel 92 erhålla prover av den tilldelade alkoholen,
7. Artikel 100.2 c skall ersättas med följande: "c) Beträffande alkohol som vid offentlig auktion tilldelas för nya industriella användningsområden i syfte att användas som bioetanol inom gemenskapens bränslesektor och som måste rektifieras före den slutliga användningen, skall en användning för de föreskrivna ändamålen anses vara fullständig när minst 90 % av de totala alkoholkvantiteter som avhämtats i samband med anbudsinfordran eller offentlig auktion har använts för ändamålen i fråga. Anbudstagaren, eller det godkända företaget, som accepterat att köpa upp alkohol skall informera kommissionen och interventionsorganet om kvantiteten, ändamålet och användningen av de produkter som erhålls genom rektifieringen. Förlusterna får emellertid inte överskrida gränserna enligt b ovan."
Kommissionens förordning (EG) nr 1681/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) För mjölkprodukter beaktas inte innehållet av sackaros när grundbeloppet för bidraget för mjölkhalten är fastställt till noll. Denna bestämmelse bör utvidgas till att gälla även om det inte fastställts något bidrag för mjölkhalten.
(6) Förvaltningskommittén för mjölk och mjölkprodukter har inte yttrat sig inom den tid som dess ordföranden har bestämt.
Förordning (EG) nr 174/1999 ändras på följande sätt:
3. Artikel 16.3 andra stycket skall ersättas med följande: "Innehållet av sackaros skall emellertid inte beaktas om grundbeloppet för den mjölkhalt som avses i punkt 2 andra stycket är fastställt till noll, eller om det inte har fastställts något grundbelopp."
De slutliga licenserna gäller endast för sådan export som avses i punkt 1.
Artikel 9.1 i förordning (EG) nr 1498/1999 skall ersättas med följande: "1. varje arbetsdag före kl. 18.00, utom för kvantiteter för vilka exportlicens begärts, antingen enligt artikel 18 eller artikel 19.5 i förordning (EG) nr 174/1999, eller för leveranser av livsmedelshjälp enligt artikel 10.4 i Uruguayrundans jordbruksavtal, översända uppgifter om följande:
b) De kvantiteter, fördelade efter begäran, efter nummer i exportbidragsnomenklaturen för mjölkprodukter och efter kod för bestämmelseort, för vilka det samma dag begärts sådan tillfällig licens som avses i artikel 8 i förordning (EG) nr 174/1999, med angivande av sista dag för att lämna in anbud samt kvantiteten i anbudsinfordran, eller, om det rör sig om en anbudsinfordran som öppnats av de väpnade styrkorna i enlighet med artikel 36.1 c i kommissionens förordning (EG) nr 800/19991(1) i vilken någon kvantitet inte specificeras, med angivande av den beräknade kvantiteten, fördelad enligt vad som sägs ovan (kod för IDES-meddelande: 2).
Artikel 3
av den 23 oktober 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
av följande skäl:
(3) Särskilt eftersom nya dyra tekniska metoder har införts genom rådets förordning (EG) nr 1593/2000 av den 17 juli 2000 om ändring av förordning (EEG) nr 3508/92 om ett integrerat system för administration och kontroll av vissa stödsystem inom gemenskapen(4), i form av förbättringar av systemet för identifiering av jordbruksskiften med hjälp av GIS-system och digitala ortofotosystem, är ett bidrag från gemenskapen motiverat för att täcka en del av medlemsstaternas kostnader för de nya åtgärdsprogrammen inom detta område. För den juridiska tydlighetens skull bör därför sista strecksatsen i artikel 5 i förordning (EG) nr 723/97 strykas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. I första meningen i artikel 4.1 skall orden "fem år i följd" ersättas med orden "sju år i följd".
om komplettering av bilagan till förordning (EG) nr 2400/96 om upptagandet av vissa namn i Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar som föreskrivs i rådets förordning (EEG) nr 2081/92 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel(1), senast ändrad genom kommissionens förordning (EG) nr 2796/2000(2), särskilt artikel 6.3 och 6.4 i denna, och
(2) Det har i enlighet med artikel 6.1 i nämnda förordning konstaterats att de två ansökningarna är förenliga med den förordningen, särskilt eftersom de omfattar alla komponenter som avses i artikel 4.
(5) Bilagan till denna förordning kompletterar bilagan till kommissionens förordning (EG) nr 2400/96(4), senast ändrad genom förordning (EG) nr 2372/2001(5).
Bilagan till förordning (EG) nr 2400/96 skall kompletteras med de produktnamn som anges i bilagan till denna förordning och dessa namn skall tas upp i Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar såsom skyddad ursprungsbeteckning (SUB) eller skyddad geografisk beteckning (SGU) i enlighet med artikel 6.3 i förordning (EEG) nr 2081/92.
Kommissionens beslut
(2002/79/EG)
med beaktande av rådets direktiv 93/43/EEG av den 14 juni 1993 om livsmedelshygien(1), särskilt artikel 10.1 i detta, och
(2) Vetenskapliga livsmedelskommittén har konstaterat att aflatoxin B1 även i extremt låga doser orsakar levercancer och dessutom är genotoxisk.
(5) Den 8-21 maj 2001 besökte kommissionens kontor för livsmedels- och veterinärfrågor Kina för att bedöma de befintliga kontrollsystemen för att hindra aflatoxinkontaminering av jordnötter avsedda för export till Europeiska gemenskapen. Vid detta besök konstaterades bland annat att kontrollen av aflatoxinhalten i jordnötter var minimal såväl i produktionen som i den allmänna bearbetningen. Brister i laboratoriehanteringen konstaterades också. För att garantera ett fullgott skydd för folkhälsan bör därför särskilda villkor införas för jordnötter och produkter framställda av jordnötter som har sitt ursprung i eller försänds från Kina.
(8) Av resultaten från det ovannämnda besöket framgår att de kinesiska myndigheterna för närvarande inte kan garantera att provresultaten är tillförlitliga eller att certifieringen avser hela sändningen. Det är därför mycket tveksamt hur tillförlitliga intyg är som avser jordnötter med ursprung i Kina.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Jordnötter som omfattas av KN-nummer 1202 10 90 eller 1202 20 00.
2. Sändningar får importeras till gemenskapen endast genom de införselplatser som anges i bilaga II.
5. Medlemsstaterna skall ta prover ur alla sändningar och analysera halterna av aflatoxin B1 och den totala aflatoxinhalten i sändningen innan denna släpps ut på marknaden från införselplatsen, och skall underrätta kommissionen om resultaten.
av den 14 mars 2002
EUROPAPARLAMENTET HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska kol- och stålgemenskapen, särskilt artikel 107 d.4,
med rådets godkännande, och
(2) Genom rådets förordning (EG, EKSG, Euratom) nr 2673/1999 om ändring av budgetförordningen inrättades ett särskilt avsnitt för ombudsmannen i Europeiska unionens allmänna budget och i konsekvens med detta ändrades berörda bestämmelser i budgetförordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
om att bilda Europeiska gruppen av regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
(1) Ett nytt regelverk för nät och tjänster inom området elektronisk kommunikation har inrättats i enlighet med följande direktiv från Europaparlamentet och rådet: 2002/21/EG av den 7 mars 2002 om ett gemensamt regelverk för elektroniska kommunikationsnät och kommunikationstjänster ("ramdirektivet")(1), 2002/19/EG av den 7 mars 2002 om tillträde till och samtrafik mellan elektroniska kommunikationsnät och tillhörande utrustning ("samtrafikdirektivet")(2), 2002/20/EG av den 7 mars 2002 om auktorisation för elektroniska kommunikationsnät och kommunikationstjänster ("tillståndsdirektivet")(3) samt 2002/22/EG av den 7 mars 2002 om samhällsomfattande tjänster och användares rättigheter avseende elektroniska kommunikationsnät och kommunikationstjänster ("direktivet om samhällsomfattande tjänster")(4).
(4) Att bestämmelserna tillämpas på ett enhetligt sätt i alla medlemsstater är av avgörande betydelse för att man skall lyckas med att utveckla en gemensam marknad för nät och tjänster inom området elektronisk kommunikation. I det nya regelverket fastställs mål och ramar för de nationella regleringsmyndigheternas åtgärder, samtidigt som de får handlingsutrymme för att inom bestämda områden väga in nationella särdrag vid tillämpningen av bestämmelserna.
(7) Gruppen bör fungera som ett organ som bistår kommissionen med utredningar, diskussioner och rådgivning inom området elektronisk kommunikation, däribland även i frågor som rör genomförande och revidering av rekommendationer avseende relevanta produkt- och tjänstemarknader samt när det gäller att utforma beslutet om transnationella marknader.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Härmed inrättas en rådgivande grupp som skall bestå av oberoende nationella regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation och vars namn skall vara Europeiska gruppen av regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation (nedan kallad gruppen).
I detta direktiv avses med regleringsmyndighet: myndighet som inrättats i respektive medlemsstat för övervakning av den löpande tolkningen och tillämpningen av bestämmelserna i de direktiv som rör elektroniska kommunikationsnät och elektroniska kommunikationstjänster såsom de är definierade i ramdirektivet.
Gruppen skall vara rådgivare till kommissionen och bistå den när det gäller att befästa den inre marknaden för nät och tjänster inom området elektronisk kommunikation.
Ledamöter
Artikel 5
Gruppen skall inom sig utse en ordförande. Verksamheten får i tillämpliga fall organiseras så att den fördelas på undergrupper och sakkunniggrupper.
Kommissionen skall vara företrädd vid gruppens samtliga möten och ha möjlighet att närvara vid samtliga de möten som undergrupperna och sakkunniggrupperna håller.
Samråd
Sekretess
Årsberättelse
Ikraftträdande
av den 21 november 2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) Uppdateringen av inventeringen av uppgifterna bör ta hänsyn till behovet av människors hälsa inom gemenskapen och till gemenskapslagstiftningens krav inom livsmedelssektorn.
(6) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga livsmedelskommittén.
Bilagan till beslut 94/652/EG ersätts med texten i bilagan till det här beslutet.
Europaparlamentets och rådets direktiv 2002/14/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) Kommissionen har samrått med arbetsmarknadens parter på gemenskapsnivå om den möjliga inriktningen av en gemenskapsåtgärd för information till och samråd med arbetstagare i företag inom gemenskapen.
(6) De rättsliga ramar som finns på nationell nivå och på gemenskapsnivå för att säkerställa arbetstagarnas deltagande i företagets angelägenheter och i de beslut som berör dem har inte alltid kunnat förhindra att ingripande beslut som påverkar arbetstagarna har fattats och offentliggjorts utan att lämpliga förfaranden för information och samråd ägt rum i förväg.
(9) Det är en förutsättning att information ges och samråd äger rum i god tid i förväg om företagens omstrukturering och anpassning till de nya villkor som globaliseringen av ekonomin skapar skall kunna bli framgångsrik, bland annat genom att nya former för arbetets organisation utvecklas.
(12) Inträdet i den tredje etappen av den ekonomiska och monetära unionen har medfört en fördjupad och ökad konkurrens på europeisk nivå. Detta kräver att stödåtgärder vidtas på nationell nivå.
(15) Detta direktiv påverkar inte de nationella system inom vilkas ram det konkreta utövandet av denna rättighet förutsätter en kollektiv viljeyttring från rättsinnehavarnas sida.
(18) Denna allmänna ram har till syfte att fastställa minimiföreskrifter som skall tillämpas i hela gemenskapen men den hindrar inte medlemsstaterna från att anta bestämmelser som är förmånligare för arbetstagarna.
(21) Emellertid bör medlemsstater där det inte finns något lagstadgat system för information till och samråd med arbetstagare eller arbetstagarrepresentanter ha möjlighet att under en övergångsperiod ytterligare begränsa tillämpningsområdet för detta direktiv vad gäller antalet anställda.
(24) Man bör undvika att påverka vissa specifika regler om information till och samråd med arbetstagare i vissa nationella lagstiftningar, vilka gäller företag och driftställen som ägnar sig åt politik, yrkessammanslutningars verksamhet, religiös verksamhet, välgörenhet, utbildning, vetenskap, konst, information eller opinionsbildning.
(27) Information och samråd innebär rättigheter och skyldigheter för arbetsmarknadens parter på företags- eller driftställenivå.
(30) Övriga rättigheter till information och samråd, inklusive de rättigheter som följer av rådets direktiv 94/45/EG av den 22 september 1994 om inrättandet av ett europeiskt företagsråd eller ett förfarande i gemenskapsföretag och grupper av gemenskapsföretag för information till och samråd med arbetstagare(7), bör inte påverkas av detta direktiv.
Artikel 1
2. Formerna för information och samråd skall fastställas och genomföras i enlighet med nationell lagstiftning och den praxis för relationerna mellan arbetsmarknadens parter som finns i de enskilda medlemsstaterna på ett sådant sätt att ändamålet med desamma säkerställs.
Definitioner
b) driftställe: en verksamhetsenhet som definieras enligt nationell lagstiftning och nationell praxis där ekonomisk verksamhet som inbegriper mänskliga och materiella resurser bedrivs kontinuerligt och som är belägen inom en medlemsstats territorium,
e) arbetstagarrepresentanter: företrädare för arbetstagare enligt definitionen i nationell lagstiftning och/eller nationell praxis,
Artikel 3
a) företag som i en medlemsstat sysselsätter minst 50 arbetstagare, eller
2. I enlighet med principerna och målen i detta direktiv får medlemsstaterna fastställa särskilda bestämmelser, som skall tillämpas på företag eller driftställen som direkt och huvudsakligen ägnar sig åt politik, yrkessammanslutningars verksamhet, religiös verksamhet, välgörenhet, utbildning, vetenskap, konst, information eller opinionsbildning, under förutsättning att sådana bestämmelser redan förekommer i nationell lagstiftning vid det datum då detta direktiv träder i kraft.
Former för information och samråd
a) Information om den senaste och den förväntade utvecklingen av företagets eller driftställets verksamhet och ekonomiska situation.
3. Informationen skall överlämnas vid ett sådant tillfälle, på ett sådant sätt och med ett sådant innehåll som gör det möjligt för särskilt arbetstagarrepresentanterna att granska informationen på ett adekvat sätt och vid behov förbereda samråd.
b) på den lednings- och representationsnivå som är relevant med hänsyn till den fråga som behandlas,
e) i syfte att söka nå en överenskommelse när det gäller de beslut som omfattas av arbetsgivarens befogenheter och som avses i punkt 2 c).
Medlemsstaterna får ge arbetsmarknadens parter tillåtelse att på lämplig nivå, inbegripet på företags- eller driftställesnivå, fritt och när som helst genom avtal fastställa formerna för information till och samråd med arbetstagare. Dessa avtal och de avtal som redan finns vid den tidpunkt som anges i artikel 11 samt alla därpå följande förnyelser av sådana avtal får på de villkor och med de begränsningar som fastställs av medlemsstaterna innehålla bestämmelser som avviker från bestämmelserna i artikel 4, om de överensstämmer med principerna i artikel 1.
1. Medlemsstaterna skall på de villkor och med de begränsningar som fastställs i nationell lagstiftning föreskriva att de arbetstagarrepresentanter och experter som eventuellt biträder dem inte har rätt att för arbetstagare eller tredje man röja information som de i företagets eller driftställets legitima intresse uttryckligen fått i förtroende. Denna förpliktelse skall fortsätta att gälla oavsett var experterna eller företrädarna befinner sig, även efter det att deras mandatperiod har löpt ut. En medlemsstat kan emellertid tillåta arbetstagarrepresentanter eller någon som biträder dem att vidarebefordra konfidentiell information till arbetstagare eller tredje man som är bundna av tystnadsplikt.
Artikel 7
Artikel 8
2. Medlemsstaterna skall föreskriva lämpliga påföljder, som skall tillämpas när arbetsgivaren eller arbetstagarrepresentanterna överträder bestämmelserna i detta direktiv. Dessa påföljder skall vara effektiva, proportionella och avskräckande.
1. Detta direktiv skall inte påverka tillämpningen av de särskilda förfaranden för information och samråd som avses i artikel 2 i direktiv 98/59/EG och i artikel 7 i direktiv 2001/23/EG.
4. Genomförandet av detta direktiv skall inte utgöra något tillräckligt skäl för tillbakagång i förhållande till den nuvarande situationen i medlemsstaterna och i förhållande till arbetstagarnas allmänna skyddsnivå på det område som omfattas av direktivet.
Om det i en medlemsstat, vid den tidpunkt då detta direktiv träder i kraft, varken finns något allmänt, varaktigt och lagstadgat system för information till och samråd med arbetstagare eller något allmänt, varaktigt och lagstadgat system för arbetstagarrepresentation på arbetsplatsen, genom vilket de anställda kan företrädas, får denna medlemsstat, trots vad som sägs i artikel 3, såvitt avser detta ändamål begränsa tillämpningen av de nationella genomförandebestämmelserna för direktivet till
Artikel 11
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Senast den 23 mars 2007 skall kommissionen i samråd med medlemsstaterna och arbetsmarknadens parter på gemenskapsnivå se över tillämpningen av detta direktiv och vid behov föreslå nödvändiga ändringar.
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Detta direktiv riktar sig till medlemsstaterna.
om ändring för nittonde gången av rådets direktiv 76/769/EEG om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar) (azofärger)
med beaktande av kommissionens förslag(1),
av följande skäl:
(3) Fullbordandet av den inre marknaden och dess funktion påverkas av att vissa medlemsstater redan har begränsat eller planerat att begränsa användningen av azofärgade textilier och läderartiklar. Det är därför nödvändigt att tillnärma medlemsstaternas lagstiftning på detta område, och bilaga I till rådets direktiv 76/769/EEG av den 27 juli 1976 om tillnärmning av medlemsstaternas lagar och andra författningar om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar)(4) måste därför ändras.
(6) För textilier som framställts av återanvända fibrer bör en maximikoncentration på 70 ppm tillämpas för de aminer som är förtecknade i punkt 43 i tillägget till direktiv 76/769/EEG. Detta bör gälla under en övergångsperiod fram till den 1 januari 2005 om aminerna avges via rester från tidigare färgning av samma fibrer. Detta kommer att möjliggöra återanvändning av textilier, vilket generellt sett är gynnsamt för miljön.
(9) Mot bakgrund av nya vetenskapliga rön bör bestämmelserna om vissa azofärger ses över, särskilt när det gäller behovet av att inbegripa andra material som inte omfattas av detta direktiv och andra aromatiska aminer. Särskild uppmärksamhet bör ägnas eventuella risker för barn.
Artikel 1
Kommissionen skall i enlighet med förfarandet i artikel 2a i direktiv 76/769/EEG anta analysmetoder för tillämpning av punkt 43 i bilaga I till det direktivet.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
om ändring av rådets direktiv 92/6/EEG om montering och användning av hastighetsbegränsande anordningar i vissa kategorier av motorfordon inom gemenskapen
med beaktande av kommissionens förslag(1),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) Användningen av hastighetsbegränsande anordningar för de tyngsta motorfordonskategorierna har haft en gynnsam inverkan på trafiksäkerheten. Den har också bidragit till miljöskyddet.
(5) Tillämpningsområdet för direktiv 92/6/EEG bör utvidgas till att omfatta motorfordon i kategori M2, fordon i kategori M3 med en totalvikt på över 5 ton men högst 10 ton samt till fordon i kategori N2.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artiklarna 1-5 skall ersättas med följande:
Med kategori M2, M3, N2 och N3 avses de kategorier som anges i bilaga II till direktiv 70/156/EEG(6).
Fordon i kategori M3 vars totalvikt överstiger 10 ton och som registrerades före den 1 januari 2005 får även i fortsättningen vara utrustade med anordningar där den högsta hastigheten ställts in på 100 km/h.
2. När det gäller den hastighetsbegränsande anordningen i fordon som är registrerade inom medlemsstaternas territorium och som endast används för transport av farligt gods har medlemsstaterna rätt att kräva att denna är inställd så att dessa fordon inte kan överskrida en högsta hastighet som understiger 90 km/h.
a) fordon som registrerats den 1 januari 1994 eller senare, från och med den 1 januari 1994,
ii) från och med den 1 januari 1996 om det rör sig om fordon som endast används för nationella transporter.
b) fordon som uppfyller de gränsvärden som anges i direktiv 88/77/EEG(7) och registrerats mellan den 1 oktober 2001 och den 1 januari 2005,
3. Varje medlemsstat får bevilja undantag från tillämpningen av artiklarna 2 och 3 under högst tre år från och med den 1 januari 2005 för fordon som tillhör kategori M2 eller som tillhör kategori N2 med en totalvikt på över 3,5 ton men högst 7,5 ton, är registrerade i det nationella fordonsregistret och inte används på en annan medlemsstats territorium.
2. Hastighetsbegränsande anordningar skall monteras av sådana verkstäder eller organ som är godkända av medlemsstaterna.".
Kommissionen skall i samband med åtgärdsprogrammet om trafiksäkerhet för perioden 2002-2010 utvärdera återverkningarna på trafiksäkerheten och vägtrafiken av att de hastighetsbegränsande anordningar som föreskrivs i detta direktiv används i fordon i kategori M2 och fordon i kategori N2 med en totalvikt av högst 7,5 ton.
Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 2005. De skall genast underrätta kommissionen om detta.
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets direktiv 2002/87/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
i enlighet med förfarandet i artikel 251 i fördraget(4), och
(2) Den senaste utvecklingen på finansmarknaderna har lett till skapandet av finansiella grupper som tillhandahåller tjänster och produkter inom olika sektorer av finansmarknaderna - så kallade finansiella konglomerat. Hittills har det inte förekommit någon form av tillsyn på gruppnivå över kreditinstitut, försäkringsföretag och värdepappersföretag som ingår i ett sådant konglomerat, särskilt vad gäller solvensställning och riskkoncentration på konglomeratnivå, transaktioner inom det finansiella konglomeratet, processer för intern riskhantering på konglomeratnivå och ledningens lämplighet. Några av dessa konglomerat är bland de största finansiella grupper som verkar på finansmarknaderna, och de tillhandahåller tjänster i en global omfattning. Om sådana konglomerat, och särskilt kreditinstitut, försäkringsföretag och värdepappersföretag som ingår i ett sådana konglomerat, skulle stöta på finansiella problem kan de allvarligt destabilisera det finansiella systemet och påverka enskilda insättare, försäkringstagare och investerare.
(5) För att den extra tillsynen över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat skall bli effektiv bör den tillämpas på alla sådana konglomerat, vars sektorsöverskridande finansiella verksamhet är betydande, vilket är fallet när vissa trösklar har uppnåtts oavsett hur de är strukturerade. Denna extra tillsyn bör täcka all finansiell verksamhet som anges i den finansiella särlagstiftningen och alla enheter som huvudsakligen ägnar sig åt sådan verksamhet bör omfattas av den extra tillsynen, inklusive kapitalförvaltningsbolagen.
(8) Finansiella konglomerat leds ofta utifrån affärsområden som inte helt motsvarar konglomeratets juridiska strukturer. För att beakta denna tendens bör kraven på ledningen utvidgas ytterligare, särskilt när det gäller ledningen av blandade finansiella holdingföretag.
(11) De berörda behöriga myndigheterna och särskilt samordnaren bör ha de erforderliga medlen för att från enheterna i ett finansiellt konglomerat eller från andra behöriga myndigheter kunna erhålla de upplysningar som krävs för att utöva sin extra tillsyn.
(14) Det kan antas att det finns en likvärdig och lämplig ordning för extra tillsyn endast om tillsynsmyndigheterna i tredje land har samtyckt till att samarbeta med de berörda behöriga myndigheterna om metoderna och målen för att utöva extra tillsyn över reglerade enheter i ett finansiellt konglomerat.
(17) I detta direktiv iakttas de grundläggande rättigheter och principer som erkänns särskilt i Europeiska unionens stadga om grundläggande rättigheter.
(20) De befintliga särreglerna för kreditinstitut, försäkringsföretag och värdepappersföretag bör kompletteras upp till en miniminivå, särskilt för att undvika tillsynsarbitrage mellan särreglerna och reglerna för finansiella konglomerat. Rådets första direktiv 73/239/EEG av den 24 juli 1973 om samordning av lagar och andra författningar angående rätten att etablera och driva verksamhet med annan direkt försäkring än livförsäkring(6), rådets första direktiv 79/267/EEG av den 5 mars 1979 om samordning av lagar och andra författningar om rätten att starta och driva direkt livförsäkringsrörelse(7), rådets direktiv 92/49/EEG av den 18 juni 1992 om samordning av lagar och andra författningar som avser annan direkt försäkring än livförsäkring (tredje direktivet om annan direkt försäkring än livförsäkring)(8), rådets direktiv 92/96/EEG av den 10 november 1992 om samordning av lagar och andra författningar som avser direkt livförsäkring (tredje livförsäkringsdirektivet)(9), rådets direktiv 93/6/EEG av den 15 mars 1993 om kapitalkrav för värdepappersföretag och kreditinstitut(10) och rådets direktiv 93/22/EEG av den 10 maj 1993 om investeringstjänster inom värdepappersområdet(11) samt Europaparlamentets och rådets direktiv 98/78/EG av den 27 oktober 1998 om extra tillsyn över försäkringsföretag som ingår i en försäkringsgrupp(12) och Europaparlamentets och rådets direktiv 2000/12/EG av den 20 mars 2000 om rätten att starta och driva verksamhet i kreditinstitut(13) bör därför ändras på motsvarande sätt. Målet om ytterligare harmonisering kan dock bara uppnås stegvis och måste baseras på en grundlig analys.
KAPITEL I
Mål
Definitioner
2. försäkringsföretag: ett försäkringsföretag i den mening som avses i artikel 6 i direktiv 73/239/EEG, artikel 6 i direktiv 79/267/EEG eller artikel 1 b i direktiv 98/78/EG.
5. kapitalförvaltningsbolag: ett förvaltningsbolag i den mening som avses i artikel 1a.2 i rådets direktiv 85/611/EEG av den 20 december 1985 om samordning av lagar och andra författningar som avser företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag)(14), samt ett företag vars säte är beläget utanför gemenskapen, vilket, om det hade sitt säte i gemenskapen, skulle behöva auktorisation i enlighet med artikel 5.1 i det direktivet.
8. finansiell sektor: en sektor som består av en eller flera av följande enheter:
c) Ett värdepappersföretag eller ett finansiellt institut enligt artikel 2.7 i direktiv 93/6/EEG (sektorn för investeringstjänster).
10. dotterföretag: ett dotterföretag i den mening som avses i artikel 1 i direktiv 83/349/EEG och varje företag över vilket ett moderföretag enligt de behöriga myndigheterna i praktiken utövar ett bestämmande inflytande. Alla dotterföretag till dotterföretag skall också betraktas som dotterföretag till det moderföretag som är överordnat dessa företag.
13. nära förbindelser: en situation där två eller flera fysiska eller juridiska personer är förenade genom
Som nära förbindelse skall även anses en situation där två eller flera fysiska eller juridiska personer kontrolleras genom en varaktig förbindelse till en och samma person.
b) Om en reglerad enhet i den mening som avses i artikel 1 finns i toppen av gruppen, är den antingen ett moderföretag till en enhet i den finansiella sektorn, en enhet med ägarintresse i en enhet i den finansiella sektorn eller en enhet som har ett sådant samband med en enhet i den finansiella sektorn som avses i artikel 12.1 i direktiv 83/349/EEG.
e) Den konsoliderade och/eller aggregerade verksamheten i gruppens enheter inom försäkringssektorn och den konsoliderade och/eller aggregerade verksamheten i gruppens enheter inom bank- och värdepapperssektorn är betydande enligt artikel 3.2 eller 3.3.
16. behöriga myndigheter: de nationella myndigheter i medlemsstaterna som enligt lag eller annan författning har behörighet att utöva tillsyn över kreditinstitut, försäkringsföretag och/eller värdepappersföretag såväl enskilt som på gruppnivå.
b) samordnaren som utsetts i enlighet med artikel 10, om annan än de myndigheter som anges under a,
19. riskkoncentration: alla exponeringar med förlustpotential som bärs av enheter inom ett finansiellt konglomerat, vilka är tillräckligt stora för att hota dessa reglerade enheters solvens eller deras finansiella ställning i allmänhet; sådana exponeringar kan orsakas av motpartsrisk/kreditrisk, investeringsrisk, försäkringsrisk, marknadsrisk eller andra risker, eller en kombination av eller samverkan mellan dessa risker.
1. För att en grupp skall bedömas bedriva verksamhet huvudsakligen inom den finansiella sektorn i den mening som avses i artikel 2.14 c, skall balansomslutningen inom gruppens reglerade och icke reglerade enheter inom den finansiella sektorn utgöra mer än 40 % av hela gruppens balansomslutning.
3. Sektorsövergripande verksamhet skall också bedömas som betydande i den mening som avses i artikel 2.14 e, om balansomslutningen för den minsta finansiella sektorn i gruppen överstiger 6 miljarder euro. Om gruppen inte uppnår det tröskelvärde som anges i punkt 2, får de relevanta behöriga myndigheterna i samförstånd besluta sig för att inte betrakta gruppen som ett finansiellt konglomerat eller att inte tillämpa bestämmelserna i artiklarna 7, 8 eller 9, om de anser att det inte är nödvändigt eller att det vore olämpligt eller vilseledande att låta gruppen omfattas av detta direktivs räckvidd eller att tillämpa sådana bestämmelser med hänsyn till de mål som skall uppnås genom extra tillsyn, till exempel med beaktande av följande:
Beslut som fattas i överensstämmelse med denna punkt skall anmälas till övriga berörda behöriga myndigheter.
b) beakta att de trösklar som anges i punkterna 1 och 2 har iakttagits under tre år i följd, så att plötsliga byten av det tillämpliga regelverket kan undvikas, och bortse ifrån att så har skett, om väsentliga förändringar i gruppens struktur uppstår.
6. Om de procentsatser som avses i punkterna 1 och 2 hamnar under 40 % respektive 10 % för konglomerat som redan är föremål för extra tillsyn, skall vid tillämpningen av dessa punkter en lägre procentsats på 35 % respektive 8 % tillämpas under de tre följande åren, för att plötsliga byten av tillämpligt regelverk skall undvikas.
7. De beräkningar som anges i denna artikel och som rör balansräkningen skall utföras på grundval av den aggregerade balansomslutningen för gruppens enheter enligt deras årsbokslut. Vid denna beräkning skall företag som är föremål för ett ägarintresse ingå till det belopp i deras balansomslutning som motsvarar den aggregerade proportionella andel som gruppen innehar. Om sammanställd redovisning emellertid finns tillgänglig, skall denna användas i stället för aggregerad redovisning.
Identifiering av ett finansiellt konglomerat
- skall de behöriga myndigheter som har auktoriserat reglerade enheter i denna grupp, om så är nödvändigt, ha ett nära samarbete,
KAPITEL II
RÄCKVIDD
1. Utan att det påverkar särreglernas bestämmelser om tillsyn skall medlemsstaterna ombesörja extra tillsyn över de reglerade enheter som avses i artikel 1, i den omfattning och på det sätt som föreskrivs i detta direktiv.
b) Varje reglerad enhet vars moderföretag är ett blandat finansiellt holdingföretag med huvudkontor inom gemenskapen.
3. Varje reglerad enhet som inte är föremål för extra tillsyn enligt punkt 2 och vars moderföretag är en reglerad enhet eller ett blandat finansiellt holdingföretag med huvudkontor utanför gemenskapen skall vara föremål för extra tillsyn på nivån finansiellt konglomerat i den omfattning och på det sätt som föreskrivs i artikel 18.
Vid tillämpning av det första stycket på "kooperativa grupper" skall de behöriga myndigheterna beakta de offentliga finansieringsåtaganden som dessa grupper har gentemot andra finansiella enheter.
FINANSIELL STÄLLNING
1. Utan att särreglerna åsidosätts skall extra tillsyn över kapitaltäckningen i de reglerade enheterna i ett finansiellt konglomerat utövas enligt de regler som anges i punkterna 2-5, i artikel 9, i avsnitt 3 i detta kapitel och i bilaga I.
De krav som avses i första och andra stycket skall vara föremål för samordnarens tillsyn enligt avsnitt 3.
3. För den beräkning av kapitaltäckningskraven som avses i punkt 2 första stycket skall följande enheter omfattas av extra tillsyn i den form och utsträckning som fastställs i bilaga I:
c) Värdepappersföretag eller finansiella institut i den mening som avses i artikel 2.7 i direktiv 93/6/EEG.
Vid tillämpning av metod 2 eller 3 (Avräknings- och totalmetoden respektive Metod för kravavräkning eller avräkning av bokfört värde) vilka avses i bilaga I skall hänsyn tas till den proportionella andel som moderföretaget eller företaget med ägarintresse innehar i en annan enhet i gruppen. Med "proportionell andel" avses den del av det tecknade kapitalet som direkt eller indirekt innehas av detta företag.
b) Om enheten är av försumbar betydelse i förhållande till målen för den extra tillsynen över reglerade enheter i ett finansiellt konglomerat.
I det fall som nämns i c i första stycket skall samordnaren, utom i brådskande fall, samråda med de andra relevanta behöriga myndigheterna innan beslut fattas.
Riskkoncentration
Samordnaren skall övervaka dessa riskkoncentrationer i enlighet med avsnitt 3.
Artikel 8
2. Medlemsstaterna skall kräva att reglerade enheter eller blandade finansiella holdingföretag regelbundet och minst en gång per år till samordnaren rapporterar samtliga transaktioner inom det finansiella konglomeratet enligt reglerna i denna artikel och i bilaga II. I den mån de tröskelvärden som anges i sista meningen i första stycket i bilaga II inte har fastställts, skall en transaktion inom det finansiella konglomeratet åtminstone anses som betydande, om beloppet överstiger 5 % av det totala belopp som kapitaltäckningskraven uppgår till på nivån finansiellt konglomerat.
3. Till dess att gemenskapens lagstiftning har samordnats ytterligare får medlemsstaterna fastställa kvantitativa gränser och kvalitativa krav eller tillåta sina behöriga myndigheter att fastställa kvantitativa gränser och kvalitativa krav eller vidta andra tillsynsåtgärder som skulle kunna uppfylla målen för extra tillsyn när det gäller transaktioner inom det finansiella konglomeratet av reglerade enheter i ett finansiellt konglomerat.
Rutiner för intern kontroll och metoder för riskhantering
a) Ett sunt styre och en sund förvaltning, varvid lämpliga ledande organ på nivån finansiellt konglomerat skall godkänna och regelbundet övervaka strategier och inriktningar med beaktande av alla risker de tar.
3. Rutinerna för intern kontroll skall innehålla följande:
4. Medlemsstaterna skall se till att det i alla företag som omfattas av extra tillsyn enligt artikel 5 finns erforderliga rutiner för intern kontroll för att ta fram de uppgifter och upplysningar som kan vara av betydelse för den extra tillsynen.
ÅTGÄRDER FÖR ATT UNDERLÄTTA EXTRA TILLSYN
1. För att säkerställa korrekt extra tillsyn över de reglerade enheterna i ett finansiellt konglomerat skall en enda samordnare med ansvar för samordning och utövande av den extra tillsynen utses bland de berörda medlemsstaternas behöriga myndigheter, inbegripet dem som finns i den medlemsstat i vilken det blandade finansiella holdingföretaget har sitt huvudkontor.
b) Om ett finansiellt konglomerat inte leds av en reglerad enhet, skall den behöriga myndighet som identifieras enligt följande principer fungera som samordnare:
Om två eller flera reglerade enheter som verkar inom olika finansiella sektorer har auktoriserats i den medlemsstat där det blandade finansiella holdingföretaget har sitt huvudkontor, skall samordningen utövas av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som verkar inom den största finansiella sektorn.
iv) Om det finansiella konglomeratet utgör en grupp utan något moderföretag i toppen, eller i övriga fall, skall samordningen utövas av den behöriga myndighet som har auktoriserat den reglerade enhet som har den största balansomslutningen inom den största finansiella sektorn.
Samordnarens uppgifter
b) Övervakning av och bedömning av ett finansiellt konglomerats finansiella ställning.
e) Planering och samordning av tillsynen, såväl löpande som i krissituationer, i samarbete med de berörda behöriga myndigheterna.
2. Samordnaren bör, när den behöver uppgifter som redan överlämnats till en annan behörig myndighet i enlighet med särreglerna, vända sig till denna myndighet närhelst detta är möjligt i syfte att undvika dubblering av rapporteringen till de olika myndigheter som utövar tillsyn.
Samarbete och utbyte av uppgifter mellan behöriga myndigheter
a) Identifiering av hur alla större enheter som tillhör det finansiella konglomeratet är grupperade och av de behöriga myndigheter som ansvarar för tillsynen över de reglerade enheterna i gruppen.
d) Det finansiella konglomeratets största aktieägare och ledning.
g) Negativ utveckling i reglerade enheter eller i andra enheter i det finansiella konglomeratet som skulle kunna påverka de reglerade enheterna allvarligt.
2. Utan att det påverkar dessa myndigheters respektive ansvar enligt särreglerna skall de berörda behöriga myndigheterna innan de fattar beslut samråda med varandra i följande fall, om deras beslut är av betydelse för andra behöriga myndigheters tillsynsuppgifter:
En behörig myndighet får besluta att inte samråda i brådskande situationer eller när ett sådant samråd kan äventyra effektiviteten i besluten. Den behöriga myndigheten skall i detta fall utan dröjsmål informera de andra behöriga myndigheterna.
4. Medlemsstaterna skall godkänna att deras behöriga myndigheter utbyter de uppgifter som avses i punkterna 1, 2 och 3 med varandra och med andra myndigheter. Insamling eller innehav av uppgifter om en enhet inom ett finansiellt konglomerat vilken inte är en reglerad enhet skall inte på något sätt anses innebära att de behöriga myndigheterna är skyldiga att utöva någon tillsynsfunktion i förhållande till den enskilda enheten.
Ledningsorgan för blandade finansiella holdingföretag
Tillgång till uppgifter
Artikel 15
De myndigheter som får en sådan begäran skall inom ramen för sin behörighet tillgodose begäran, antingen genom att själva utföra kontrollen, genom att låta en revisor eller expert utföra den eller genom att låta den begärande myndigheten själv utföra den.
Verkställande åtgärder
- av de behöriga myndigheterna när det gäller reglerade enheter. I detta syfte skall samordnaren underrätta de behöriga myndigheterna om sina upptäckter.
Artikel 17
2. Utan att det påverkar tillämpningen av nationella straffrättsliga bestämmelser skall medlemsstaterna se till att påföljder eller åtgärder, vars syfte är att konstaterade överträdelser eller orsakerna till desamma skall upphöra, kan utdömas respektive vidtas gentemot blandade finansiella holdingföretag eller deras faktiska ledare, när dessa bryter mot lagar och andra författningar som antagits för att genomföra bestämmelserna i detta direktiv. I vissa fall kan sådana åtgärder kräva domstols medverkan. De behöriga myndigheterna skall ha ett nära samarbete för att se till att dessa påföljder och åtgärder får avsedd effekt.
Artikel 18
2. I brist på sådan likvärdig tillsyn som avses i punkt 1 skall de behöriga myndigheterna på dessa reglerade myndigheter analogt tillämpa de bestämmelser om extra tillsyn över reglerade enheter som avses i artikel 5.2. Alternativt får de behöriga myndigheterna tillämpa en av de metoder som anges i punkt 3.
Samarbete med behöriga myndigheter i tredje land
KAPITEL III
Kommissionens befogenheter
b) En mer precis formulering av definitionerna i artikel 2 i syfte att säkerställa en enhetlig tillämpning av detta direktiv i gemenskapen.
e) Samordning av bestämmelserna enligt artiklarna 7 och 8 och bilaga II, så att enhetlig tillämpning inom gemenskapen uppmuntras.
Kommitté
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
5. Kommittén får ge allmän vägledning om huruvida det är sannolikt att de system för extra tillsyn som tillämpas av behöriga myndigheter i tredje land kommer att uppfylla det mål för den extra tillsynen som ställs upp i detta direktiv, när det gäller reglerade enheter i ett finansiellt konglomerat vars ledande enhet har sitt huvudkontor utanför gemenskapen. Kommittén skall fortlöpande se över all sådan vägledning och beakta varje förändring i den extra tillsyn som utförs av sådana behöriga myndigheter.
ÄNDRINGAR AV NUVARANDE DIREKTIV
Direktiv 73/239/EEG ändras på följande sätt:
1. Samråd med behöriga myndigheter i den andra berörda medlemsstaten skall genomföras innan auktorisation beviljas för ett försäkringsföretag som
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett försäkringsföretag som är auktoriserat i en annan medlemsstat.
b) är dotterföretag till moderföretaget till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen, eller
2. I artikel 16.2 skall följande stycken läggas till:
- försäkringsföretag i den mening som avses i artikel 6 i detta direktiv, artikel 6 i första direktivet 79/267/EEG av den 5 mars 1979 om samordning av lagar och andra författningar om rätten att starta och driva direkt livförsäkringsrörelse(17) eller artikel 1 b i Europaparlamentets och rådets direktiv 98/78/EG(18),
- kreditinstitut och finansiella institut i den mening som avses i artiklarna 1.1 och 1.5 i Europaparlamentets och rådets direktiv 2000/12/EG(19),
- De instrument som avses i punkt 3.
Om aktier i ett annat kreditinstitut, värdepappersföretag, finansiellt institut, försäkringsföretag, återförsäkringsföretag eller försäkringsholdingbolag innehas tillfälligt i syfte att ge finansiellt bistånd för att rekonstruera och rädda denna enhet, får den behöriga myndigheten bevilja undantag från bestämmelserna om avdrag enligt a och b i fjärde stycket.
Med det avdrag av ägarintresse som anges i detta stycke menas här ägarintresse i den mening som avses i artikel 1 f i direktiv 98/78/EG.".
Direktiv 79/267/EEG ändras på följande sätt:
1. Samråd med behöriga myndigheter i den andra berörda medlemsstaten skall genomföras innan auktorisation beviljas för ett livförsäkringsföretag som
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett försäkringsföretag som är auktoriserat i en annan medlemsstat.
b) är dotterföretag till moderföretaget till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen, eller
2. I artikel 18.2 skall följande stycken läggas till:
- försäkringsföretag i den mening som avses i artikel 6 i detta direktiv, artikel 6 i direktiv 73/239/EEG(23)eller artikel 1 b i Europaparlamentets och rådets direktiv 98/78/EG(24),
- kreditinstitut och finansiella institut i den mening som avses i artiklarna 1.1 och 1.5 i Europaparlamentets och rådets direktiv 2000/12/EG(25),
- De instrument som avses i punkt 3.
För beräkningen av solvensmarginalen enligt detta direktiv får medlemsstaterna föreskriva att försäkringsföretag som är föremål för extra tillsyn enligt direktiv 98/78/EG eller enligt direktiv 2002/87/EG inte behöver dra ifrån poster enligt a och b i tredje stycket i de kreditinstitut, värdepappersföretag, finansiella institut, försäkrings- eller återförsäkringsföretag eller försäkringsholdingbolag som ingår i den extra tillsynen.
Ändring av direktiv 92/49/EEG
"1a. Om köparen av det innehav som avses i punkt 1 är ett försäkringsföretag, ett kreditinstitut eller ett värdepappersföretag med auktorisation i en annan medlemsstat eller moderföretag till en sådan enhet, eller en fysisk eller juridisk person som har ägarkontroll över en sådan enhet, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av ett sådant samråd som avses i artikel 12a i direktiv 73/239/EEG.".
- till centralbanker och andra organ med liknande funktion i egenskap av monetära myndigheter,
Artikel 25
1. I artikel 14 skall följande punkt införas:
"5c. Denna artikel skall inte hindra en behörig myndighet från att
överföra uppgifter för att dessa skall kunna utföra sina uppgifter, och den skall inte heller hindra sådana myndigheter eller organ från att vidarebefordra sådana uppgifter som de kan behöva enligt punkt 4. Uppgifter som erhålls i detta sammanhang skall omfattas av de bestämmelser om tystnadsplikt som fastställs i denna artikel.".
I artikel 7.3 i direktiv 93/6/EEG skall första och andra strecksatsen ersättas med följande text:
Artikel 27
1. I artikel 6 skall följande stycken läggas till:
b) är dotterföretag till moderföretaget till ett kreditinstitut eller försäkringsföretag som är auktoriserat i gemenskapen, eller
2. Artikel 9.2 skall ersättas med följande:
Ändringar i direktiv 98/78/EG
"g) företag med ägarintresse: ett företag som är antingen moderföretag eller ett annat företag som har ett ägarintresse eller ett företag som är knutet till ett annat företag genom ett sådant förhållande som avses i artikel 12.1 i direktiv 83/349/EEG.
j) försäkringsholdingföretag med blandad verksamhet: ett annat moderföretag än ett försäkringsföretag, ett försäkringsföretag i tredje land, ett återförsäkringsföretag, ett försäkringsholdingföretag eller ett blandat finansiellt holdingföretag i den mening som avses i direktiv 2002/87/EG, vilket har minst ett försäkringsföretag bland sina dotterföretag.".
3. I artikel 8.2 skall det första stycket ersättas med följande:
"Artikel 10a
a) försäkringsföretag bland vars delägare det finns företag i den mening som avses i artikel 2 med huvudkontor i tredje land, och
a) att de behöriga myndigheterna i medlemsstaterna kan få fram den information som krävs för att utöva extra tillsyn över försäkringsföretag med huvudkontor inom gemenskapen och med dotterföretag eller ägarintressen i företag utanför gemenskapen, och
Artikel 10b
5. I punkt 1 B i bilaga I skall följande stycke läggas till:
"2.4a Berörda kreditinstitut, värdepappersföretag och finansiella institut
Ändringar av direktiv 2000/12/EG
a) Punkt 9 skall ersättas med följande:
"21. finansiellt holdingföretag: ett finansiellt institut vars dotterföretag uteslutande eller huvudsakligen är kreditinstitut eller finansiella institut, varvid minst ett av dotterföretagen skall vara ett kreditinstitut, och som inte är ett blandat finansiellt holdingföretag i den mening som avses i Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(31).
"Samråd med den behöriga myndighet som har ansvar för tillsynen över försäkringsföretag eller värdepappersföretag skall genomföras innan auktorisation beviljas för ett kreditinstitut som
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett försäkringsföretag som är auktoriserat i gemenskapen.
"2. Om förvärvaren av det innehav som avses i punkt 1 är ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag med auktorisation i en annan medlemsstat eller moderföretag till ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag med auktorisation i en annan medlemsstat, eller en fysisk eller juridisk person som har ägarkontroll över ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag med auktorisation i en annan medlemsstat, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av sådant samråd som avses i artikel 12.".
"12. Sådana ägarposter i andra kreditinstitut och finansiella institut som motsvarar mer än 10 % av deras kapital.
15. Ägarintresse av det slag som avses i artikel 1.9, vilket ett kreditinstitut innehar i
- försäkringsholdingföretag i den mening som avses i artikel 1 led i i direktiv 98/78/EG.
- de instrument som avses i artikel 18.3 i direktiv 79/267/EEG.".
Som ett alternativ till avdrag av poster enligt punkterna 15 och 16 får medlemsstaterna tillåta att deras kreditinstitut också tillämpar metoderna 1, 2 eller 3 i bilaga I i direktiv 2002/87/EG. Metod 1 (metod baserad på sammanställd redovisning) skall endast tillämpas om den behöriga myndigheten är säker på graden av samordnad förvaltning och intern kontroll avseende de enheter som skall inbegripas i tillämpningsområdet för sammanställningen. Den valda metoden skall tillämpas konsekvent över tiden.
5. Artikel 51.3 skall ersättas med följande:
"Utan att det påverkar tillämpningen av artikel 54a skall sammanställningen inte på något sätt anses innebära att de behöriga myndigheterna har skyldighet att utöva tillsyn i förhållande till det enskilda finansiella holdingföretaget.".
"Om företagen står i ett sådant samband som avses i artikel 12.1 i direktiv 83/349/EEG skall de behöriga myndigheterna bestämma hur sammanställningen skall ske.".
"Artikel 54a
9. Följande artikel skall läggas till:
Utan att detta påverkar bestämmelserna i avdelning V kapitel 2 avsnitt 3 i detta direktiv skall medlemsstaterna, då moderföretaget till ett eller flera kreditinstitut är ett holdingföretag med blandad verksamhet, se till att de behöriga myndigheter som ansvarar för tillsynen över dessa kreditinstitut utövar allmän tillsyn över transaktioner mellan kreditinstitutet och holdingföretaget med blandad verksamhet samt dess dotterföretag.
10. I artikel 56.7 skall följande mening läggas till:
"Artikel 56a
Den rådgivande bankrörelsekommittén får ge allmän vägledning om huruvida det är sannolikt att de system för gruppbaserad tillsyn som tillämpas av behöriga myndigheter i tredje land kommer att uppfylla de mål för den gruppbaserade tillsynen som ställs upp i detta kapitel, när det gäller kreditinstitut vars moderföretag har sitt huvudkontor utanför gemenskapen. Kommittén skall fortsätta att se över all sådan vägledning och beakta varje förändring i de system för den gruppbaserade tillsynen som tillämpas av sådana behöriga myndigheter.
KAPITALFÖRVALTNINGSBOLAG
Till dess att särreglerna har samordnats ytterligare skall medlemsstaterna föreskriva att kapitalförvaltningsbolag skall omfattas av
För tillämpningen av det första stycket skall medlemsstaterna föreskriva eller ge sina behöriga myndigheter behörighet att besluta om enligt vilka särregler (för banksektorn, försäkringssektorn eller värdepapperssektorn) kapitalförvaltningsbolag skall omfattas av den gruppbaserade tillsyn och/eller den extra tillsyn som avses i första stycket a. I denna bestämmelse skall särreglerna om i vilken form och utsträckning finansiella institut (om kapitalförvaltningsbolag omfattas av tillämpningsområdet för gruppbaserad tillsyn över kreditinstitut och värdepappersföretag) och återförsäkringsföretag (om kapitalförvaltningsbolag omfattas av tillämpningsområdet för extra tillsyn över försäkringsföretag) skall omfattas också tillämpas på kapitalförvaltningsbolag. Vad avser den extra tillsyn som avses i första stycket b skall kapitalförvaltningsbolaget behandlas som en del av den sektor som det skall räknas till i enlighet med första stycket a.
ÖVERGÅNGS- OCH SLUTBESTÄMMELSER
1. Senast 11 augusti 2007 skall kommissionen till den kommitté för finansiella konglomerat som avses i artikel 21 överlämna en rapport om medlemsstaternas praxis och i förekommande fall om behovet av ytterligare harmonisering i fråga om
- hur betydande transaktioner inom det finansiella konglomeratet och betydande riskkoncentration bör definieras samt om tillsynen över transaktioner inom det finansiella konglomeratet och riskkoncentration som avses i bilaga II, särskilt i fråga om införandet av kvantitativa gränser och kvalitativa krav i detta syfte,
2. Inom ett år efter det att en överenskommelse träffats på internationell nivå om bestämmelserna om eliminering av dubbelt utnyttjande av poster i kapitalbasen i finansiella grupper skall kommissionen undersöka hur bestämmelserna i detta direktiv kan anpassas till dessa internationella överenskommelser och vid behov lägga fram lämpliga förslag.
När medlemsstaterna antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare bestämmelser om hur denna hänvisning skall göras skall varje medlemsstat själv utfärda.
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska unionens officiella tidning.
Detta direktiv riktar sig till medlemsstaterna.
om ändring av bilagorna till rådets direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG beträffande fastställande av gränsvärden för bekämpningsmedelsrester (2,4-D, triasulfuron och tifensulfuronmetyl) i och på spannmål, livsmedel av animaliskt ursprung och vissa produkter av vegetabiliskt ursprung, inklusive frukt och grönsaker
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/642/EEG av den 27 november 1990 om fastställande av gränsvärden för bekämpningsmedelsrester i och på produkter av vegetabiliskt ursprung inklusive frukt och grönsaker(4), senast ändrat genom direktiv 2002/79/EG, särskilt artikel 7 i detta,
(1) Genom kommissionens direktiv 2001/103/EG(7), 2000/66/EG(8) respektive 2001/99/EG(9) infördes de befintliga verksamma ämnena 2,4-D, triasulfuron och tifensulfuronmetyl i bilaga I till direktiv 91/414/EEG för att användas som herbicider, utan att det angavs några särskilda förhållanden som skulle kunna inverka på grödor som eventuellt behandlades med växtskyddsmedel innehållande dessa verksamma ämnen.
(4) I samband med införandet av de berörda verksamma ämnena i bilaga I till direktiv 91/414/EEG avslutades de tekniska och vetenskapliga utvärderingarna genom kommissionens granskningsrapport. Rapporten avslutades den 2 oktober 2001 för 2,4-D, den 13 juli 2000 för triasulfuron och den 29 juni 2001 för tifensulfuronmetyl. I rapporterna fastställs det acceptabla dagliga intaget (ADI) för 2,4-D till 0,05 mg per kg kroppsvikt och dag, för triasulfuron till 0,01 mg per kg kroppsvikt och dag och för tifensulfuronmetyl till 0,01 mg per kg kroppsvikt och dag. Konsumenternas livstidsexponering genom livsmedel som behandlats med de berörda verksamma ämnena har uppskattats och utvärderats med hjälp av de metoder som används inom gemenskapen. Hänsyn har också tagits till de riktlinjer som offentliggjorts av Världshälsoorganisationen(10) samt yttrandet om de använda metoderna från den Vetenskapliga kommittén för växter(11). Det har fastslagits att de föreslagna gränsvärdena inte leder till att de acceptabla dagliga intagen överskrids. Under de utvärderingar och diskussioner som föregick införandet av de berörda verksamma ämnena i bilaga I till direktiv 91/414/EEG noterades inga akuta toxiska effekter som skulle kräva att det fastställs en akut referensdos.
(7) Bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
">Plats för tabell>"
">Plats för tabell>"
Artikel 4
När en medlemsstat antar dessa bestämmelser, skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 6
av den 19 december 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I förordning (EEG) nr 3696/93 fastställs en statistisk indelning av produkter efter näringsgren, nedan kallad CPA, för att tillgodose behovet av statistik inom gemenskapen.
(4) Det är nödvändigt att ändra CPA, behålla det internationellt integrerade systemet och skapa konvergens globalt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 20 februari 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Genom förordning (EG) nr 2529/2001 införs ett nytt bidragssystem som ersätter det system som infördes genom rådets förordning (EG) nr 2467/98 av den 3 november 1998 om den gemensamma organisationen av marknaden för får- och getkött(2), ändrad genom förordning (EG) nr 1669/2000(3). För att ta hänsyn till de nya förfarandena och av tydlighetsskäl är det nödvändigt att införa nya regler som ersätter reglerna i kommissionens förordning (EEG) nr 1481/86 av den 15 maj 1986 om fastställande av priser på färska eller kylda slaktkroppar av lamm på gemenskapens representativa marknader och om registrering av priserna på vissa andra slaktkroppskvaliteter för får inom gemenskapen(4), senast ändrad genom förordning (EG) nr 2877/2000(5).
(4) Det pris som noterats på marknaden skall grunda sig på priser på slaktkroppar exklusive mervärdeskatt men utan avdrag för andra pålagor. Marknadspriset skall noteras med avseende på "slaktkroppsvikten" enligt definitionen i kommissionens beslut 94/434/EG av den 30 maj 1994 om tillämpningsföreskrifter för rådets direktiv 93/25/EEG vad avser statistiska undersökningar av får- och getbestånd och får- och getproduktion(6), senast ändrad genom beslut 1999/47/EG(7). En avvikelse från denna definition bör dock tillåtas för slaktkroppar av unga lamm som väger mellan 9 och 16 kg av hänsyn till marknadspraxis som ger ett högre handelsvärde åt hela slaktkroppar med huvud och slaktbiprodukter.
(7) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för får och getter.
1. Medlemsstater vars fårköttproduktion överstiger 200 ton per år skall senast varje torsdag meddela kommission priserna på färska eller kylda slaktkroppar av lamm och tackor.
1. Marknadspriserna skall noteras med avseende på "slaktvikt" enligt definitionen i beslut 94/434/EG.
När priserna noteras på grundval av priserna för levande djur skall priset per kg levande vikt divideras med en omräkningskoefficient på högst 0,5. Om det är allmän praxis att sälja slaktkroppen med huvud och slaktbiprodukter kan medlemsstaten fastställa en högre koefficient för lamm med en levande vikt upp till 28 kg.
1. När det förekommer marknader mer än en gång under den period på sju dagar som anges i artikel 2.1 skall priset på varje kategori vara det aritmetiska genomsnittet av de priser som har noterats vid varje marknadstillfälle.
Artikel 4
b) Kategorierna av slaktkroppar av lamm.
Artikel 5
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om komplettering av bilagan till förordning (EG) nr 2400/96 om upptagandet av vissa namn i "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar" som föreskrivs i rådets förordning (EEG) nr 2081/92 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel(1), senast ändrad genom kommissionens förordning (EG) nr 2796/2000(2), särskilt artikel 6.3 och 6.4 i denna, och
(2) Det har i enlighet med artikel 6.1 i nämnda förordning konstaterats att ansökan är förenlig med den förordningen, särskilt eftersom den omfattar alla komponenter som avses i artikel 4.
(5) Bilagan till denna förordning kompletterar bilagan till kommissionens förordning (EG) nr 2400/96(4) senast ändrad genom förordning (EG) nr 245/2002(5).
Bilagan till förordning (EG) nr 2400/96 skall kompletteras med det produktnamn som anges i bilagan till denna förordning och detta namn skall tas upp i "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar" såsom skyddad geografisk beteckning (SGB) i enlighet med artikel 6.3 i förordning (EEG) nr 2081/92.
Kommissionens förordning (EG) nr 780/2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Förordning (EG) nr 3063/93 bör därför ändras.
2. I artikel 2.2 skall den första meningen ersättas med följande: "Sammanslutningarna av biodlare skall förelägga den behöriga myndigheten sina program för godkännande.".
b) I punkt 2 skall första strecksatsen ersättas med följande: "- Sammanslutningarnas eller biodlarens namn och adress,".
a) I första stycket skall första och andra strecksatserna ersättas med följande: "- Antal sammanslutningar av biodlare och antal enskilda biodlare som inkommit med stödansökningar.
6. I artikel 6.2 första stycket skall andra meningen utgå.
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om inrättande av en europeisk sjösäkerhetsbyrå
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2 i detta,
med beaktande av Regionkommitténs yttrande(3),
(1) Ett stort antal lagstiftningsåtgärder har antagits inom gemenskapen för att förbättra säkerheten och förhindra förorening i samband med sjötransporter. För att vara effektiv måste sådan lagstiftning tillämpas korrekt och enhetligt i hela gemenskapen. På så sätt säkerställs likvärdiga konkurrens- och marknadsvillkor, minskas den snedvridning av konkurrensen som följer av de ekonomiska fördelar som fartyg som inte uppfyller normerna åtnjuter och gynnas de rederier och andra som bedriver sjöfartsverksamhet på ett seriöst sätt.
(4) För att målsättningarna med byråns inrättande skall uppnås bör byrån utföra ett antal andra viktiga arbetsuppgifter avsedda att höja sjösäkerheten och förhindra förorening från fartyg i de vatten som tillhör medlemsstaterna. I detta avseende bör byrån i samarbete med medlemsstaterna anordna lämplig utbildningsverksamhet beträffande frågor som gäller hamnstatskontroll och flaggstat och tillhandahålla tekniskt stöd i samband med genomförandet av gemenskapslagstiftningen. Den bör underlätta samarbete mellan medlemsstaterna och kommissionen enligt Europaparlamentets och rådets direktiv 2002/59/EG av den 27 juni 2002 om inrättandet av ett övervaknings- och informationssystem för sjötrafik i gemenskapen och om upphävande av rådets direktiv 93/75/EEG(5) genom att utveckla och sköta det informationssystem som behövs dels för att uppnå de mål som uppställs i direktivet, dels i verksamhet som gäller utredningar av allvarliga olyckor till sjöss. Den bör ge kommissionen och medlemsstaterna objektiva, tillförlitliga och jämförbara uppgifter och data om sjösäkerhet och förhindrande av förorening från fartyg, så att dessa kan vidta nödvändiga åtgärder för att förbättra befintliga åtgärder och utvärdera åtgärdernas effektivitet. Den bör se till att den kunskap om sjösäkerhet som finns inom gemenskapen står till förfogande för de stater som ansöker om anslutning. Dessa stater och andra tredjeländer som ingått avtal med Europeiska gemenskapen, genom vilka de antar och genomför gemenskapslagstiftningen inom området för sjösäkerhet och förhindrande av förorening från fartyg, bör ha möjlighet att delta i byråns verksamhet.
(7) Byrån bör tillämpa den relevanta gemenskapslagstiftningen rörande allmänhetens tillgång till handlingar och skydd för enskilda vid databehandling av personuppgifter. Den bör ge allmänheten och alla berörda parter objektiv, tillförlitlig och lättbegriplig information om sin verksamhet.
(10) För att byrån skall fungera väl måste den verkställande direktören vara utsedd på grundval av meriter och dokumenterad skicklighet i förvaltning och ledarskap samt kompetens och erfarenheter som är relevanta för sjösäkerhet och förhindrande av förorening från fartyg och han/hon måste vid utförandet av sina arbetsuppgifter vara helt oavhängig och flexibel när det gäller byråns inre organisation. Den verkställande direktören bör därför förbereda och vidta alla åtgärder som är nödvändiga för att se till att byråns arbetsprogram genomförs, varje år utarbeta ett utkast till allmän rapport och lägga fram det för styrelsen, göra beräkningar av byråns intäkter och utgifter samt genomföra budgeten.
(13) Senast fem år från det att byrån inlett sin verksamhet bör styrelsen beställa en oberoende extern utvärdering för att bedöma i vilken utsträckning förordningen, byrån och dess arbetsmetoder bidragit till att etablera en hög sjösäkerhetsnivå och en hög nivå på förhindrandet av förorening från fartyg.
MÅL OCH UPPGIFTER
1. Genom denna förordning inrättas en europeisk sjösäkerhetsbyrå, (byrån), i syfte att skapa en hög, enhetlig och effektiv sjösäkerhetsnivå och en hög nivå på förhindrandet av förorening från fartyg inom gemenskapen.
Uppgifter
b) Den skall bistå kommissionen i arbetet med att effektivt genomföra gemenskapslagstiftningen om sjösäkerhet och förhindrande av förorening från fartyg i hela gemenskapen. Byrån skall särskilt
iii) bistå kommissionen i genomförandet av de arbetsuppgifter som den har tilldelats av kommissionen genom befintlig och kommande gemenskapslagstiftning om sjösäkerhet och förhindrande av förorening från fartyg, särskilt lagstiftning om klassificeringssällskap, säkerheten på passagerarfartyg, säkerheten för fartygsbesättningar samt sjöfolks utbildning, certifiering och vakthållning.
ii) utveckla tekniska lösningar och ge tekniskt stöd avseende genomförandet av gemenskapslagstiftningen.
ii) utveckla och sköta de informationssystem som är nödvändiga för att uppnå det direktivets syften.
g) Under förhandlingarna med de stater som ansöker om anslutning får byrån tillhandahålla tekniskt stöd för genomförandet av gemenskapslagstiftningen om sjösäkerhet och förhindrande av förorening från fartyg. Denna uppgift skall samordnas med befintliga regionala samarbetsprogram och vid behov omfatta anordnande av relevant utbildningsverksamhet.
1. För att sköta sina uppgifter får byrån genomföra besök i medlemsstaterna i enlighet med de riktlinjer som styrelsen fastställt. Medlemsstaternas nationella myndigheter skall underlätta arbetet för byråns personal.
Artikel 4
2. Byrån får på eget initiativ kommunicera på de områden som ingår i dess uppdrag. Den skall särskilt se till att allmänheten och alla berörda parter snabbt får objektiv, tillförlitlig och lättbegriplig information om dess arbete.
KAPITEL II
Rättslig status, regionala centrum
3. På begäran från kommissionen och med samtycke från de berörda medlemsstaterna får styrelsen besluta att inrätta de regionala centrum som byrån behöver för att kunna utföra de arbetsuppgifter avseende övervakning av navigation och sjötrafik som anges i direktiv 2002/59/EG.
Personal
3. Byråns personal skall bestå av tjänstemän som utsetts eller avdelats temporärt av kommissionen eller medlemsstaterna och av andra anställda som vid behov skall anställas av byrån för att fullgöra dess uppgifter.
Byrån och dess personal skall omfattas av protokollet om Europeiska gemenskapernas immunitet och privilegier.
1. Byråns avtalsrättsliga ansvar skall regleras av den lagstiftning som är tillämplig på avtalet i fråga.
4. Domstolen skall vara behörig att avgöra tvister om sådant skadestånd som avses i punkt 3.
Språk
Artikel 10
2. Styrelsen skall
c) inom ramen för utarbetandet av arbetsprogrammet behandla ansökningar från medlemsstater om tekniskt stöd enligt artikel 2 c ii,
e) anta byråns slutliga budget innan räkenskapsåret börjar och vid behov anpassa den till gemenskapens bidrag och byråns övriga intäkter,
h) utföra de av sina åligganden som hör samman med byråns budget i enlighet med artiklarna 18, 19 och 21,
Artikel 11
Styrelseledamöter skall utses på grundval av relevant erfarenhet och sakkunskap inom området för sjösäkerhet och förhindrande av förorening från fartyg.
4. I förekommande fall skall deltagande av företrädare för tredje land och villkoren för detta fastställas genom de förfaranden som avses i artikel 17.2.
1. Styrelsen skall utse en ordförande och en vice ordförande bland sina ledamöter. Vice ordföranden skall automatiskt ersätta ordföranden om denne är förhindrad att fullgöra sina åligganden.
Sammanträden
3. Styrelsen skall hålla två ordinarie sammanträden per år. Den skall dessutom sammanträda på initiativ av ordföranden eller på begäran av kommissionen eller en tredjedel av medlemsstaterna.
6. Styrelseledamöterna får, med förbehåll för bestämmelserna i arbetsordningen, biträdas av rådgivare eller experter.
Röstning
I en ledamots frånvaro skall suppleanten ha rätt att utöva dennes rösträtt.
Den verkställande direktörens arbetsuppgifter och befogenheter
a) Han/hon skall utarbeta arbetsprogrammet och lägga fram det för styrelsen efter samråd med kommissionen. Han/hon skall vidta nödvändiga åtgärder för att genomföra programmet. Han/hon skall besvara alla ansökningar om stöd från någon medlemsstat i enlighet med artikel 10.2 c eller från kommissionen.
d) Han/hon skall organisera ett effektivt övervakningssystem för att kunna jämföra byråns resultat med verksamhetens mål. På grundval därav skall den verkställande direktören varje år utarbeta ett utkast till allmän rapport och lägga fram det för styrelsen. Han/hon skall fastställa förfaranden för regelbunden utvärdering baserade på erkända branschnormer.
3. Den verkställande direktören får biträdas av en eller flera enhetschefer. Om den verkställande direktören är frånvarande eller har förhinder, skall han/hon ersättas av någon av enhetscheferna.
1. Byråns verkställande direktör skall utnämnas av styrelsen på grundval av meriter, dokumenterad skicklighet i förvaltning och ledarskap samt kompetens och erfarenheter som är relevanta för sjösäkerhet och förhindrande av förorening från fartyg. Styrelsen skall fatta sitt beslut med fyra femtedels majoritet av alla ledamöter som har rösträtt. Kommissionen får föreslå en eller flera kandidater.
Artikel 17
2. Inom ramen för dessa avtal skall förfaranden utarbetas genom vilka bl.a. skall fastställas karaktären och omfattningen av de detaljerade bestämmelserna för dessa länders deltagande i byråns arbete, inbegripet bestämmelser om ekonomiska bidrag och personal.
Artikel 18
a) bidrag från gemenskapen,
2. Byråns utgifter skall omfatta kostnader för personal, administration, infrastruktur och drift.
5. Styrelsen skall senast den 30 april varje år anta ett budgetförslag, tillsammans med ett preliminärt arbetsprogram, och överlämna det till kommissionen och de tredjeländer som deltar i byråns arbete i enlighet med artikel 17.
Artikel 19
2. Kontroll av byråns åtaganden, betalningar av alla utgifter samt kontroll av alla intäkters existens och inkassering av alla intäkter skall utföras av kommissionens styrekonom.
4. Europaparlamentet skall på styrelsens rekommendation bevilja byråns verkställande direktör ansvarsfrihet för genomförandet av budgeten.
1. För bekämpning av bedrägeri, korruption och annan olaglig verksamhet skall bestämmelserna i Europaparlamentets och rådets förordning (EG) nr 1073/1999 tillämpas utan begränsning när det gäller byrån.
Artikel 21
KAPITEL IV
Utvärdering
3. Styrelsen skall ta emot utvärderingen och utfärda rekommendationer till kommissionen om hur förordningen, byrån och dess arbetsmetoder eventuellt bör ändras. Utvärderingsresultatet och rekommendationerna skall överlämnas av kommissionen till Europaparlamentet och rådet samt offentliggöras.
Byrån skall vara verksam senast tolv månader efter det att förordningen trätt i kraft.
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
av den 3 oktober 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 152.4 b i detta,
efter att ha hört Regionkommittén,
(1) I rådets direktiv 90/667/EEG av den 27 november 1990 om fastställande av veterinära bestämmelser om bortskaffande och bearbetning av animaliskt avfall och dess utsläppande på marknaden samt om förhindrande av sjukdomsalstrande organismer i foder av animaliskt ursprung samt om ändring av direktiv 90/425/EEG(4) fastställs principen att alla typer av animaliskt avfall, oavsett källa, efter lämplig behandling får användas för produktion av foderråvaror.
(4) Mot bakgrund av de senaste årens erfarenheter är det lämpligt att klargöra förhållandet mellan direktiv 90/667/EEG och gemenskapens miljölagstiftning. Denna förordning bör inte påverka tillämpningen av gällande miljölagstiftning eller förhindra utarbetandet av nya regler om miljöskydd, särskilt inte när det gäller biologiskt nedbrytbart avfall. I detta avseende har kommissionen åtagit sig att i slutet av 2004 utarbeta ett direktiv om bioavfall, inklusive matavfall, och vars syfte kommer att vara dels att fastställa bestämmelser om användning, återvinning, återanvändning och omhändertagande av detta avfall, dels att kontrollera eventuella föroreningar.
(7) Vetenskapliga utlåtanden pekar på att utfodring av en djurart med protein som härrör från kroppar, eller delar av kroppar, från samma djurart medför risk för spridning av sjukdomar. Som en försiktighetsåtgärd bör sådan utfodring således förbjudas. Genomförandebestämmelser bör antas för att säkerställa nödvändigt avskiljande av animaliska biprodukter avsedda för användning i foder i alla bearbetnings-, lagrings- och transportstadier. Det bör emellertid finnas utrymme för undantag från detta allmänna förbud för fisk och pälsdjur, om vetenskapliga utlåtanden motiverar detta.
(10) För att eliminera risken för att patogener och/eller restsubstanser av ämnen sprids bör animaliska biprodukter bearbetas, lagras och hållas avskilda i godkända och övervakade anläggningar som den berörda medlemsstaten utsett, eller bortskaffas på lämpligt sätt. I vissa fall kan en bearbetnings-, förbrännings- eller samförbränningsanläggning som ligger i en annan medlemsstat användas, särskilt när detta är motiverat på grund av avstånd, transporttid eller kapacitetsproblem.
(13) Undantag från reglerna för användning av animaliska biprodukter kan vara lämpliga för att underlätta utfodring av djur som inte är avsedda att användas som livsmedel. De behöriga myndigheterna bör övervaka sådan användning.
(16) Gemenskapens hälsolagstiftning bygger på etablerade vetenskapliga rön. De behöriga vetenskapliga kommittéer som inrättats genom kommissionens beslut 97/404/EG(7) och 97/579/EG(8) bör därför alltid vid behov höras. I synnerhet behövs det ytterligare vetenskapliga utlåtanden om användning av produkter av animaliskt ursprung i organiska gödningsmedel och jordförbättringsmedel. I avvaktan på att gemenskapsregler antas mot bakgrund av dessa utlåtanden, får medlemsstaterna behålla eller anta nationella regler som är strängare än de som återfinns i denna förordning om dessa regler överensstämmer med annan tillämplig gemenskapslagstiftning.
(19) Animaliska biprodukter som inte är avsedda att användas som livsmedel (särskilt bearbetat animaliskt protein, utsmält fett, sällskapsdjursfoder, hudar, skinn och ull) finns upptagna i produktförteckningen i bilaga I till fördraget. För vissa delar av jordbruksbefolkningen utgör avyttringen av sådana produkter en viktig inkomstkälla. För att säkerställa att denna sektor utvecklas på ett ändamålsenligt sätt och kan öka sin produktion, bör det fastställas hälsobestämmelser för människor och djur för dessa produkter på gemenskapsnivå. Med tanke på att djur lätt smittas av olika sjukdomar bör särskilda krav gälla när animaliska biprodukter släpps ut på marknaden, särskilt i regioner med hög hälsostatus.
(22) Det lämpligaste sättet för den behöriga myndigheten på destinationsorten att få garantier för att en sändning med animaliska produkter uppfyller bestämmelserna i denna förordning är via det dokument som skall åtfölja en sådan sändning. Hälsointyget bör sparas för att det skall vara möjligt att kontrollera vart vissa importerade produkter sänds.
(25) En sådan förenkling kommer att leda till större öppenhet när det gäller vissa hälsobestämmelser om sådana animaliska produkter som inte är avsedda som livsmedel. En förenkling av detaljbestämmelserna i hälsolagstiftningen får dock inte leda till att området avregleras. Det är därför nödvändigt att behålla och, för att garantera människors och djurs hälsa, skärpa de detaljerade hälsobestämmelserna för animaliska produkter som inte är avsedda som livsmedel.
(28) Direktiv 90/667/EEG, rådets beslut 95/348/EG av den 22 juni 1995 om fastställande av veterinära bestämmelser och djurhälsobestämmelser gällande Förenade kungariket och Irland för bearbetning av vissa typer av avfall avsedda att saluföras lokalt som foder för vissa kategorier av djur(13) och rådets beslut 1999/534/EG av den 19 juli 1999 om åtgärder för bearbetning av visst animaliskt avfall till skydd mot transmissibel spongiform encefalopati och om ändring av kommissionens beslut 97/735/EG(14) bör därför upphävas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Denna förordning skall inte tillämpas på följande:
c) Hela kroppar eller delar från vilda djur som inte misstänks vara infekterade med sjukdomar som kan överföras till människor eller djur, med undantag av fisk som fiskas i kommersiellt syfte och kroppar eller delar av vilda djur som används för att tillverka jakttroféer.
i) härrör från transportmedel i internationell trafik,
f) Ägg, embryon och sperma avsedda för avel.
Artikel 2
a) animaliska biprodukter: hela kroppar eller delar från djur eller animaliska produkter som avses i artiklarna 4-6 som inte är avsedda att användas som livsmedel, inbegripet ägg, embryon och sperma.
d) kategori 3-material: animaliska biprodukter som avses i artikel 6.
g) vilda djur: djur som inte hålls av människor.
j) utsläppande på marknaden: all verksamhet som syftar till att sälja sådana animaliska biprodukter eller därav framställda produkter som omfattas av denna förordning till tredje man i gemenskapen eller varje annan form av överlåtelse mot betalning eller utan motprestation till sådan tredje man eller lagring för leverans till sådan tredje man.
m) producent: alla producenter vars verksamhet genererar animaliska biprodukter.
2. De särskilda definitionerna i bilaga I skall också gälla.
1. Animaliska biprodukter och produkter som framställts av dessa skall samlas in, transporteras, lagras, hanteras, bearbetas, bortskaffas, släppas ut på marknaden, exporteras, transiteras och användas i enlighet med denna förordning.
Artikel 4
ii) Djur som avlivats som ett led i utrotningen av TSE.
v) Vilda djur som misstänks vara infekterade med sjukdomar som kan överföras till människor eller djur.
c) Produkter framställda från djur som tillförts ämnen som är förbjudna enligt direktiv 96/22/EG samt produkter av animaliskt ursprung som innehåller rest av miljöföroreningar och andra ämnen som förtecknas i grupp B.3 i bilaga I till rådets direktiv 96/23/EG av den 29 april 1996 om införande av kontrollåtgärder för vissa ämnen och restsubstanser av dessa i levande djur och i produkter framställda därav och om upphävande av direktiv 85/358/EEG och 86/469/EEG samt beslut 89/187/EEG och 91/664/EEG(19), om restsubstanserna av dessa ämnen överskrider de gränsvärden som fastställs i gemenskapens lagstiftning eller, om gemenskapsgränsvärden saknas, i nationell lagstiftning.
f) Blandningar av kategori 1-material med antingen kategori 2-material eller kategori 3-material eller med båda, inbegripet allt material som är avsett för bearbetning i en bearbetningsanläggning för kategori 1-material.
b) bearbetas enligt någon av metoderna 1-5 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, eller enligt metod 1 om den behöriga myndigheten kräver detta, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI och slutligen bortskaffas som avfall genom förbränning eller samförbränning i en förbrännings- eller samförbränningsanläggning som godkänts i enlighet med artikel 12,
e) mot bakgrund av nya vetenskapliga rön bortskaffas med någon annan metod som godkänts i enlighet med förfarandet i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén. Denna metod kan antingen komplettera eller ersätta de metoder som föreskrivs i punkterna a-d.
Artikel 5
a) Naturgödsel och mag- och tarminnehåll.
d) Produkter av animaliskt ursprung utom, kategori 1-material, som importeras från tredje land och som under sådana inspektioner som föreskrivs i gemenskapslagstiftningen inte uppfyller veterinärmedicinska bestämmelser för import till gemenskapen, om de inte återsänds eller importen godtas med vissa förbehåll som fastställts i gemenskapslagstiftningen.
g) Animaliska biprodukter som inte består av kategori 1- eller kategori 3-material.
b) bearbetas enligt någon av metoderna 1-5 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, eller om den behöriga myndigheten kräver detta, enligt bearbetningsmetod 1, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI, och
c) bearbetas enligt bearbetningsmetod 1 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI, och
iii) bortskaffas som avfall genom nedgrävning på en deponi som godkänts i enlighet med direktiv 1999/31/EG,
i) användas utan föregående bearbetning som råvara i en biogas- eller komposteringsanläggning som godkänts i enlighet med artikel 15 eller behandlas i en teknisk anläggning som godkänts för detta ändamål i enlighet med artikel 18,
f) när det gäller hela kroppar eller delar från vilda djur som inte misstänks vara infekterade med sjukdomar som kan överföras till människor eller djur, användas för att tillverka jakttroféer i en teknisk anläggning som godkänts för detta ändamål i enlighet med artikel 18, eller
4. Kategori 2-material får endast släppas ut på marknaden eller exporteras i enlighet med denna förordning eller enligt regler som fastställts i enlighet med förfarandet i artikel 33.2.
1. Kategori 3-material skall omfatta animaliska biprodukter som motsvarar följande beskrivning och allt material som innehåller sådana biprodukter:
c) Hudar, skinn, hovar, horn, svinborst och fjädrar från djur som slaktas i ett slakteri och som har genomgått en före slaktbesiktning där de befunnits lämpade för slakt för att användas som livsmedel i enlighet med gemenskapslagstiftningen.
f) Livsmedel av animaliskt ursprung eller som innehåller produkter av animaliskt ursprung, med undantag av matavfall, som inte längre är avsedda att användas som livsmedel av kommersiella skäl eller på grund av tillverkningsproblem eller förpackningsdefekter eller andra defekter som inte innebär någon risk för människor eller djur.
i) Färska biprodukter från fisk från anläggningar som tillverkar fiskprodukter som är avsedda att användas som livsmedel.
l) Matavfall, med undantag av matavfall enligt artikel 4.1 e.
b) bearbetas i en bearbetningsanläggning som godkänts i enlighet med artikel 13 med tillämpning av någon av bearbetningsmetoderna 1-5, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI och bortskaffas som avfall, antingen genom förbränning eller samförbränning i en förbrännings- eller samförbränningsanläggning som godkänts i enlighet med artikel 12, eller på en deponi som godkänts i enlighet med direktiv 1999/31/EG,
e) användas som råvara i en anläggning för framställning av sällskapsdjursfoder som godkänts i enlighet med artikel 18,
h) när det gäller material som kommer från fisk, ensileras eller komposteras i enlighet med bestämmelser som fastställts enligt förfarandet i artikel 33.2, eller
Artikel 7
2. Under transporten skall ett handelsdokument, eller, när det krävs enligt denna förordning, ett hälsointyg åtfölja animaliska biprodukter och bearbetade produkter. Handelsdokument och hälsointyg skall uppfylla de krav och bevaras under den tid som anges i bilaga II. De skall särskilt innehålla uppgifter om mängden och en beskrivning av materialet och dess märkning.
5. Bearbetade produkter får endast lagras vid lagringsanläggningar som godkänts enligt artikel 11.
Avsändande av animaliska biprodukter och bearbetade produkter till andra medlemsstater
3. Animaliska biprodukter och de bearbetade produkter som avses i punkt 2 skall
4. När medlemsstater sänder kategori 1-material, kategori 2-material, bearbetade produkter som härrör från kategori 1- eller kategori 2-material och bearbetat animaliskt protein till andra medlemsstater skall den behöriga myndigheten på ursprungsorten underrätta den behöriga myndigheten på bestämmelseorten om varje avgående sändning via Animo-systemet, eller med hjälp av någon annan överenskommen metod. Meddelandet skall innehålla de upplysningar som anges i kapitel I.2 i bilaga II.
Artikel 9
Artikel 10
2. För att kunna godkännas skall ett hanteringsställe för kategori 1- eller kategori 2-material
c) genomgå hanteringsställets egenkontroll på det sätt som föreskrivs i artikel 25,
a) uppfylla kraven i kapitel I i bilaga III,
d) kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
1. Lagringsanläggningar skall godkännas av den behöriga myndigheten.
b) ha kontrollerats av den behöriga myndigheten i enlighet med artikel 26.
1. Förbränning och samförbränning av bearbetade produkter skall genomföras i enlighet med bestämmelserna i direktiv 2000/76/EG. Förbränning och samförbränning av animaliska biprodukter skall antingen genomföras i enlighet med bestämmelserna i direktiv 2000/76/EG eller, då det direktivet inte är tillämpligt, i enlighet med bestämmelserna i denna förordning. Förbrännings- och samförbränningsanläggningar skall godkännas i enlighet med det direktivet eller i enlighet med punkt 2 eller 3.
b) villkoren för verksamheten i kapitel II i bilaga IV,
e) temperaturmätningskraven i kapitel V i bilaga IV,
a) användas endast för bortskaffande av döda sällskapsdjur och/eller kategori 2- och kategori 3-material,
d) uppfylla de tillämpliga villkoren för verksamheten i kapitel II i bilaga IV,
g) uppfylla kraven för onormala driftsförhållanden i kapitel VI i bilaga IV.
Artikel 13
2. För att kunna godkännas skall bearbetningsanläggningar för kategori 1- eller kategori 2-material
c) valideras av den behöriga myndigheten i enlighet med kapitel V i bilaga V,
f) kunna säkerställa att de bearbetade produkterna uppfyller kraven i kapitel I i bilaga VI.
Godkännande av oleokemiska anläggningar för kategori 2- och kategori 3-material
b) införa och genomföra rutiner för övervakning och kontroll av kritiska kontrollpunkter i de processer som används,
3. För att kunna godkännas skall en oleokemisk anläggning för kategori 3-material bearbeta utsmält fett som härrör endast från kategori 3-material och uppfylla de relevanta kraven i punkt 2.
Godkännande av biogas- och komposteringsanläggningar
a) uppfylla kraven i kapitel II del A i bilaga VI,
d) införa och genomföra rutiner för övervakning och kontroll av kritiska kontrollpunkter,
Artikel 16
2. De åtgärder som avses i punkt 1 skall säkerställa att produkterna har framställts från djur som
3. Förutsatt att de villkor som gäller sådana åtgärder för sjukdomsbekämpning som avses i punkt 2 a är uppfyllda, skall det vara tillåtet att på marknaden släppa ut animaliska biprodukter, och sådana därav framställda produkter som avses i bilagorna VII och VIII, som kommer från ett område eller en del av ett område som är föremål för djurhälsorestriktioner men som inte är infekterade eller misstänks vara infekterade, förutsatt att produkterna, allt efter omständigheterna
c) har identifierats på ett korrekt sätt,
Artikel 17
2. För att kunna godkännas skall en bearbetningsanläggning för kategori 3-material
c) valideras av den behöriga myndigheten i enlighet med kapitel V i bilaga V,
f) kunna säkerställa att de bearbetade produkterna uppfyller kraven i kapitel I i bilaga VII.
Godkännande av anläggningar för tillverkning av sällskapsdjursfoder och av tekniska anläggningar
a) I enlighet med de särskilda kraven i bilaga VIII för de produkter som anläggningen framställer skall den åta sig att
iii) beroende på vilken produkt det gäller, ta prover som sedan analyseras på ett laboratorium som godkänts av den behöriga myndigheten, så att det kan kontrolleras att kraven i denna förordning är uppfyllda,
b) Anläggningen skall kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
Utsläppande på marknaden och export av bearbetat animaliskt protein och andra bearbetade produkter som skulle kunna användas som foderråvara
b) har framställts enbart av sådant kategori 3-material som förtecknas i bilaga VII,
Artikel 20
a) antingen
b) kommer från anläggningar som har godkänts och står under tillsyn i enlighet med artikel 18 eller, när det gäller de animaliska biprodukter som avses i bilaga VIII, från andra anläggningar som har godkänts i enlighet med gemenskapens veterinärlagstiftning.
a) har framställts av utsmält fett som kommer från bearbetning av kategori 2-material i en bearbetningsanläggning för kategori 2-material som godkänts i enlighet med artikel 13 med tillämpning av någon av bearbetningsmetoderna 1-5 i en oleokemisk anläggning för kategori 2-material som har godkänts i enlighet med artikel 14,
Artikel 21
Artikel 22
a) Utfodring av ett djurslag med animaliskt protein som härrör från djurkroppar eller delar av djur av samma art.
2. Genomförandebestämmelser till denna artikel, inbegripet bestämmelser som rör kontrollåtgärder, skall antas i enlighet med det förfarande som avses i artikel 33.2. Undantag från punkt 1 a får beviljas för fisk och pälsdjur i enlighet med samma förfarande, efter samråd med den berörda vetenskapliga kommittén.
1. Medlemsstaterna får, under de behöriga myndigheternas tillsyn, godkänna följande:
2. a) Medlemsstaterna får även godkänna användning av de animaliska biprodukter som anges i stycke b för utfodring av de djur som anges i stycke c under de behöriga myndigheternas tillsyn och i enlighet med reglerna i bilaga IX.
ii) Kategori 3-material som avses i artikel 6.1 a-6.1 j och, om inte annat följer av artikel 22, i artikel 6.1 l.
ii) cirkusdjur,
v) vilda djur vars kött inte är avsett som livsmedel,
d) Medlemsstaterna får dessutom, under de behöriga myndigheternas tillsyn, tillåta användning av sådant kategori 1-material som avses i artikel 4.1 b ii för utfodring av utrotningshotade eller skyddade arter av asätande fåglar enligt regler som har fastställts i enlighet med det förfarande som anges i artikel 33.2, efter samråd med Europeiska myndigheten för livsmedelssäkerhet.
b) de kontroller som införs för att säkerställa att de animaliska biprodukterna i fråga endast används för godkända ändamål.
Om det vid en sådan inspektion visar sig att dessa krav inte har uppfyllts skall den behöriga myndigheten vidta lämpliga åtgärder.
Undantag i fråga om bortskaffande av animaliska biprodukter
b) följande animaliska biprodukter med ursprung i avlägsna områden får bortskaffas som avfall genom förbränning eller nedgrävning på platsen:
iii) kategori 3-material,
3. När det gäller kategori 1-material som avses i artikel 4.1 b ii får förbränning och nedgrävning utföras i enlighet med punkt 1 b eller c endast om den behöriga myndigheten godkänner och övervakar den metod som används och är övertygad om att den utesluter varje risk för överföring av TSE.
b) vilka områden de kategoriserar som avlägsna områden vid tillämpning av punkt 1 b och skälen till denna kategorisering.
b) hindra att animaliska biprodukter överges, dumpas eller bortskaffas på ett okontrollerat sätt.
Anläggningarnas egenkontroll
b) införa och genomföra rutiner för övervakning och kontroll av sådana kritiska kontrollpunkter i processen,
ii) ligger inom de gränsvärden för fysisk-kemiska restsubstanser som anges i gemenskapslagstiftningen,
2. Om resultatet av ett test som utförts på ett prov som tagits enligt punkt 1 c inte uppfyller bestämmelserna i denna förordning skall den ansvarige för bearbetningsanläggningen
c) under den behöriga myndighetens tillsyn bortskaffa den kontaminerade satsen eller låta den genomgå förnyad bearbetning,
f) granska de register över obearbetade animaliska biprodukter som är av betydelse för det färdiga provet,
Artikel 26
2. Hur ofta inspektioner och tillsyn skall genomföras beror på anläggningens storlek, vilken typ av produkter som tillverkas, vilka riskbedömningar som gjorts samt vilka garantier som lämnats i enlighet med principerna för systemet för riskbedömning och kritiska kontrollpunkter (HACCP).
5. Närmare bestämmelser för genomförandet av denna artikel, inbegripet regler om hur ofta kontroller skall ske och om referensmetoder för mikrobiologiska analyser, får fastställas i enlighet med det förfarande som avses i artikel 33.2.
1. Experter från kommissionen får, när så krävs för en enhetlig tillämpning av denna förordning, i samarbete med de behöriga myndigheterna i medlemsstaterna genomföra kontroller på plats. Den medlemsstat på vars territorium en inspektion företas skall ge all nödvändig hjälp till experterna så att de kan fullgöra sina uppgifter. Kommissionen skall informera den behöriga myndigheten om resultaten av de genomförda kontrollerna.
De bestämmelser som skall tillämpas vid import från tredje land av de produkter som avses i bilagorna VII och VIII får varken vara fördelaktigare eller mindre fördelaktiga än de som gäller för produktion och saluföring av motsvarande produkter i gemenskapen.
Förbud och efterlevnad av gemenskapsbestämmelser
3. De produkter som avses i bilagorna VII och VIII skall, om inte något annat anges i dessa bilagor, komma från ett tredje land eller en del av ett tredje land som återfinns på en sådan förteckning som skall upprättas och uppdateras i enlighet med förfarandet i artikel 33.2.
a) Det tredje landets lagstiftning.
d) Vilka garantier det tredje landet kan ge för att gällande hygienkrav uppfylls.
g) Hälsostatus för livsmedelsproducerande djur samt för andra tamdjur och vilda djur i det tredje landet, med särskilt beaktande av exotiska djursjukdomar och alla sådana aspekter av den allmänna hälsosituationen i landet som skulle kunna innebära en risk för folk- eller djurhälsan i gemenskapen.
4. De produkter som avses i bilagorna VII och VIII, med undantag av tekniska produkter, skall komma från en anläggning som finns upptagen på en gemenskapsförteckning som upprättats i enlighet med det förfarande som avses i artikel 33.2, på grundval av ett meddelande till kommissionen från de behöriga myndigheterna i det tredje landet i vilket det intygas att anläggningen uppfyller gemenskapens krav och att officiella inspektörer i det tredje landet ansvarar för tillsynen av anläggningen.
b) Medlemsstaterna skall, inom sju arbetsdagar från det att de tagit emot de förslag till ändringar av förteckningen över anläggningar som avses i punkt a, skriftligen meddela kommissionen sina synpunkter på dessa förslag.
5. De tekniska produkter som avses i bilaga VIII skall komma från anläggningar som har godkänts och registrerats av de behöriga myndigheterna i det tredje landet.
Artikel 30
I beslutet skall fastställas vilka villkor som gäller för import och/eller transitering av animaliska biprodukter från denna region, detta land eller denna grupp av länder.
b) vilka särskilda hälsokrav som skall gälla för import till och/eller transitering genom gemenskapen,
Artikel 31
a) upprätta en förteckning över tredje länder eller delar av tredje länder samt för att fastställa villkor för import och/eller transitering,
ii) villkoren för import och/eller transitering,
De experter från medlemsstaterna som ansvarar för kontrollerna skall utses av kommissionen.
4. Om det vid en kontroll enligt punkt 1 uppdagas allvarliga överträdelser av hälsobestämmelserna, skall kommissionen omedelbart begära att det tredje landet vidtar lämpliga åtgärder eller tillfälligt stoppa sändningarna av produkter och genast underrätta medlemsstaterna.
1. Efter samråd med berörd vetenskaplig kommitté i frågor som kan ha betydelse för djurs och människors hälsa får bilagorna ändras eller kompletteras och lämpliga övergångsbestämmelser antas i enlighet med förfarandet i artikel 33.2.
Föreskrivande förfarande
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara 15 dagar.
Samråd med vetenskapliga kommittéer
Nationella bestämmelser
3. Medlemsstaterna får anta eller bibehålla nationella bestämmelser som i större utsträckning än denna förordning begränsar användningen av organiska gödningsmedel och jordförbättringsmedel i väntan på att gemenskapsregler skall antas för användningen av dessa medel, i enlighet med artikel 20.2. Medlemsstaterna får anta eller bibehålla nationella bestämmelser som i större utsträckning än denna förordning begränsar användningen av fettderivat som framställts ur kategori 2-material i avvaktan på ett tillägg till bilaga VIII av gemenskapsregler för deras användning i enlighet med artikel 32.
Kommissionen skall utarbeta en rapport om hur medlemsstaterna finansierar bearbetning, insamling, lagring och bortskaffande av animaliska biprodukter, och rapporten skall åtföljas av lämpliga förslag.
Direktiv 90/667/EEG samt besluten 95/348/EG och 1999/534/EG skall upphöra att gälla sex månader efter det att denna förordning trätt i kraft.
Ikraftträdande
av den 10 oktober 2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING,
av följande skäl:
(3) Under antagandeprocessen fastställdes emellertid inte något sådant datum.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
I artikel 2 i förordning (EG) nr 1282/2002 skall följande läggas till som andra stycke: "Den skall tillämpas från och med den 1 mars 2003."
Rådets förordning (EG) nr 1881/2002
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(2),
(1) I enlighet med artikel 13.1 i rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(4) beviljades en övergångsperiod på två år, med början samma dag som ikraftträdandet, under vilken bestämmelserna i avdelning IV i ovannämnda förordning skulle gälla, till producentorganisationer som erkänts enligt förordning (EEG) nr 1035/72(5), men som inte uppfyllde kraven för erkännande enligt förordning (EG) nr 2200/96. Denna tvååriga övergångsperiod kan förlängas till fem år om medlemsstaten i fråga godkänner en handlingsplan som läggs fram av producentorganisationen över hur denna skall uppfylla kraven i förordning (EG) nr 2200/96 för att erkännas av den medlemsstaten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 28 oktober 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Enligt artikel 3 i kommissionens förordning (EEG) nr 3149/92(3), senast ändrad genom förordning (EEG) nr 1098/2001(4), skall den årliga planen för utdelning av livsmedel till de sämst ställda genomföras under perioden 1 oktober-30 september följande år. För att interventionslagren skall kunna förvaltas på bästa sätt bör de produkter som skall delas ut tas ut ur lagren senast den 31 augusti under genomförandeåret.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från berörda förvaltningskommittéer.
Förordning (EEG) nr 3149/92 ändras på följande sätt:
"Artikel 5
För de medlemsstater som inte har infört euron skall interventionsprodukternas bokföringsvärde omräknas till den nationella valutan med hjälp av den växelkurs som gällde den 1 oktober.
Artikel 2
av den 31 oktober 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) De belgiska och italienska myndigheterna har meddelat kommissionen att marknaderna i Antwerpen och Bologna inte längre är representativa importmarknader för frukt och grönsaker. Dessa marknader bör därför strykas från förteckningen i artikel 3.1 i kommissionens förordning (EG) nr 3223/94(3), senast ändrad genom förordning (EG) nr 453/2002(4).
"- Belgien och Luxemburg: Bryssel".
Artikel 2
av den 5 november 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2 i detta,
med beaktande av Regionkommitténs yttrande(3),
(1) Genomförandeåtgärderna i gällande förordningar och direktiv inom sjösäkerhetsområdet har antagits genom ett föreskrivande förfarande inom ramen för den kommitté som inrättas genom rådets direktiv 93/75/EEG av den 13 september 1993 om minimikrav för fartyg som anlöper eller avgår från gemenskapens hamnar med farligt eller förorenande gods(5) och i vissa fall en ad hoc-kommitté. Dessa kommittéer har styrts av reglerna i rådets beslut 87/373/EEG av den 13 juli 1987 om närmare villkor för utövandet av kommissionens genomförandebefogenheter(6).
(4) I enlighet med resolutionen av den 8 juni 1993 bör en kommitté för sjösäkerhet och förhindrande av förorening från fartyg inrättas och tilldelas de uppgifter som tidigare hört till de kommittéer som inrättats inom ramen för nämnda lagstiftning. All ny gemenskapslagstiftning som antas inom sjösäkerhetsområdet bör innehålla hänvisning till denna kommitté.
(7) Nämnda lagstiftning bör också ändras så att COSS ersätter den kommitté som inrättats genom direktiv 93/75/EEG eller, i förekommande fall, den ad hoc-kommitté som inrättas genom en viss rättsakt. Genom denna förordning bör framför allt relevanta bestämmelser i rådets förordningar (EEG) nr 613/91 av den 4 mars 1991 om överflyttning av fartyg från ett register till ett annat inom gemenskapen(9), (EG) nr 2978/94 av den 21 november 1994 om genomförande av IMO-resolution A.747(18) om tillämpningen av mätning av dräktighet av barlastutrymmen i oljetankfartyg med segregerade barlasttankar(10) och (EG) nr 3051/95 av den 8 december 1995 om säkerhetsorganisation för roll-on/roll-off-passagerarfartyg (ro-ro-fartyg)(11) samt Europaparlamentets och rådets förordning (EG) nr 417/2002 av den 18 februari 2002 om ett påskyndat införande av krav på dubbelskrov eller likvärdig konstruktion för oljetankfartyg med enkelskrov och om upphävande av rådets förordning (EG) nr 2978/94(12) ändras för infogande av en hänvisning till COSS och för tillämpning av det föreskrivande förfarande som anges i artikel 5 i beslut 1999/468/EG.
(10) Medlemsstaterna bör därför tillåtas att tillämpa de senaste bestämmelserna i de internationella instrumenten, med undantag för bestämmelser som redan uttryckligen ingår i en gemenskapsrättsakt. Detta kan uppnås genom att man anger att den version av den internationella konvention som skall beaktas för det berörda direktivet eller den berörda förordningen skall vara "i gällande version", utan att ett datum anges.
(13) Förfarandet för kontroll av överensstämmelse kommer att få full verkan endast om de planerade åtgärderna antas så snart som möjligt, och under alla omständigheter innan den internationella ändringen träder i kraft. Följaktligen bör den tidsfrist som rådet enligt artikel 5.6 i beslut 1999/468/EG beviljas för att fatta beslut om förslag till åtgärder vara en månad.
Syfte
b) påskynda uppdateringen och underlätta senare ändringar av gemenskapens sjöfartslagstiftning mot bakgrund av utvecklingen av de internationella instrument som avses i artikel 2.1.
2. gemenskapens sjöfartslagstiftning: följande gällande gemenskapsrättsakter:
c) Rådets förordning (EG) nr 2978/94.
f) Rådets förordning (EG) nr 3051/95.
i) Rådets direktiv 98/18/EG av den 17 mars 1998 om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg.(17)
l) Europaparlamentets och rådets direktiv 2000/59/EG av den 27 november 2000 om mottagningsanordningar i hamn för fartygsgenererat avfall och lastrester.(20)
o) Europaparlamentets och rådets förordning (EG) nr 417/2002.
1. Kommissionen skall biträdas av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg, nedan kallad COSS.
3. Kommittén skall själv anta sin arbetsordning.
Gemenskapens sjöfartslagstiftning skall omfattas av de internationella instrument som har trätt i kraft, inbegripet de senaste ändringarna av dessa, med undantag för de ändringar som undantagits från tillämpningsområdet för gemenskapens sjöfartslagstiftning på grund av resultatet av det förfarande för kontroll av överensstämmelse som fastställs i artikel 5.
1. För att uppnå syftet med denna förordning och för att minska risken för en konflikt mellan gemenskapens sjöfartslagstiftning och internationella instrument skall medlemsstaterna och kommissionen samarbeta genom samordningsmöten och/eller på andra lämpliga sätt för att i förekommande fall fastställa en gemensam ståndpunkt eller strategi i behöriga internationella forum.
3. Om det föreligger sådana omständigheter som avses i punkt 2 skall förfarandet för kontroll av överensstämmelse inledas av kommissionen, eventuellt på begäran av någon medlemsstat.
4. Om en sådan risk som avses i punkt 2 första stycket föreligger skall medlemsstaterna under förfarandet för kontroll av överensstämmelse avhålla sig från varje initiativ som syftar till att genomföra ändringen i den nationella lagstiftningen eller tillämpa denna ändring av det internationella instrumentet i fråga.
Alla relevanta ändringar av de internationella instrument som är införlivade i gemenskapens sjöfartslagstiftning i enlighet med artiklarna 4 och 5 skall i informationssyfte offentliggöras i Europeiska gemenskapernas officiella tidning.
COSS skall utöva de befogenheter som den tilldelas i enlighet med gällande gemenskapslagstiftning. Artikel 2.2 får ändras genom det förfarande som anges i artikel 3.2 i syfte att infoga en hänvisning till gemenskapsrättsakter som trätt i kraft efter antagandet av denna förordning och enligt vilka COSS tillerkänns genomförandebefogenheter.
Förordning (EEG) nr 613/91 ändras på följande sätt:
2. Artiklarna 6 och 7 skall ersättas med följande:
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(24) tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 7
Ändring av förordning (EG) nr 2978/94
"g) Marpol 73/78: 1973 års internationella konvention till förhindrande av förorening från fartyg, i dess lydelse enligt det därtill hörande protokollet av år 1978, i gällande version."
"Artikel 7
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
Ändring av förordning (EG) nr 3051/95
2. Artikel 10 skall ersättas med följande:
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(28) tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 11
2. Artikel 10.1 skall ersättas med följande:
Artikel 12
av den 28 november 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Utvecklingen av tekniker och begrepp, i synnerhet vad gäller skillnaden mellan formell utbildning och andra former av undervisningsaktiviteter och genomförandet av klassificeringen av inriktningen av utbildningen, framtvingar en anpassning av förteckningen över variabler för utbildning som anges i artikel 4.1 h i förordning (EG) nr 577/98.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"h) Utbildning
- inriktning
- syfte för de senaste kurserna eller annan undervisningsaktivitet
utbildningsnivå
- år då denna utbildning framgångsrikt avslutades"
Artikel 3
av den 23 december 2002
(2003/8/EG)
med beaktande av rådets förordning (EEG) nr 1612/68 av den 15 oktober 1968 om arbetskraftens fria rörlighet inom gemenskapen(1), senast ändrad genom förordning (EEG) nr 2434/92(2), särskilt artikel 44 i denna, och
(2) Mot bakgrund av erfarenheterna sedan 1993 och för att beakta och befästa den nya utvecklingen av EURES-verksamheten, bör nätverket nu stärkas och fullt ut integreras i medlemsstaternas arbetsförmedlingsverksamhet. Den nuvarande ansvarsfördelningen och de nuvarande beslutsförfarandena bör få en ny utformning.
(5) EURES-nätverket bör därför befästas och stärkas som ett viktigt instrument för att övervaka den transnationella rörligheten, stödja arbetstagarnas fria rörlighet, integrera de europeiska arbetsmarknaderna och informera medborgarna om relevant gemenskapslagstiftning.
(8) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Tekniska kommittén för fri rörlighet för arbetstagare.
EURES-nätverket
Mål
a) utveckling av europeiska arbetsmarknader som är öppna och tillgängliga för alla,
d) utveckling av metoder och indikatorer för detta ändamål.
EURES-nätverket skall omfatta följande parter:
i) regionala arbetsförmedlingar i medlemsstaterna,
Dessa parter skall inbegripa de fackliga organisationer och arbetsgivarorganisationer som EURES medlemmar utser.
Kommissionens generaldirektorat för sysselsättning och socialpolitik skall ansvara för Europeiska samordningsbyrån.
a) analysera den geografiska och yrkesmässiga rörligheten och utarbeta en generell metod för transnationell rörlighet i enlighet med den europeiska sysselsättningsstrategin,
Artikel 5
Logotypen skall registreras som ett gemenskapsvarumärke vid Byrån för harmonisering inom den inre marknaden (varumärken och formgivning). Den får användas av EURES medlemmar och samarbetspartner.
En högnivågrupp för strategiska frågor inrättas härmed. Gruppen skall bestå av cheferna för EURES-medlemmarna och ha en företrädare för kommissionen som ordförande. Den skall bistå kommissionen med att främja och övervaka utvecklingen av EURES-nätverket.
b) EURES-nätverkets riktlinjer, enligt artikel 9.1,
Ledarna för arbetsmarknadsorganisationerna på EU-nivå skall inbjudas till att delta i gruppens möten.
Artikel 7
Artikel 8
2. Utifrån principen om att alla lediga platser och platsansökningar som offentliggörs av EURES medlemmar och samarbetspartner skall göras tillgängliga i hela Europeiska gemenskapen, skall EURES-stadgan särskilt innehålla följande information:
ii) utveckling av samarbetet mellan olika länder och i gränstrakter, inklusive arbetsförmedling och social service, arbetsmarknadens parter och andra institutioner som berörs, med sikte på att arbetsmarknaderna skall fungera bättre och integreras samt på att öka rörligheten,
i) integrering av medlemmarnas databaser för lediga platser i EURES-systemet för förmedling av lediga platser inom en tidsfrist som skall bestämmas,
iv) utarbetande, inlämnande till EURES samordningsbyrå och genomförande av verksamhetsplaner, med särskilda regler för EURES-verksamhet som bedrivs över gränserna,
c) Förfaranden för att upprätta ett enhetligt system och gemensamma former för utbyte av information om arbetsmarknaden och om transnationell rörlighet inom EURES-nätverket, i enlighet med artiklarna 14, 15 och 16 i förordning (EEG) nr 1612/68, inklusive information om lediga platser och utbildningsmöjligheter inom Europeiska unionen som skall integreras i en webbplats för information om rörlighet i arbetslivet.
1. I enlighet med den EURES-stadga som föreskrivs i artikel 8 och efter samråd med den högnivågrupp för strategiska frågor som avses i artikel 6, skall EURES samordningsbyrå fastställa riktlinjer för EURES-verksamheten för en period på tre år.
a) den huvudsakliga verksamhet som EURES-medlemmen skall bedriva inom ramen för nätverket, inklusive sådan transnationell, gränsöverskridande och branschspecifik verksamhet som avses i artikel 17 i förordning (EEG) nr 1612/68,
Verksamhetsplanerna skall även innehålla en utvärdering av verksamheten och de framsteg som gjorts under den föregående perioden.
Artikel 10
Artikel 11
Artikel 12
Europaparlamentets och rådets direktiv 2003/24/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) I syfte att harmonisera säkerhetsnivån för passagerarfartyg i hela gemenskapen bör det undantag som beviljats Grekland när det gäller tidtabellen för tillämpningen av säkerhetsbestämmelserna upphävas.
(6) Ändringar i relevanta internationella texter, t.ex. Internationella sjöfartsorganisationens (IMO) konventioner, protokoll, koder och resolutioner, måste kunna beaktas på ett flexibelt och snabbt sätt.
(9) Direktiv 98/18/EG bör därför ändras i enlighet med detta.
Direktiv 98/18/EG ändras enligt följande:
"ha) ålder: fartygets ålder uttryckt i antal år efter dess leveransdatum."
"2. Varje medlemsstat skall
c) till kommissionen anmäla var denna information finns och när förteckningen senast ändrades.".
Stabilitetskrav för och utfasning av ro-ro-passagerarfartyg
Artikel 6b
2. Medlemsstaterna skall samarbeta och samråda med organisationer som företräder personer med nedsatt rörlighet när det gäller genomförandet av riktlinjerna i bilaga III.
4. Medlemsstaterna skall senast den 17 maj 2006 rapportera till kommissionen om genomförandet av denna artikel beträffande alla passagerarfartyg som avses i punkt 1, de passagerarfartyg som avses i punkt 3 och som är certifierade för fler än 400 passagerare samt alla höghastighetspassagerarfartyg."
Artikel 6.3 g i direktiv 98/18/EG skall utgå med verkan från och med den 1 januari 2005.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
av den 3 april 2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
av följande skäl:
(3) Direktiv 96/96/EG har ändrats genom införande av skärpta utsläppsgränser för vissa kategorier av motorfordon och funktionsprovning av hastighetsbegränsande anordningar på tunga nyttofordon. Direktiv 2000/30/EG bör anpassas för att överensstämma med det direktivet genom att nya tekniska bestämmelser införs om att omborddiagnossystem och hastighetsbegränsande anordningar skall omfattas av vägkontrollerna. För att överensstämma med direktiv 96/96/EG, måste det införas nya tekniska bestämmelser i direktiv 2000/30/EG, vilket skall ske genom att omborddiagnossystem och hastighetsbegränsande anordningar skall omfattas av vägkontrollerna. Direktiv 2000/30/EG bör också uppdateras (tillsammans med direktiv 96/96/EG) så att det innehåller reviderade utsläppsgränsvärdena för vissa kategorier av motorfordon.
Artikel 1
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 2004. De skall genast underrätta kommissionen om detta.
Artikel 3
om främjande av användningen av biodrivmedel eller andra förnybara drivmedel
med beaktande av kommissionens förslag(1),
i enlighet med förfarandet i artikel 251 i fördraget(4), och
(2) Naturresurserna, som enligt artikel 174.1 i fördraget skall utnyttjas varsamt och rationellt, utgörs bland annat av olja, naturgas och fasta bränslen, vilka är viktiga energikällor, men de ger även upphov till de största koldioxidutsläppen.
(5) Kommissionen anger i sin vitbok "Den gemensamma transportpolitiken fram till 2010: Vägval inför framtiden" att koldioxidutsläppen från transportsektorn förväntas öka med 50 % mellan 1990 och 2010 till omkring 1113 miljoner ton, varvid vägtransporterna, som svarar för 84 % av de transportrelaterade koldioxidutsläppen, bär det tyngsta ansvaret. I vitboken ställs det därför av miljöskäl upp krav på att oljeberoendet (för närvarande 98 %) inom transportsektorn skall minskas genom användning av alternativa drivmedel, såsom biodrivmedel.
(8) Framsteg i tekniken har lett till att de flesta fordon som i dag är i bruk i Europeiska unionen utan problem kan använda en låg inblandning av biodrivmedel. De senaste tekniska framstegen gör det möjligt att använda högre halter av biodrivmedel i blandningen. I vissa länder används redan blandningar som innehåller halter av biodrivmedel på 10 % och däröver.
(11) Medlemsstaternas forskningspolitik om ökad användning av biodrivmedel bör i avsevärd utsträckning omfatta vätgassektorn och främja detta alternativ, och därvid beakta gemenskapens alla relevanta ramprogram.
(14) Bioetanol och biodiesel som i ren form eller i blandningar används i fordon bör uppfylla de kvalitetsstandarder som fastställts för att motorerna skall fungera optimalt. Det noteras att Europeiska standardiseringskommitténs standard prEN 14214 för fettsyrametylestrar (FAME) kan tillämpas i fråga om biodiesel för dieselmotorer, där tillverkningsalternativet är omförestring. Europeiska standardiseringskommittén bör sålunda fastställa lämpliga standarder för andra biodrivmedelsprodukter i Europeiska unionen.
(17) Kommissionens grönbok "Mot en europeisk strategi för trygg energiförsörjning" ställer upp målet att man senast år 2020 skall ha ersatt 20 % av konventionella drivmedel med alternativa drivmedel inom vägtransportsektorn.
(20) Den optimala metoden för att öka andelen biodrivmedel på de nationella marknaderna och gemenskapsmarknaderna är beroende av tillgången på resurser och råvaror, av den nationella politiken och gemenskapspolitiken för att främja biodrivmedel och av skattebestämmelser, samt av att alla intressenter/parter involveras på ett lämpligt sätt.
(23) Eftersom målet för den föreslagna åtgärden, nämligen införandet av allmänna principer för att en minimiandel biodrivmedel skall kunna marknadsföras och distribueras, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna på grund av åtgärdens omfattning och det därför bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå detta mål.
(26) Det bör föreskrivas ett förfarande för att snabbt anpassa förteckningen över biodrivmedel, andelen förnybart innehåll och tidsplanen för att införa biodrivmedel på transportmarknaden till den tekniska utvecklingen och till resultaten av en miljökonsekvensbedömning av den första introduktionsfasen.
(29) De åtgärder som är nödvändiga för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(7).
Syftet med detta direktiv är att främja användningen av biodrivmedel eller andra förnybara drivmedel som skall ersätta diesel eller bensin för transportändamål i varje medlemsstat, för att på så sätt bidra till mål som t.ex. att uppfylla åtaganden som rör klimatförändringar, bidra till försörjningstryggheten på ett miljövänligt sätt och främja förnybara energikällor.
a) biodrivmedel: flytande eller gasformigt bränsle för transport, som framställs av biomassa,
d) energiinnehåll: det nedre värmevärdet för ett drivmedel.
b) biodiesel: metylester av dieselkvalitet från vegetabilisk eller animalisk olja, som skall användas som biodrivmedel.
e) biodimetyleter: dimetyleter som framställs av biomassa och skall användas som biodrivmedel.
h) syntetiska biodrivmedel: syntetiska kolväten eller blandningar av syntetiska kolväten, som framställs av biomassa.
Artikel 3
ii) Ett referensvärde för dessa mål skall vara 5,75 %, beräknat på energiinnehållet, av all bensin och diesel för transportändamål som släpps ut på deras marknader, senast den 31 december 2010.
b) Biodrivmedel som blandats i mineraloljederivat i enlighet med de tillämpliga europeiska standarder som beskriver de tekniska specifikationerna för drivmedel (EN 228 och EN 590).
4. Medlemsstaterna bör i sina åtgärder ta hänsyn till vilken inverkan på den totala klimat- och miljöbalansen som de olika biodrivmedlen och andra förnybara drivmedel har och får prioritera främjandet av sådana drivmedel som ger en mycket god kostnadseffektiv miljöbalans med beaktande av konkurrenskraft och försörjningstrygghet.
1. Medlemsstaterna skall före den 1 juli varje år rapportera till kommissionen om
- det föregående årets totala försäljning av drivmedel samt andelen biodrivmedel, rena eller blandade, och andra förnybara drivmedel som släppts ut på marknaden. I förekommande fall skall medlemsstaterna rapportera om exceptionella förhållanden när det gäller utbudet av råolja eller oljeprodukter som har påverkat försäljningen av biodrivmedel och andra förnybara drivmedel.
a) Objektiva faktorer, t.ex. den begränsade nationella potentialen för produktion av biodrivmedel från biomassa.
2. Kommissionen skall senast den 31 december 2006 och vartannat år därefter utarbeta och till Europaparlamentet och rådet lämna en utvärderingsrapport om framstegen när det gäller användning av biodrivmedel och andra förnybara drivmedel i medlemsstaterna.
b) De ekonomiska aspekterna och miljökonsekvenserna av en ytterligare ökning av andelen biodrivmedel och andra förnybara drivmedel.
e) Bedömning av användningen av biodrivmedel och andra förnybara drivmedel med avseende på deras olika konsekvenser för klimatförändringen och deras påverkan när det gäller att minska koldioxidutsläppen.
Artikel 5
1. Kommissionen skall biträdas av en kommitté.
3. Kommittén skall själv anta sin arbetsordning.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska unionens officiella tidning.
Kommissionens direktiv 2003/60/EG
(Text av betydelse för EES)
med beaktande av rådets direktiv 76/895/EEG av den 23 november 1976 om fastställande av gränsvärden för bekämpningsmedelsrester i och på frukt och grönsaker(1), senast ändrat genom kommissionens direktiv 2002/79/EG(2), särskilt artikel 5 i detta,
med beaktande av rådets direktiv 90/642/EEG av den 27 november 1990 om fastställande av gränsvärden för bekämpningsmedelsrester i och på produkter av vegetabiliskt ursprung inklusive frukt och grönsaker(6), senast ändrat genom kommissionens direktiv 2002/100/EG, särskilt artikel 7 i detta,
(1) De befintliga verksamma ämnena amitrol, dikvat, isoproturon och etofumesat infördes i bilaga I till rådets direktiv 91/414/EEG genom kommissionens direktiv 2001/21/EG(9), 2002/18/EG(10) respektive 2002/37/EG(11).
(4) Om det inte finns något permanent eller provisoriskt gränsvärde för bekämpningsmedelsrester på gemenskapsnivå måste medlemsstaterna fastställa ett provisoriskt nationellt gränsvärde i enlighet med artikel 4.1 f i direktiv 91/414/EEG innan växtskyddsmedel som innehåller dessa verksamma ämnen kan godkännas.
(7) Gemenskapens gränsvärden och de värden som rekommenderas i Codex alimentarius fastställs och utvärderas genom liknande förfaranden. I Codex alimentarius anges ett begränsat antal gränsvärden för dikvat och fentin (-acetat eller -hydroxid). Dessa har beaktats vid fastställandet av de gränsvärden som anges i detta direktiv. De gränsvärden i Codex alimentarius som inom en nära framtid kommer att rekommenderas att dras tillbaka har inte beaktats. De gränsvärden som grundas på gränsvärden i Codex alimentarius har utvärderats med avseende på riskerna för konsumenterna, och inga risker kunde påvisas med de toxikologiska endpoints som var baserade på studier som var tillgängliga för kommissionen.
(10) Att provisoriska gränsvärden fastställs på gemenskapsnivå hindrar inte medlemsstaterna från att fastställa provisoriska gränsvärden för de ämnen som anges i det här direktivet i enlighet med artikel 4.1 f i direktiv 91/414/EEG och bilaga VI till det direktivet. Fyra år anses vara en tillräckligt lång period för att godkänna ytterligare användningsområden för de berörda verksamma ämnena. De provisoriska gränsvärdena bör därefter bli permanenta.
(13) Detta direktiv är förenligt med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
I bilaga II till direktiv 76/895/EEG skall posterna beträffande dikvat utgå.
Artikel 3
De gränsvärden för bekämpningsmedelsrester som anges i bilaga IV till detta direktiv skall läggas till i bilaga II till direktiv 90/642/EEG.
De skall tillämpa dessa bestämmelser från och med den 1 juli 2003, med undantag för bestämmelserna för fentinhydroxid, fentinacetat och klorfenapyr, som skall tillämpas från och med 1 juli 2004.
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska unionens officiella tidning.
Kommissionens förordning (EG) nr 568/2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
om ändring av Europaparlamentets och rådets förordning (EG) nr 999/2001 när det gäller snabbtest
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I förordning (EG) nr 999/2001 fastställs för tillämpningen av den förordningen en förteckning över nationella referenslaboratorier för TSE. Grekland har bytt nationellt referenslaboratorium.
(4) Vetenskapliga styrkommittén rekommenderade i sitt yttrande av den 6 och 7 mars 2003 att två nya test skulle införas i förteckningen över de snabbtest som godkänts för övervakning av bovin spongiform encefalopati (BSE). Tillverkarna av båda testen har presenterat data som visar att deras test också får användas för övervakning av TSE hos får.
(7) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
Bilaga X till förordning (EG) nr 999/2001 skall ändras i enlighet med bilagan till den här förordningen.
Kommissionens förordning (EG) nr 1139/2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Det finns en teoretisk möjlighet att bovin spongiform encefalopati (BSE) förekommer i får- och getpopulationen. Det är omöjligt att genom rutinmetoder skilja mellan BSE- och skrapiesmitta hos dessa djur. Infektiviteten i nedre delen av tunntarmen (ileum) är vid båda sjukdomarna signifikant redan i ett tidigt skede av infektionen. Som en förebyggande åtgärd bör ileum från får och getter i alla åldrar tillföras förteckningen över specificerat riskmaterial.
(6) Eftersom huvudets tillstånd huvudsakligen är beroende av att det hanteras varsamt och att skotthålet i pannan förseglas på ett säkert sätt liksom foramen magnum, måste det finnas kontrollsystem i slakterierna och i de styckningsanläggningar som särskilt godkänts.
(9) Förordning (EG) nr 999/2001 bör därför ändras.
Artikel 1
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
om ändring av rådets förordning (EG) nr 2223/96 med avseende på tidsfrister för sändningen av huvudaggregaten i nationalräkenskaperna, undantag när det gäller sändningen av huvudaggregaten i nationalräkenskaperna och sändning av uppgifter om sysselsättning angivna i arbetade timmar
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 285 i detta,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) I den rapport om statistiska krav i den ekonomiska och monetära unionen (EMU), som framlagts av Monetära kommittén, och som godkändes av Ekofinrådet den 18 januari 1999, framhålls att effektiv övervakning och samordning av den ekonomiska politiken är av största vikt för den inre marknaden, och att detta kräver ett omfattande statistiksystem genom vilket beslutsfattarna förses med ett nödvändigt beslutsunderlag. I rapporten talas också om vikten av att sådana uppgifter finns tillgängliga för gemenskapen, i synnerhet för de medlemsstater som deltar i euroområdet.
(5) Kvartalsvisa och årliga undantag som beviljats medlemsstaterna och som hindrar sammanställandet av huvudaggregaten i nationalräkenskaperna för euroområdet och gemenskapen bör avskaffas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Texten som följer på rubriken "Leveransprogram för nationalräkenskapsdata" skall ändras på följande sätt:
2. Texten som följer på rubriken: "Avvikelser beträffande de tabeller som skall sändas i enlighet med frågeformuläret "ESA-95" per land" skall ersättas med texten i bilaga III.
Kommissionens förordning (EG) nr 1914/2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
(1) I artikel 11.1 i förordning (EG) nr 3448/93 föreskrivs att de ekonomiska villkor som anges i artikel 117 c i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3), senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 2700/2000(4), skall betraktas som uppfyllda för att tillåta att vissa kvantiteter av vissa basprodukter får hänföras till förfarandet för aktiv förädling för att användas vid framställning av varor. De detaljerade tillämpningsföreskrifter till denna bestämmelse som gör det möjligt att fastställa vilka basjordbruksprodukter som får hänföras till förfarandet för aktiv förädling samt att kontrollera och planera kvantiteterna därav, skall antas i enlighet med artikel 16 i förordning (EG) nr 3448/93.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 2 skall punkt 2 ersättas av följande:
3. Artikel 24 skall ersättas av följande:
Kommissionens förordning (EG) nr 2151/2003
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Genom förordning (EG) nr 2195/2002 fastställdes ett enda klassificeringssystem för offentlig upphandling i syfte att standardisera de referenser som används av upphandlande myndigheter och enheter för att beskriva föremålet för upphandlingen.
(4) De tekniska ändringar och förbättringar som kartlagts under lagstiftningsprocessen inför antagandet av förordning (EG) nr 2195/2002 men som inte kunde tas med i den förordningen, bör införas i samma förordnings bilagor.
(7) Uppdateringen av CPV-koderna och CPV-strukturen bör även återspeglas i de vägledande konverteringstabellerna mellan CPV och FN:s centrala produktindelning (CPC Prov.), Europeiska gemenskapens statistiska näringsgrensindelning (NACE Rev. 1) och Kombinerade nomenklaturen (KN).
(10) I gemensam ståndpunkt (EG) nr 33/2003 antagen av rådet den 20 mars 2003 inför antagandet av Europaparlamentets och rådets direktiv om samordning av förfarandena vid offentlig upphandling av byggentreprenader, varor och tjänster(4) och gemensam ståndpunkt (EG) nr 34/2003, antagen av rådet den 20 mars 2003 inför antagandet av Europaparlamentets och rådets direktiv om samordning av förfarandena vid upphandling på områdena vatten, energi, transporter och posttjänster(5), fastställs inte varuområden efter den statistiska indelningen av produkter efter näringsgren (CPA).
(13) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Rådgivande kommittén för offentlig upphandling.
Förordning (EG) nr 2195/2002 skall ändras enligt följande:
Bilaga III skall ersättas med texten i bilaga III till denna förordning.
Artikel 2
av den 23 februari 2004
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Österrikes begäran av den 30 juni 2003,
av följande skäl,
(3) Åtgärderna som fastställs i den här förordningen överensstämmer med yttrandet från Kommittén för det statistiska programmet som inrättades genom rådets beslut 89/382/EEG, Euratom(2).
1. Följande undantag från bestämmelserna i förordning (EG) nr 2150/2002 beviljas härmed:
c) Luxemburg beviljas undantag för redovisning av resultat avseende avsnitt 8.1.1, posterna 1 (jordbruk, jakt och skogsbruk) och 2 (fiske) i bilaga I.
Artikel 2
