EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av följande: Antagandet av en gemensam transportpolitik innebär bland annat att man fastställer gemensamma regler för internationella godstransporter på väg till eller från en medlemsstat eller genom en eller flera medlemsstater.
Artikel 1
3. De typer av transporter som är förtecknade i bilaga 2 skall inte längre regleras av något kvoteringssystem. Dock får tillståndskrav behållas som villkor för denna transportverksamhet, förutsatt att ingen restriktion av kvantitativ natur förekommer; i sådant fall skall medlemsstaterna ombesörja att beslut i tillståndsärenden fattas senast fem dagar efter mottagandet av tillståndsansökan.
Medlemsstaterna skall senast tre månader efter detta direktivs ikraftträdande och i vart fall före utgången av år 1962 underrätta kommissionen om de åtgärder som vidtagits för att genomföra det.
Artikel 4
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Enligt artikel 17.4 i förordning nr 359/67/EEG får det exportbidrag som gäller den dag då ansökan om exportlicens inlämnas, tillämpas vid export som sker inom licensens giltighetstid och att ett korrektionsbelopp i så fall skall användas för exportbidraget. Enligt artikel 1 i kommissionens förordning nr 474/67/EEG om förutfastställelse av exportbidraget för ris och brutet ris(2), är korrektionsbeloppet lika med skillnaden mellan cif-priset och cif-priset vid terminsköp.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
I artikel 1 i förordning nr 474/67/EEG skall första och andra stycket ersättas med följande:
Under tiden mellan de veckovisa fastställelserna skall det bidragsbelopp som gäller vid förutfastställelse endast justeras om tillämpningen av ovannämnda bestämmelse medför att beloppet ändras med mer än 0,025 räkneenheter per 100 kg."
RÅDETS DIREKTIV av den 20 mars 1970 om tillnärmning av medlemsstaternas lagstiftning om åtgärder mot luftförorening genom avgaser från motorfordon (70/220/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: Förordningen av den 14 oktober 1968 med ändring i Straßenverkehrs-Zulassungs-Ordnung publicerades i Tyskland i Bundesgesetzblatt Del 1 den 18 oktober 1968. Denna förordning innehåller bestämmelser om åtgärder mot luftföroreningar från förbränningsmotorer i motorfordon. Bestämmelserna kommer att träda i kraft den 1 oktober 1970.
Varje medlemsstat som skall utfärda ett nationellt typgodkännande för en fordonstyp måste genom det nämnda meddelandet kunna förvissa sig om att fordonstypen genomgått de prov som krävs enligt detta direktiv. Därför bör varje medlemsstat underrätta övriga medlemsstater om sina resultat genom att sända dem en kopia av det meddelande som upprättats för varje motorfordonstyp som provats.
Artikel 1
Ingen medlemsstat får vägra att bevilja EEG-typgodkännande eller nationellt typgodkännande för ett fordon av skäl som hänför sig till luftförorening genom gaser från förbränningsmotorer med styrd tändning i fordonet - från och med den 1 oktober 1970, om fordonet uppfyller både kraven i bilaga 1, med undantag för kraven i punkt 3.2.1.1 och 3.2.2.1, och kraven i bilagorna 2, 4, 5 och 6,
1. När en ansökan kommer in från en tillverkare eller dennes representant skall de behöriga myndigheterna i den berörda medlemsstaten fylla i uppgifterna i meddelandet enligt bilaga 7. En kopia av meddelandet skall sändas till övriga medlemsstater och till sökanden. Andra medlemsstater som får en ansökan om nationellt typgodkännande för samma fordonstyp skall godta det nämnda dokumentet som bevis för att de föreskrivna proven har utförts.
Den medlemsstat som har beviljat ett typgodkännande skall vidta de åtgärder som krävs för att säkerställa att den underrättas om varje ändring i fråga om delar eller egenskaper som avses i punkt 1.1 i bilaga 1. De behöriga myndigheterna i medlemsstaten skall avgöra om nya prov måste utföras på den ändrade prototypen och om en ny rapport måste upprättas. Om dessa prov visar att kraven i detta direktiv inte uppfylls skall ändringen inte godkännas.
Artikel 6
Artikel 7
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande,
Råolja och petroleumprodukter är av allt större betydelse för gemenskapens försörjning med energi. Varje svårighet, även om den är tillfällig, som väsentligt begränsar leveranserna av dessa produkter, skulle kunna vålla allvarliga störningar i gemenskapens ekonomiska verksamhet. Gemenskapen bör därför kunna upphäva eller i vart fall minska de skadliga verkningar som skulle kunna uppstå i ett sådant fall.
En viss överensstämmelse mellan dessa befogenheter är nödvändig för att underlätta en samordning av de enskilda staternas åtgärder inom ramen för samråd på gemenskapsnivå.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Om svårigheter i försörjningen med råolja eller petroleumprodukter uppkommer i gemenskapen eller i en av medlemsstaterna skall kommissionen på begäran av en medlemsstat eller på eget initiativ snarast sammankalla en grupp av företrädare för medlemsstaterna, i vilken kommissionens företrädare skall vara ordförande.
Artikel 6
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag, och
Artikel 1
Artikel 2
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
Gemensamma krav för inre backspeglar har lagts fram genom rådets direktiv av den 1 mars 1971(4) och krav bör också utarbetas för passagerarutrymmets inredningsdetaljer, manöverorganens utformning, taket och ryggstöden och sätenas baksida. Ytterligare krav avseende inredning kommer att antas senare, särskilt i fråga om förankringspunkter för bilbälten och säten, huvudstöd, skydd för föraren mot styranordningen och identifikation av manöverorganen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
- taket eller det öppningsbara taket,
Artikel 3
- taket eller det öppningsbara taket,
Artikel 4
De ändringar som är nödvändiga för att anpassa kraven i bilagorna till den tekniska utvecklingen skall beslutas enligt det förfarande som föreskrivs i artikel 13 i rådets direktiv av den 6 februari 1970 om en anpassning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon.
2. Medlemsstaterna ska se till att till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
RÅDETS FÖRORDNING (EEG) nr 668/74 av den 28 mars 1974 om ändring av förordning (EEG) nr 922/72 om allmänna tillämpningsföreskrifter för stöd till silkesodling
med beaktande av rådets förordning (EEG) nr 845/72(1) av den 24 april 1972 om särskilda åtgärder för att främja silkesodling, särskilt artikel 2.4 i denna,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
RÅDETS DIREKTIV av den 17 december 1974 om utvidgande av tillämpningsområdet för direktiv nr 64/221/EEG om samordningen av särskilda åtgärder som gäller utländska medborgares rörlighet och bosättning och som är berättigade med hänsyn till allmän ordning, säkerhet eller hälsa till att även omfatta medborgare i en medlemsstat som begagnar sig av rätten att stanna kvar inom en annan medlemsstats territorium efter att ha verkat där som egna företagare (75/35/EEG)
med beaktande av Europaparlamentets yttrande (1),
Direktiv nr 64/221/EEG bör därför gälla för personer som omfattas av direktiv 75/34/EEG.
Direktiv nr 64/221/EEG skall gälla för medborgare i medlemsstaterna och deras familjemedlemmar som har rätt att stanna kvar inom en medlemsstats territorium i enlighet med direktiv nr 75/34/EEG
RÅDETS DIREKTIV av den 20 maj 1975 om tillnärmning av medlemsstaternas lagar och andra författningar beträffande aerosolbehållare (75/324/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: I vissa medlemsstater är det ett obligatoriskt krav att aerosolbehållare motsvarar vissa tekniska specifikationer. Sådana specifikationer varierar från medlemsstat till medlemsstat, vilket hindrar handeln inom gemenskapen.
De tekniska specifikationer som anges i bilagan till detta direktiv kommer inom kort att behöva anpassas till tekniska framsteg. För att underlätta att nödvändiga åtgärder genomförs på ett effektivt sätt skall former fastställas för ett nära samarbete mellan medlemsstaterna och kommissionen inom ramen för en kommitté för anpassning av direktivet om aerosolbehållare till teknisk utveckling.
Artikel 1
I detta direktiv avses med aerosolbehållare varje behållare som inte kan återanvändas, är tillverkad av metall, glas eller plast, innehåller gas som komprimerats, kondenserats eller lösts under tryck, med eller utan vätska, pasta eller pulver, och som är försedd med en utlösningsanordning för att spruta ut innehållet som en suspension av fasta eller flytande partiklar i gas, som lödder, pasta eller pulver eller i flytande tillstånd.
Artikel 4
1. En kommitté för anpassning av direktivet om aerosolbehållare till teknisk utveckling, nedan kallad "kommittén", inrättas härmed. Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
1. När det förfarande som anges i denna artikel skall tillämpas, skall ordföranden hänskjuta ärendet till kommittén, antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
b) Om förslaget inte har tillstyrkts av kommittén eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet åtgärder. Rådet skall fatta sitt beslut med kvalificerad majoritet.
1. Varje aerosolbehållare skall vara försedd med följande uppgifter i väl synlig, läslig och varaktig skrift som, om förpackningen är av liten volym (högst 150 ml), kan anbringas på en vidfäst etikett; denna bestämmelse gäller utöver krav i andra av gemenskapens direktiv, särskilt direktiven om farliga ämnen och beredningar: a) Namn och adress eller varumärke för den person som svarar för utsläppandet på marknaden av aerosolbehållaren.
d) De uppgifter som anges i punkt 2.2 i bilagan.
Artikel 9
1. Om någon medlemsstat uppmärksammar att en eller flera aerosolbehållare på goda grunder kan antas medföra fara för hälsa och säkerhet, trots att den eller de motsvarar kraven i detta direktiv, har denna stat rätt att provisoriskt förbjuda försäljning av dessa behållare inom sina nationsgränser eller förena försäljningen med särskilda villkor. Medlemsstaten skall omedelbart underrätta de andra medlemsstaterna och kommissionen om detta och ange skälen till sitt beslut.
Artikel 11
Artikel 12
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(1),
Under den tid då direktiven tillämpats har det framkommit att små förpackningar av betutsäde och utsäde av foderväxter utgör en handelsvara inom gemenskapen.
Vissa av ovannämnda direktiv innehåller bestämmelser om att likvärdighet hos utsäde som skördats i andra länder, särskilt i tredje land, fr.o.m. den 1 juli 1975 inte längre får beslutas nationellt av medlemsstaterna. Eftersom det inte har varit möjligt att utföra gemensam undersökning av utsäde av foder-, olje- och spånadsväxter i samtliga fall bör dock ovannämnda period förlängas för dessa utsäden för att undvika att nuvarande handelsförbindelser störs.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"G. EEG-småförpackningar: förpackningar med följande certifikatutsäden: - Monogermt frö eller tekniskt monogermfrö (precisionsfrö): högst 100 000 frögyttringar eller frön eller med en nettovikt om 2,5 kg, exklusive, i förekommande fall, pesticider i pulverform, pelleteringsmedel eller andra fasta tillsatser.
2. Medlemsstaterna skall kräva, förutom för EEG-småförpackningar, att förpackningar inte omplomberas, varken en eller flera gånger, annat än genom officiell plombering. Om förpackningar omplomberas, skall detta samt ansvarig myndighet och datum för omplombering anges på den etikett som krävs enligt artikel 11.1.
4. Det inledande avsnittet i artikel 11.1 skall ersättas med följande:
"b) anta bestämmelser om undantag från punkt 1 för småförpackningar med basutsäde om dessa är märkta med: "Endast godkänt för saluföring i . . . . . . (den berörda medlemsstaten)"."
RÅDETS FÖRORDNING (EEG) nr 2777/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för fjäderfäkött
med beaktande av kommissionens förslag,
För att den gemensamma marknaden för jordbruksprodukter skall kunna fungera och utvecklas måste den kompletteras av en gemensam jordbrukspolitik som framför allt innefattar gemensam organisation av marknaderna för olika jordbruksprodukter. En sådan organisation kan utformas på olika sätt beroende på vilket produkt det är fråga om.
För att uppnå detta syfte bör det i regel vara tillräckligt att i samband med import från tredje land införa importavgifter som bestäms med hänsyn till effekten på foderkostnaderna av den skillnad som råder mellan priserna på foderspannmål inom gemenskapen och på världsmarknaden, och till behovet att skydda gemenskapens förädlingsindustri.
Utöver det ovan beskrivna systemet bör möjligheter skapas att, när marknadssituationen så kräver, helt eller delvis förbjuda tillämpningen av aktiv förädling.
De utgifter som medlemsstaterna ådrar sig till följd av förpliktelser som uppstår vid tillämpningen av denna förordning skall finansieras av gemenskapen i enlighet med bestämmelserna i artikel 2 och 3 i rådets förordning (EEG) nr 729/70(2) av den 21 april 1970 om finansieringen av den gemensamma jordbrukspolitiken, ändrad genom förordning (EEG) nr 1566/72(3).
b) kycklingar: levande höns, ankor, gäss, kalkoner och pärlhöns med en högsta vikt på 185 gram.
2. produkter enligt punkt 1 b utom slaktade fjäderfä och ätbara slaktbiprodukter så kallade styckningsdelar av fjäderfä,
5. produkter enligt punkt 1 d och e,
Artikel 2
- Åtgärder för att underlätta registreringen av prisutvecklingen på marknaden.
- får antas för de produkter som anges i artikel 1.1 a, c, d, e och f.
Artikel 3
1. Importavgiften på slaktat fjäderfä skall bestå av följande delar: a) En del som motsvarar skillnaden mellan gemenskapens och världsmarknadens priser på den kvantitet fodersäd, differentierad med hänsyn till art av fjäderfä, som åtgår till att inom gemenskapen producera 1 kg slaktat fjäderfä.
Vid fastställande av de importavgifter som skall tillämpas från och med den 1 november, den 1 februari och den 1 maj, skall emellertid hänsyn tas till utvecklingen av världsmarknadspriserna på foderspannmål endast om ett nytt slusspris fastställs samtidigt.
- anta tillämpningsföreskrifter för denna artikel.
2. Trots bestämmelserna i punkt 1 skall importavgiften för de produkter som anges under Gemensamma tulltaxans nummer 02.03, 15.01 B och 16.02 B I och för vilka tullsatsen har bundits inom GATT, begränsas till det belopp som följer av denna bundenhet.
Om en betydande prisökning noteras på gemenskapsmarknaden och denna situation sannolikt kommer att bestå och därigenom stör eller hotar att störa marknaden, får nödvändiga åtgärder vidtas.
1. Slusspriserna skall fastställas på förhand för varje kvartal i enlighet med artikel 17.
Världsmarknadspriset på kvantiteten av foderspannmål skall fastställas kvartalsvis på basis av priserna på sådan spannmål under de sex månader som föregår det kvartal under vilket slusspriset fastställs.
4. För de produkter som anges i artikel 1.2 d skall slusspriserna härledas från slusspriset på slaktat fjäderfä på basis av de koefficienter som fastställts för sådana produkter i enlighet med artikel 5.3.
1. Om anbudspriset fritt gränsen för en produkt ligger under slusspriset, skall importavgiften för denna vara höjas med en tilläggsavgift som motsvarar skillnaden mellan slusspriset och anbudspriset fritt gränsen.
Om exporten från ett eller flera tredje länder sker till onormalt låga priser, lägre än de priser som gäller i andra tredje länder, skall ett andra anbudspris fritt gränsen fastställas för export från dessa länder.
Artikel 9
Exportbidraget skall beviljas på ansökan av berörd part.
Exportbidrag skall fastställas med jämna mellanrum i enlighet med förfarandet i artikel 17. Vid behov får kommissionen, på begäran av en medlemsstat eller på eget initiativ, ändra exportbidragen under mellanperioderna.
I den mån det är nödvändigt för att den gemensamma organisation av marknaden för fjäderfäkött skall fungera väl, får rådet, på förslag av kommissionen, med kvalificerad majoritet helt eller delvis förbjuda tillämpningen av bestämmelserna för aktiv förädling för produkter enligt artikel 1.1 som skall användas till framställningen av de produkter som anges i den punkten.
2. Såvida inte annat föreskrivs i denna förordning eller rådet, på förslag av kommissionen, med kvalificerad majoritet fattar beslut om undantag från denna förordning, skall följande vara förbjudet:
Artikel 12
2. Om den situation som avses i punkt 1 uppstår skall kommissionen, på begäran av en medlemsstat eller på eget initiativ, fatta beslut om nödvändiga åtgärder. Medlemsstaterna skall underrättas om beslutet som skall gälla med omedelbar verkan. Om kommissionen mottar en begäran från en medlemsstat, skall den fatta beslut om denna begäran inom 24 timmar efter det att den mottagits.
De produkter som anges i artikel 1.1 och som framställs av eller utvinns ur produkter som inte är angivna i artikel 9.2 och 10.1 i fördraget skall inte få omsättas fritt inom gemenskapen.
Artikel 15
1. Härmed inrättas en förvaltningskommitté för fjäderfäkött och ägg (nedan kallad "kommittén"). Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
1. När förfarandet som föreskrivs i denna artikel skall tillämpas, skall ordföranden hänskjuta ärendet till kommittén, antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
Rådet får inom en månad fatta ett annat beslut med kvalificerad majoritet.
Artikel 19
Denna förordning skall tillämpas så att hänsyn tas samtidigt och på lämpligt sätt till de mål som fastställs i artiklarna 39 och 110 i fördraget.
Artikel 22
Hänvisningar till artiklar i den upphävda förordningen skall läsas enligt den jämförelsetabell som finns i bilagan.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Europaparlamentets yttrande(1),
Dessa krav skiljer sig åt från en medlemsstat till en annan. Det är därför nödvändigt att alla medlemsstater antar samma krav, antingen som tillägg till eller i stället för sina nuvarande regler, för att därmed för alla fordonstyper medge det förfarande för EEG-typgodkännande som behandlats i rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(3).
Artikel 1
Ingen medlemsstat får vägra att bevilja EEG-typgodkännande eller nationellt typgodkännande för ett fordon av skäl som hänför sig till de föreskrivna skyltarna och märkningarna eller deras placering och fastsättningsmetod om de uppfyller kraven i bilagan.
Artikel 4
2. Efter anmälan av detta direktiv skall medlemsstaterna underrätta kommissionen om alla förslag till lagar och andra författningar som de avser att anta inom det område som omfattas av detta direktiv; underrättelsen skall lämnas i så god tid att kommissionen hinner lämna synpunkter på förslaget.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(1),
Kontroll av badvatten är nödvändig för att inom ramen för den gemensamma marknaden uppnå gemenskapens mål vad avser en förbättring av levnadsvillkoren, en harmonisk utveckling av ekonomiska verksamheter inom gemenskapen som helhet och en fortgående och balanserad tillväxt.
För att uppnå dessa kvalitetsmål måste medlemsstaterna fastställa gränsvärden enligt vissa parametrar. Badvatten måste överensstämma med dessa värden inom tio år efter anmälan av detta direktiv.
Den tekniska utvecklingen gör det nödvändigt med en snabb anpassning av de tekniska krav som fastställs i bilagan. För att underlätta beslut om de åtgärder som krävs för detta ändamål, bör ett förfarande fastställas genom vilket ett nära samarbete upprättas mellan medlemsstaterna och kommissionen inom en kommitté för anpassning till den tekniska utvecklingen.
a) "badvatten": allt rinnande eller stillastående sötvatten och havsvatten, i vilket - badning är uttryckligen tillåten av de behöriga myndigheterna i varje medlemsstat, eller
c) "badsäsong": den period under vilken ett stort antal badare kan förutses med hänsyn till lokalt bruk, inbegripet eventuella lokala regler för badning och väderleksförhållanden.
Artikel 3
Kommissionen får delta i dessa överläggningar.
och om, i fråga om de 5, 10 eller 20 % av proven som inte överensstämmer med värdena
Artikel 7
b) om badvatten berikas på naturlig väg med vissa ämnen och detta orsakar avvikelse från de värden som föreskrivs i bilagan.
Om en medlemsstat åsidosätter bestämmelserna i detta direktiv skall den omedelbart meddela kommissionen detta med uppgift om skälen och den förväntade tidsperioden.
- de G- och I-parametervärden som anges i bilagan.
Artikel 11
c) Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Kommissionen kan offentliggöra den erhållna informationen efter det att den berörda medlemsstaten har gett sitt tillstånd.
RÅDETS DIREKTIV av den 27 juli 1976 om tillnärmning av medlemsstaternas lagstiftning om alkoholmätare och alkoholaerometrar (76/765/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: Definition, konstruktion och metoder för godkännande och provning av alkoholmätare och alkoholaerometrar är i medlemsstaterna underkastade tvingande bestämmelser som skiljer sig mellan medlemsstaterna och därmed utgör hinder för rörligheten av och handeln med dessa mätdon inom gemenskapen. Dessa bestämmelser måste därför närmas till varandra.
I sin resolution av den 17 december 1973(4) om industripolitik uppmanade rådet kommissionen att före den 1 december 1974 till rådet lämna ett förslag till ett direktiv om alkoholmätning och alkoholmätare.
Detta direktiv fastställer egenskaper hos alkoholmätare och alkoholaerometrar som används för att bestämma alkoholhalten i blandningar av vatten och etanol.
Ingen medlemsstat får begränsa, vägra eller förbjuda att någon alkoholmätare eller alkoholaerometer släpps ut på marknaden eller tas i drift, under åberopande av dess metrologiska egenskaper, om den försetts med märkning för EEG-typgodkännande eller första EEG-verifikation.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
RÅDETS DIREKTIV av den 16 december 1976 om minimikrav på utbildning av vissa förare av vägfordon (76/914/EEG)
med beaktande av rådets förordning (EEG) nr 543/69 av den 25 mars 1969 om harmonisering av viss social lagstiftning rörande transporter på väg(), senast ändrad genom förordning (EEG) nr 515/72(), och särskilt artikel 5.1 b andra strecksatsen och artikel 2 c i denna,
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Kursinnehåll och uppläggning i fråga om den yrkesutbildning som avses i punkt 1 skall fastställas av medlemsstaten. Att sådan utbildning har genomgåtts skall styrkas genom examen eller kunskapskontroll som ombesörjs av staten eller av de organ som staten har utsett att utföra kontrollen under direkt överinseende av staten.
1. Det intyg om yrkeskompetens som avses i andra strecksatsen i artikel 5.1 b och artikel 5.2 c i förordning (EEG) nr 543/69 skall utfärdas till de personer som uppfyller de villkor som föreskrivs i artikel 1 i detta direktiv av den stat eller av de organ som staten utsett att ombesörja utfärdandet under direkt överinseende av staten.
1. Efter samråd med kommissionen skall medlemsstaterna inom två år efter anmälan av detta direktiv genomföra de åtgärder som är nödvändiga för att följa direktivet.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 113 i detta,
Artikel 1
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 54.3 g i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
Inom gemenskapen måste ett aktiebolags bolagsordning eller stiftelseurkund utformas på ett sådant sätt att varje intressent ur dessa handlingar kan inhämta grundläggande uppgifter om bolaget, däribland en detaljerad redovisning av kapitalets sammansättning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE
- I Danmark: aktieselskabet.
Med "förvaltningsbolag med rörligt kapital" avses i detta direktiv endast bolag - som uteslutande har till föremål för sin verksamhet att placera sina medel i olika värdepapper, fastigheter eller andra tillgångar med enda syfte att sprida investeringsriskerna och fördela resultatet av kapitalförvaltningen mellan aktieägarna,
Artikel 2
c) - om bolaget inte har något "auktoriserat" kapital, det tecknade kapitalets storlek;
e) tiden för bolagets bestånd om inte denna tid är obestämd.
b) de tecknade aktiernas nominella belopp och, minst en gång om året, deras antal;
e) om det finns aktier av olika slag, uppgifter enligt b, c och d för varje aktieslag med uppgift om de rättigheter som är förenade med varje aktieslag;
h) det nominella värdet av de aktier eller, i avsaknad av sådant värde, det antal aktier som ges ut mot tillskott av annan egendom än pengar (apportegendom) samt beskrivning av denna egendom och namnet på den som tillskjuter egendomen;
k) särskilda förmåner som vid bolagsbildningen eller före tillståndet att börja verksamheten har tillerkänts någon som har deltagit i bolagsbildningen eller i åtgärder som har lett fram till tillståndet.
2. Punkt 1 tillämpas inte på förbindelser med anledning av avtal som bolaget har ingått på villkor att det får tillstånd att börja sin verksamhet.
2. Om enligt lagstiftningen i en medlemsstat ett bolag i fall som avses i punkt 1 kan upplösas genom förordnande av rätten, får behörig domstol ge bolaget den frist som detta behöver för att vidta rättelse.
1. Medlemsstaternas lagstiftning skall föreskriva att ett kapital på minst 25 000 europeiska beräkningsenheter måste tecknas för att bolaget skall få bildas eller få tillstånd att börja sin verksamhet.
Artikel 7
1. Aktierna får inte ges ut mot vederlag som understiger det nominella beloppet eller, om sådant saknas, det bokförda parivärdet.
1. Aktier som ges ut mot vederlag måste då bolaget bildas eller får tillstånd att börja sin verksamhet vara betalda till minst 25 procent av det nominella beloppet eller, om sådant saknas, av det bokförda parivärdet.
1. En eller flera av bolaget oberoende sakkunniga, som utses eller godkänns av en förvaltningsmyndighet eller en domstol, skall avge ett utlåtande om apportegendomen innan bolaget bildas eller får tillstånd att börja sin verksamhet. Beroende på varje medlemsstats lagstiftning kan de sakkunniga vara fysiska eller juridiska personer eller bolag.
4. En medlemsstat får underlåta att tillämpa denna artikel om samtliga aktier till 90 procent av sitt nominella värde eller, i avsaknad av sådant värde, av sitt bokförda parivärde utges mot apportegendom från ett eller flera bolag och följande villkor är uppfyllda: a) de i artikel 3 i avsedda personerna eller bolagen med anknytning till det bolag som tar emot apportegendomen har avstått från att kräva sakkunnigutlåtande;
d) de bolag som lämnar apportegendomen förklarar, att de med belopp som motsvarar det vid c angivna värdet åtar sig ansvar för skulder som kan uppkomma för det mottagande bolaget från det att detta bolag har gett ut aktierna mot apportegendom till dess att ett år har förflutit från bolagets offentliggörande av årsredovisningen för det räkenskapsår under vilket apportegendomen lämnades; överlåtelse av aktierna får inte ske under denna tid;
Artikel 11
2. Punkt 1 tillämpas inte i fråga om förvärv som sker inom ramen för bolagets löpande verksamhet, på begäran eller under kontroll av en förvaltningsmyndighet eller en domstol eller på en fondbörs.
Artikel 13
Artiklarna 2-13 skall inte inverka på medlemsstaternas föreskrifter om kompetens och tillvägagångssätt vid ändring av en bolagsordning eller en stiftelseurkund.
b) Det vid a angivna tecknade beloppet skall minskas med sådan icke inbetald del därav som inte redovisas på balansräkningens aktivsida.
2. Om lagstiftningen i en medlemsstat tillåter förskottsutdelning av vinst skall minst följande villkor iakttas: a) ett delårsbokslut skall upprättas som visar att tillräckliga medel finns tillgängliga för utdelningen;
4. Lagstiftningen i en medlemsstat får föreskriva undantag från punkt 1 a i fråga om förvaltningsbolag med fast kapital.
I den omfattning den nu angivna möjligheten används i medlemsstaternas lagstiftning a) skall denna ålägga bolagen ifråga att föra in ordet "förvaltningsbolag" i alla dokument som anges i artikel 4 i direktiv 68/151/EEG;
Artikel 16
1. Vid betydande förlust av det tecknade kapitalet skall kallelse inom den tid som anges i medlemsstaternas lagstiftning ske till en bolagstämma, som skall pröva om bolaget skall upplösas eller om andra åtgärder skall vidtas.
1. Ett bolag får inte teckna sina egna aktier.
Lagstiftningen i en medlemsstat får dock bestämma att den skall befrias från betalningsansvar som kan visa att han inte har försummat något.
b) Det nominella värdet eller, om sådant värde saknas, det bokförda parivärdet hos de förvärvade aktierna inräknat de aktier som bolaget tidigare har förvärvat och fortfarande innehar samt de aktier som har förvärvats av någon som handlat i eget namn men för bolagets räkning, får inte överstiga tio procent av det tecknade kapitalet.
2. Lagstiftningen i en medlemsstat får medge undantag från punkt 1 a första meningen, om ett förvärv av egna aktier är nödvändigt för att bolaget skall undgå en betydande och nära förestående skada. I ett sådant fall skall styrelsen eller direktionen informera den närmast följande bolagsstämman om grunden för förvärvet och syftet med detta, om de förvärvade aktiernas antal och nominella värde eller, i avsaknad av sådant värde, bokförda parivärde, om den andel av det tecknade kapitalet som de förvärvade aktierna utgör samt om vederlaget för aktierna.
1. Medlemsstaterna behöver inte tillämpa artikel 19 på: a) aktier som förvärvas för att genomföra ett beslut om nedsättning av kapitalet eller i fall som avses i artikel 39;
d) aktier som förvärvas på grund av en lagstadgad skyldighet eller till följd av ett rättsligt avgörande till skydd för en aktieägarminoritet, särskilt vid fusion, ändring av föremålet för bolagets verksamhet eller av bolagets form, byte av säte till utlandet eller införandet av begränsningar i rätten att överlåta aktier;
g) helt betalda aktier som förvärvas vid en exekutiv aktion som äger rum för att infria en fordran som bolaget har mot en aktieägare;
3. Om aktierna inte avyttras inom den tid som anges i punkt 2 skall de förklaras ogiltiga. Lagstiftningen i en medlemsstat kan bestämma att ogiltigförklaringen skall åtföljas av en motsvarande nedsättning av det tecknade kapitalet. En sådan nedsättning skall föreskrivas i den mån förvärvet av de aktier som skall förklaras ogiltiga har medfört att nettotillgångarna kommit att understiga det belopp som anges i artikel 15.1 a.
Artikel 22
2. Om lagstiftningen i en medlemsstat tillåter ett bolag att förvärva egna aktier, direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall lagstiftningen kräva att förvaltningsberättelsen innehåller minst följande uppgifter: a) skälen för de förvärv som har skett under räkenskapsåret;
d) antal och nominellt värde eller, i avsaknad av sådant värde, bokfört parivärde beträffande samtliga aktier som har förvärvats och som innehas av bolaget samt den andel av det tecknade kapitalet som dessa aktier utgör.
2. Punkt 1 tillämpas inte på åtgärder som utgör led i en banks eller något annat finansinstituts löpande verksamhet eller som vidtas i syfte att aktier skall förvärvas av eller till förmån för de anställda i bolaget eller ett detta närstående bolag. Sådana åtgärder får dock inte leda till att nettotillgångarna understiger det belopp som anges i artikel 15.1 a.
1. Om ett bolag direkt eller genom någon som handlar i eget namn men för bolagets räkning tar emot egna aktier som säkerhet, jämställs detta med förvärv som avses i artiklarna 19 och 20.1 samt artiklarna 22 och 23.
1. Alla kapitalökningar skall beslutas av bolagsstämman. Ett sådant beslut, liksom genomförandet av kapitalökningen, skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
4. Denna artikel tillämpas vid emission av alla värdepapper som kan bytas ut mot aktier eller som är förenade med teckningsrätt till aktier, men inte vid själva utbytet av värdepapperen eller vid utnyttjandet av teckningsrätten.
Artikel 27
4. Medlemsstaterna behöver inte tillämpa punkt 2 när alla aktier som emitteras som ett led i ökningen av det tecknade kapitalet ges ut mot apportegendom från ett eller flera bolag, om alla aktieägare i det bolag som tar emot apportegendomen har avstått från sakkunnigutlåtande samt villkoren i artikel 10.4b-f är uppfyllda.
Artikel 29
b) får - om i ett bolag med aktier av olika slag i fråga om rösträtt eller rätt till utdelning enligt artikel 15 eller vid utskiftning i samband med likvidation, det tecknade kapitalet ökas genom att nya aktier av endast ett av dessa aktieslag ges ut - tillåta att ägarna till aktier av annat slag får utöva sin företrädesrätt att teckna nya aktier först efter ägarna till aktier av det slag som emissionen avser.
5. Lagstiftningen i en medlemsstat får bestämma att bolagsordningen, stiftelseurkunden eller bolagsstämman, den senare med iakttagande av bestämmelserna i punkt 4 angående beslutförhet, majoritet och offentliggörande, kan bemyndiga det bolagsorgan att begränsa eller upphäva företrädesrätten som har rätt att besluta om ökning av aktiekapitalet inom gränserna för det "auktoriserade" kapitalet. Ett sådant bemyndigande får inte gälla för längre tid än ett bemyndigande enligt artikel 25.2.
Artikel 30
Artikel 32
3. Denna artikel tillämpas även när nedsättningen av det tecknade kapitalet sker genom att bolaget helt eller delvis avstår från betalning av aktieägarnas insatser.
2. I de fall som avses i punkt 1 skall medlemsstaternas lagstiftning minst föreskriva de åtgärder som behövs för att belopp som härrör från nedsättningen av det tecknade kapitalet inte skall kunna användas för utbetalningar till aktieägarna eller för att befria dessa från skyldigheten att betala sina insatser.
Artikel 35
c) De aktieägare som har fått sina aktier inlösta har kvar sina rättigheter i bolaget med undantag för rätten att återfå insatserna och rätten att delta i en första vinstutdelning avseende icke inlösta aktier.
a) Tvångsindragningen skall föreskrivas eller tillåtas i bolagsordningen eller stiftelseurkunden innan teckning sker av de aktier som skall dras in. b) I det fallet att tvångsindragningen endast tillåts i bolagsordningen eller stiftelseurkunden skall den beslutas av bolagstämman, om inte samtliga berörda aktieägare har godkänt indragningen.
e) Beslutet om tvångsindragning skall offentliggöras enligt varje lands lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
1. Om det tecknade kapitalet sätts ned genom indragning av aktier som bolaget har förvärvat direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall bolagsstämman alltid besluta om indragningen.
Artikel 38
Om lagstiftningen i en medlemsstat tillåter bolagen att ge ut aktier som kan återköpas, skall lagstiftningen för återköp av aktierna minst kräva att följande villkor är uppfyllda: a) återköpet skall tillåtas i bolagsordningen eller stiftelseurkunden innan teckning sker av de aktier som kan återköpas;
d) återköpet får endast ske med medel som kan delas ut enligt artikel 15.1 eller med intäkter från en nyemission som sker i och för återköpet;
g) om det har beslutats att en överkurs skall betalas till aktieägarna med anledning av återköpet, får överkursen endast erläggas med medel som får delas ut enligt artikel 15.1 eller med medel ur en reserv, annan än den som avses i e, som inte får delas ut till aktieägarna i annat fall än då det tecknade kapitalet sätts ned; denna reserv får endast användas för att öka det tecknade kapitalet genom överföring av reserver, för att täcka kostnader som avses i artikel 3 j eller emissionskostnader för aktier eller obligationer eller för att betala en överkurs till innehavare av aktier eller obligationer som skall återköpas;
1. Medlemsstaternas lagstiftning skall föreskriva att de beslut som avses i artikel 29.4 och 5 samt artiklarna 30, 31, 35 och 38 skall kräva minst en majoritet som inte får understiga två tredjedelar av de röster som är förenade med de företrädda värdepapperen eller det företrädda tecknade kapitalet.
1. Medlemsstaterna får frångå artikel 9.1, artikel 19.1 a första ledet och b samt artiklarna 25, 26 och 29 i den mån det behövs för att bestämmelser skall kunna antas eller tillämpas som har till ändamål att underlätta för anställda och andra i den nationella lagstiftningen angivna personkategorier att få del i företagens kapital.
För att detta direktiv skall kunna genomföras måste medlemsstaternas lagstiftning behandla de aktieägare lika som befinner sig i samma ställning.
RÅDETS DIREKTIV av den 25 juli 1977 om renrasiga avelsdjur av nötkreatur (77/504/EEG)
med beaktande av Europaparlamentets yttrande(1),
De flesta medlemsstater har hittills strävat efter att som ett led i den nationella avelspolitiken främja produktionen av husdjur av ett begränsat antal raser som uppfyller särskilda avelsmässiga normer. Raser och normer skiljer sig åt från en medlemsstat till en annan och dessa skillnader hindrar handeln inom gemenskapen.
Inom vissa tekniska områden bör åtgärder för genomförande vidtas. För att besluta om sådana åtgärder bör ett förfarande fastställas som leder till ett nära samarbete mellan medlemsstaterna och kommissionen inom Ständiga kommittén för husdjursavel. Till dess att beslut fattas om dessa åtgärder för genomförande skall nu gällande bestämmelser på de områden det är fråga om förbli oförändrade.
Artikel 1
- där renrasiga avelsdjur av en viss ras av nötkreatur är införda eller registrerade med uppgifter om deras härstamning.
- Handel med sperma och embryon från renrasiga avelsdjur av nötkreatur inom gemenskapen.
- Handel inom gemenskapen med tjurar som används för artificiell insemination, om inte annat följer av artikel 3.
Till dess att sådana bestämmelser träder i kraft skall godkännande av renrasiga djur av nötkreatur för avelsändamål, godkännande av tjurar för artificiell insemination samt användning av sperma och embryon lyda under nationell rätt, förutsatt att denna inte är mer restriktiv än den lagstiftning som är tillämplig på renrasiga avelsdjur av nötkreatur, sperma och embryon i den medlemsstat som är destinationsland.
Artikel 5
1. Följande skall bestämmas enligt det förfarande som fastställs i artikel 8:
- Villkor för införande i stamböcker.
b) skall godkännandet av avelsorganisationer eller avelsföreningar även fortsättningsvis regleras av de föreskrifter som för närvarande gäller i varje medlemsstat,
Till dess att gemenskapsregler införs på området får de villkor som gäller import av renrasiga avelsdjur av nötkreatur från icke-medlemsländer inte vara mer gynnsamma än de som gäller för handeln inom gemenskapen.
1. När det förfarande som fastställs i denna artikel skall tillämpas skall ordföranden utan dröjsmål hänskjuta ärendet till Ständiga kommittén för husdjursavel (i det följande kallad "kommittén"), upprättad genom rådets beslut 77/505/EEG, antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
4. Kommissionen skall själv anta förslaget och genomföra det omedelbart om det har tillstyrkts av kommittén. Om förslaget inte har tillstyrkts av kommittén eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 1979 och skall genast underrätta kommissionen om detta.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning nr 162/66/EEG av den 27 oktober 1966 om handeln med oljor och fetter mellan gemenskapen och Grekland(3),
Kontantbidraget beviljas endast för vissa kvaliteter av olivolja och vissa presentationsformer av oljan. För att förhindra vissa uppgörelser som inte svarar mot sedvanliga exportmönster, bör det föreskrivas att rätten att importera med befrielse från avgift bör medges endast när exporten omfattar varor och presentationsformer för vilka ett kontantbidrag verkligen kan beviljas.
Artikel 1
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av följande: Mot bakgrund av den tekniska och vetenskapliga kunskapsutvecklingen bör bilagorna 1, 2 och 3 till ovannämnda direktiv ändras av de skäl som anges nedan.
I syfte att höja det genetiska värdet på utsäde bör bestämmelser om standarder för sortrenhet som måste uppfyllas av grödan antas för ytterligare ett antal arter.
I den situation som för närvarande råder har det inte varit möjligt att uppnå fullständig harmonisering inom gemenskapen av de villkor som gäller för förekomst a
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: Den internationella standardiseringsorganisationen ISO har nu antagit två internationella standarder om ett världstäckande klassificeringssystem, som gör det möjligt att identifiera tillverkaren av ett fordon(3) och även fordonet(4). Det är därför lämpligt att införa i direktiv 76/114/EEG detta system för identifiering av tillverkare, och samtidigt anpassa kraven om identifiering av fordon i direktivet med ISO-standarden.
Artikel 1
1. Från den 1 oktober 1978 får ingen medlemsstat, av skäl som hänför sig till föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt, - vägra att bevilja EEG-typgodkännande för en fordonstyp, vägra att utfärda det dokument som anges i artikel 10.1 sista strecksatsen i direktiv 70/156/EEG, eller vägra att bevilja nationellt typgodkännande, eller
2. Från den 1 oktober 1981 gäller följande: - Medlemsstaterna får inte längre utfärda den handling som anges i artikel 10.1 sista strecksatsen i direktiv 70/156/EEG för en typ av fordon för vilka föreskrivna skyltar och märkningar samt deras placering och fastsättning inte överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av Europaparlamentets yttrande(3), och
Det bör fastställas att utgifter i samband med interventionsåtgärder för vilka ett belopp per enhet bestäms inom ramen för en gemensam organisation av marknaderna helt skall täckas av gemenskapsmedel.
De allmänna bestämmelserna för gemenskapsfinansiering av interventioner bör samlas i en enda förordning. Rådets förordning (EEG) nr 2824/72 av den 28 december 1972 om allmänna bestämmelser för finansiering av interventioner genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket(4) bör därför upphävas.
De åtgärder som förtecknas i bilagan motsvarar begreppet intervention för stabilisering av jordbruksmarknaderna enligt artikel 3.1 i förordning (EEG) nr 729/70.
Artikel 3
2. För övriga interventionsåtgärder som anges i artikel 3 skall finansieringen vara lika med utgifterna med avdrag för eventuella intäkter som interventionsåtgärden medför.
Artikel 6
Om de aktuella produkterna till följd av lagringen minskar i värde, skall den finansiella effekten av denna värdeminskning fastställas och bokföras när produkten övergår i intervention. För detta ändamål skall värdeminskningskoefficienterna och de priser för vilka de skall tillämpas bestämmas enligt förfarandet i artikel 26 i rådets förordning (EEG) nr 2727/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för spannmål(14), senast ändrad genom förordning (EEG) nr 1254/78(15), eller motsvarande artikel i övriga förordningar om den gemensamma organisationen av jordbruksmarknaderna, och vid behov efter granskning i EUGFJ-kommittén.
Om det beräknade priset för en given produkt när interventionen upphör är väsentligt lägre än värdet av de lager som skall överföras, värderade enligt det förfarande som anges i första stycket, får dock beslut fattas om att ersätta det inköpspris som interventionsorganen betalat med ett annat pris. Detta pris skall fastställas enligt förfarandet i artikel 13 i förordning (EEG) nr 729/70, vid behov efter granskning i den berörda förvaltningskommittén. Det får inte vara lägre än de genomsnittliga inköpspriserna och de priser som erhålls vid avyttring av interventionslager.
Artikel 10
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av rådets direktiv 71/320/EEG av den 26 juli 1971 om tillnärmning av medlemsstaternas lagstiftning om bromsutrustning på vissa kategorier av motorfordon och släpvagnar till dessa fordon(3), i dess lydelse enligt kommissionens direktiv 75/524/EEG(4), och med beaktande av följande:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. I väntan på att särskilda bestämmelser angående låsningsfria bromssystem skall träda i kraft, skall fordon i kategorierna M1, M2, M3, N1, N2, N3, O3 och O4 som är utrustade med sådana system underkastas bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
- vägra att bevilja EEG-typgodkännande eller att utfärda det exemplar av det intyg som anges i sista strecksatsen i artikel 10.1 i direktiv 70/156/EEG eller att bevilja ett nationellt typgodkännande med avseende på en fordonstyp, eller
2. Från den 1 oktober 1980 skall medlemsstaterna
3. Från den 1 oktober 1981 får medlemsstaterna förbjuda ibruktagande av fordon vars bromsutrustning inte överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
Artikel 3
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
För att säkerställa att den olja som anbudet gäller och den olja som tilldelats är identiska, bör det vara möjligt att ta ytterligare ett prov innan det tilldelade partiet plomberas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"3. Under perioden från och med den 1 januari till och med 31 december 1979 skall minimipriset vara exklusive skatt och hänföra sig till 100 kg olivolja som levereras fritt lager, antingen i köparens egna fat och lastad på ett fordon som tillhandahållits av honom, eller i köparens tankfordon."
"Artikel 10Interventionsorganet skall genast meddela varje anbudsgivare med rekommenderat brev med mottagningsbevis om resultatet av hans deltagande i anbudsförfarandet."
1. Köparen skall, innan han avhämtar oljan, betala det preliminära försäljningspriset till interventionsorganet. Detta skall beräknas genom att multiplicera den kvantitet som enligt uppgift fanns i partiet med det pris som erbjudits för partiet.
8. Artikel 21 andra stycket skall utgå.
RÅDETS ELFTE DIREKTIV av den 26 mars 1980 om harmonisering av medlemsstaternas lagstiftning om omsättningsskatt - uteslutning av de franska utomeuropeiska departementen från tillämpningsområdet för direktiv 77/388/EEG (80/368/EEG)
med beaktande av kommissionens förslag, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
de utomeuropeiska departementen."
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Enligt kommissionens förordning (EEG) nr 797/80 av den 31 mars 1980 om justering av förutfastställda exportavgifter och exportbidrag för socker() skall exportbidragen höjas och exportavgifterna sänkas i fråga om exportlicenser som utfärdats före den 1 juli 1980 men som utnyttjas först efter detta datum.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. I punkt 2 skall följande läggas till som ett tredje stycke:
Denna förordning träder i kraft den 1 juli 1980.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(2),
Av trafiksäkerhetsskäl bör hädanefter montering av bilbälten och fasthållningsanordningar som överensstämmer med direktiv 77/541/EEG krävas i fordon i vissa M- och N-kategorier, och monteringen av dessa tillåtas och främjas i fordon i de övriga M- och N-kategorierna genom en utvidgning av räckvidden för detta direktiv. En sådan utvidgning har möjliggjorts av den tekniska utvecklingen i fråga om konstruktion av motorfordon.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. I bilaga 1: a) Avsnitt 3.1 skall ersättas med följande:
I de fall där andra fordon som omfattas av artikel 9 är utrustade med bilbälten eller fasthållningsanordningar skall dessa uppfylla alla krav i detta direktiv med undantag av avsnitten 3.1.1-3.1.3."
3.1.1.2 För passagerarsätet i fordon i kategori M2 anses höftbälten, med eller utan upprullningsdon, som tillräckliga om vindrutan befinner sig utanför den referenszon som definieras i bilaga 2 till direktiv 74/60/EEG.
"3.1.3 På bakre sittplatser i fordon i kategori M1, höftbälten eller trepunktsbälten antingen de är försedda med upprullningsdon eller inte."
Artikel 2
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 och 235 i detta,
med beaktande av följande: Artikel 11.2 i rådets direktiv 79/869/EEG av den 9 oktober 1979 om mätmetoder samt provtagnings- och analysfrekvenser avseende ytvatten för dricksvattenframställning i medlemsstaterna(2) bör ändras av hänsyn till Greklands anslutning till Europeiska gemenskaperna.
Artikel 1
Detta direktiv träder i kraft den 1 januari 1981.
RÅDETS FÖRORDNING (EEG) nr 654/81 av den 10 mars 1981 om ändring av rådets förordning (EEG) nr 3179/78 om Europeiska ekonomiska gemenskapens antagande av konventionen om framtida multilateralt samarbete om fisket i Nordvästatlanten
med beaktande av kommissionens förslag,
Den 7 juni 1979 antog Nordvästatlantiska fiskeriorganisationens allmänna råd, i enlighet med artikel 20 punkt 2 i den konventionen, med ikraftträdande den 1 januari 1980 sådana ändringar i bilaga 3 till konventionen om framtida multilateralt samarbete om fisket i Nordvästatlanten som rör avgränsningen mellan de statistiska delområdena i farvattnen mellan Grönlands västkust och Kanadas kust.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
med beaktande av kommissionens förslag (),
med beaktande av följande: Genom förordning nr 79/65/EEG (), senast ändrad genom förordning (EEG) nr 2910/73 () inrättade rådet ett informationssystem för jordbruksföretagens redovisningsuppgifter för att belysa inkomstförhållanden och andra ekonomiska förhållanden i jordbruksföretag i Europeiska ekonomiska gemenskapen.
Alla rapporterande företag som undersöks i medlemsstaterna för registrering av inkomster i jordbruket som underlag för jordbrukspolitiken bör tillhöra gemenskapens informationssystem och antalet rapporterande företag bör därför ökas. Detta antal bör kunna variera inom vissa gränser och beroende på utvecklingen inom jordbruket och kraven på uppgifter från den gemensamma jordbrukspolitiken.
Informationssystemets områden skall i största möjliga mån vara identiska med dem som används för att redovisa andra regionala uppgifter som är väsentliga för att skapa riktlinjer för den gemensamma jordbrukspolitiken. I detta avseende bör bilagan till förordning nr 79/65/EEG ändras.
"b) " () EGT nr L 148, 5.6.1978, s. 1."
1. Det undersökningsområde som avses i artikel 1.2 a skall omfatta de jordbruksföretag som är av en storlek som i ekonomiskt avseende är lika med eller större än det tröskelvärde, uttryckt i europeiska storleksenheter (ESE) som definieras genom beslut 78/463/EEG.
b) drivas av en jordbrukare som vill och kan sköta redovisningen för jordbruket och är beredd att ställa redovisningsuppgifter från sitt företag till kommissionens förfogande,
4. Tillämpningsföreskrifter till denna artikel, särskilt tröskelvärdet för företagens ekonomiska storlek och antalet rapporterande företag per område, skall fastställas enligt förfarandet i artikel 19."
1. Varje medlemsstat skall före den 1 februari 1982 inrätta en nationell kommitté för informationssystemet, nedan kallad "den nationella kommittén".
b) rapporten om tillämpningen av planen för val av rapporterande företag.
4. Medlemsstater som har flera områden får för varje område under sin jurisdiktion upprätta en regional kommitté för informationssystemet; nedan kallad "den regionala kommittén".
4) Artikel 6 skall ersättas med följande:
a) att underrätta den nationella kommittén, de regionala kommittéerna och bokföringsbyråerna om de gällande tillämpningsföreskrifterna och att säkerställa att dessa föreskrifter tillämpas korrekt,
P rapporten om genomförandet av planen för val av rapporterande företag,
P förteckningen över bokföringsbyråer som vill och kan upprätta företagsredovisningar, enligt de avtalsvillkor som anges i artiklarna 9 och 14, d) att sammanställa de företagsredovisningar som bokföringsbyråerna översänt och med hjälp av ett gemensamt kontrollprogram kontrollera att de är korrekt ifyllda,
2. Tillämpningsföreskrifterna till denna artikel skall utarbetas enligt förfarandet i artikel 19."
"1. Den nationella kommittén, de regionala kommittéerna, samordningsorganet och bokföringsbyråerna skall vara skyldiga att, inom sina respektive ansvarsområden, ge kommissionen alla uppgifter som den begär av dem om hur de utför sina arbetsuppgifter vid tillämpningen av denna förordning.
med beaktande av kommissionens förslag,
Förordning (EEG) nr 1108/70 (), i dess lydelse enligt förordning nr 1384/79 () skall ändras på så sätt att Greklands järnvägsnät tas in i bilagan till sistnämnda förordning.
Följande tillägg skall göras till förteckningen i bilaga 2 till förordning (EEG) nr 1108/70 under punkt "A.1.JÄRNVÄG - Huvudnät" efter rubriken "Förbundsrepubliken Tyskland":
Artikel 2
med beaktande av rådets direktiv 66/401/EEG av den 14 juni 1966 om saluföring av utsäde av foderväxter(), senast ändrat genom direktiv 81/126/EEG(), särskilt artikel 21 a i detta,
De villkor som skall uppfyllas för gröda och utsäde, även standarder för sortrenhet, bör ändras så att de överensstämmer med de system för certifiering av utsäde avsett för internationell handel som fastställts av Organisationen för europeiskt ekonomiskt samarbete (OECD). De datum för genomförandet som fastställts i artikel 2, andra strecksatsen, i kommissionens direktiv 78/386/EEG av den 18 april 1978 om ändring av bilagorna till direktiv 66/401/EEG om saluföring av utsäde av foderväxter(), senast ändrat genom direktiv 81/126/EEG, samt i artikel 2.1 första strecksatsen i kommissionens direktiv 78/388/EEG av den 18 april 1978 om ändring av bilagorna till direktiv 69/208/EEG om saluföring av utsäde av olje- och spånadsväxter(), senast ändrat genom direktiv 81/126/EEG, bör följaktligen anpassas till den aktuella situationen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I andra och tredje meningen i punkt 4 skall orden "Vicia faba" tilläggas efter "Pisum sativum".
Bilaga 2 till direktiv 66/401/EEG ändras på följande sätt:
Artikel 3
- en per 30 m² vid produktion av basutsäde,
Bilaga 2 till direktiv 69/208/EEG ändras på följande sätt:
>Plats för tabell>
I artikel 2.1 andra strecksatsen i direktiv 78/386/EEG skall "den 1 januari 1982" ersättas med "vid ett datum som kommer att fastställas senare".
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa:
- de övriga bestämmelserna i detta direktiv, senast den 1 januari 1983.
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS BESLUT av den 26 oktober 1983 om motåtgärder inom den internationella handelssjöfarten (83/573/EEG)
med beaktande av följande: Utfallet av det informationssystem för sjöfarten som inrättades genom föreskrifterna i besluten 78/774/EEG (), 79/4/EEG (), 80/1181/EEG (), 81/189/EEG () och 82/870/EEG () samt vissa medlemsstaters erfarenhet visar att det skulle vara välbetänkt att inom gemenskapen inrätta ett lämpligt förfarande för motåtgärder inom den internationella handelssjöfarten som berörda medlemsstater kan vidta gentemot tredje länder.
Vid samrådsförfarande enligt artikel 1 bör medlemsstaterna om så är lämpligt i största möjliga utsträckning ange a) den utveckling som har orsakat att motåtgärder vidtagits,
d) den typ av motåtgärder som har vidtagits eller skall vidtas,
Artikel 4
Beslutet riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 54.3 g i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
Kvalifikationskraven måste harmoniseras i fråga om de personer som är behöriga att genomföra lagstadgad revision av räkenskaper. Det bör säkerställas att sådana personer är oberoende och har ett gott anseende.
Medlemsstaterna måste även ges rätt att besluta om övergångsbestämmelser till förmån för yrkesmässigt verksamma personer.
En medlemsstat får godkänna personer som utanför den staten har förvärvat kvalifikationer som är likvärdiga med dem som föreskrivs i detta direktiv.
Frågan om att erkänna ett sådant godkännande att utföra revision som har meddelats en medborgare i en annan medlemsstat kommer att regleras särskilt i direktiv om etablering och utövande av verksamhet inom områdena företagsekonomi, nationalekonomi och redovisning samt i direktiv om frihet att tillhandahålla tjänster inom dessa områden.
Artikel 1
2. Beroende på varje medlemsstats lagstiftning kan de i punkt 1 angivna personerna vara fysiska personer eller juridiska personer eller andra former av bolag eller sammanslutningar (revisionsbolag enligt definitionen i detta direktiv).
1. Lagstadgad revision av de i artikel 1.1 angivna handlingarna får endast utföras av godkända personer. Medlemsstaternas myndigheter får endast godkänna: a) Fysiska personer som uppfyller minst de villkor som anges i artikel 3-19.
iii) En majoritet av ledamöterna i revisionsbolagets förvaltnings- eller ledningsorgan måste vara fysiska personer eller revisionsbolag som uppfyller minst de i artikel 3-19 uppställda villkoren; medlemsstaterna får föreskriva att sådana personer eller revisionsbolag även skall vara godkända. Om ett organ inte har fler än två ledamöter, måste en av dessa minst uppfylla de angivna villkoren.
Artikel 3
En fysisk person får godkännas att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna, endast om han efter att ha kvalificerat sig för tillträde till universitetsstudier har genomgått en teoretisk och praktisk utbildning samt avlagt en statligt organiserad eller godkänd yrkesexamen som är jämförbar med slutexamen från ett universitet.
- balansanalys,
- kostnadsbokföring och internredovisning,
- rättsliga och yrkesmässiga normer för lagstadgad revision och för dem som utför sådan revision,
- beskattningsrätt,
- informations- och databehandling,
- grundläggande principer för ekonomisk styrning av företag.
2. Med avvikelse från bestämmelserna i artikel 5 får en medlemsstat föreskriva att den som har en akademisk examen eller motsvarande kompetens i ett eller flera av de i artikel 6 angivna ämnena får befrias från att avlägga prov som avser hans förmåga att praktiskt tillämpa kunskaperna i dessa ämnen, om han har fått en praktisk utbildning i ämnena som dokumenteras genom av staten erkända examen eller betyg.
2. Medlemsstaterna skall säkerställa att hela den praktiska utbildningen fullgörs hos personer som erbjuder tillräckliga garantier med avseende på utbildningen.
b) att de under sju år har utövat yrkesmässig verksamhet inom de angivna områdena och dessutom har erhållit praktisk utbildning enligt artikel 8 samt har godkänts vid en sådan yrkesexamen som avses i artikel 4.
2. Tiden för den yrkesmässiga verksamheten och den praktiska utbildningen får inte understiga tiden för den teoretiska och praktiska yrkesutbildning som har föreskrivits enligt artikel 4.
b) de skall ha styrkt att de har sådana juridiska kunskaper som i medlemsstaten krävs för lagstadgad revision av de i artikel 1.1 angivna handlingarna. Myndigheterna i medlemsstaten behöver dock inte fordra att sådana kunskaper styrks, om myndigheterna finner att de juridiska kunskaper som har förvärvats i en annan stat är tillräckliga.
1. En medlemsstat får anse sådana yrkesutövare som godkända enligt detta direktiv, vilka har godkänts genom ett förvaltningsbeslut av en behörig myndighet i den medlemsstaten innan de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas.
Till dess att de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas får en medlemsstat anse sådana yrkesutövare som godkända enligt detta direktiv, vilka visserligen inte har godkänts genom förvaltningsbeslut av en behörig myndighet men som dels har samma kvalifikationer i medlemsstaten som de personer vilka har godkänts genom sådana beslut och dels vid tidpunkten för dessa godkännanden utför lagstadgad revision av de i artikel 1.1 angivna handlingarna på de godkända personernas vägnar.
2. Villkoren enligt artikel 2.1 b ii och iii måste uppfyllas senast inom en tidsfrist som inte får överstiga fem år räknat från den tidpunkt då de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas.
Intill ett år efter den tidpunkt då de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas får de yrkesutövare som inte har godkänts genom förvaltningsbeslut av en behörig myndighet, men som i en medlemsstat ändå har rätt att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna och som faktiskt har utfört sådan revision fram till den nämnda tidpunkten, godkännas av medlemsstaten enligt detta direktiv.
1. I sex år räknat från den tidpunkt då de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas får medlemsstaterna vidta övergångsåtgärder för att reglera förhållandena för sådana personer som vid nämnda tidpunkt är i färd med sin teoretiska eller praktiska utbildning, men som då utbildningen avslutas inte skulle uppfylla de villkor som detta direktiv ställer upp och därför inte skulle få utföra den lagstadgade revision av de i artikel 1.1 angivna handlingarna för vilken de har utbildats.
De i artikel 15 och 16 nämnda yrkesutövarna och de i artikel 18 nämnda personerna får med avvikelse från artikel 4 godkännas, endast om de enligt behöriga myndigheters uppfattning är lämpliga att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna och har kvalifikationer som är likvärdiga med dem som innehas av personer som godkänns enligt artikel 4.
b) redan har utfört lagstadgad revision i det ifrågavarande bolaget, innan detta överskred gränserna för två av de tre kriterierna enligt artikel 11 i direktiv 78/660/EEG.
I avvaktan på en senare samordning av den lagstadgade revisionen av räkenskapshandlingar får en medlemsstat - som inte utnyttjar den i artikel 6.1 i direktiv 83/349/EEG angivna möjligheten och i vilken stat, då detta direktiv antas, flera kategorier fysiska personer enligt nationell lagstiftning är behöriga att utföra lagstadgad revision av de i artikel 1.1 b angivna handlingarna - lämna särskilt tillstånd för en person som har godkänts enligt artikel 20 i detta direktiv att utföra lagstadgad revision av de i artikel 1.1 b angivna handlingarna, om på moderbolagets bokslutsdag den grupp av företag vars räkenskaper skall sammanställas sammanlagt enligt företagens senaste årsbokslut inte överskrider gränserna för två av de tre kriterierna i artikel 27 i direktiv 78/660/EEG, förutsatt att personen i fråga är behörig att utföra lagstadgad revision av de i artikel 1.1 a i detta direktiv angivna handlingarna i samtliga de företag som ingår i sammanställningen.
AVSNITT III Yrkesmässig omsorg och oberoende
Artikel 24
Artikel 23 och 24 skall även tillämpas på fysiska personer som uppfyller villkoren i artikel 3-19 och som utför lagstadgad revision av de i artikel 1.1 angivna handlingarna på ett revisionsbolags vägnar.
Artikel 27
Artikel 28
b) Namn och adress för aktieägare eller andra delägare i revisionsbolaget.
AVSNITT V Avslutande bestämmelser
b) vid behov ge kommissionen råd om tillägg till eller ändringar i detta direktiv.
2. Medlemsstaterna får föreskriva att de i punkt 1 avsedda bestämmelserna skall tillämpas först från den 1 januari 1990.
Artikel 31
med beaktande av kommissionens förslag, och
För att säkerställa att stödsystemet fungerar på rätt sätt är det nödvändigt att bestämma för vilka typer av olivolja stöd skall beviljas.
I artikel 20c i den förordningen anges att producentorganisationer och sammanslutningar av producentorganisationer bör utföra vissa kontroll- och samordningsuppgifter. Dessa uppgifter bör därför exakt anges.
Artikel 20d.2 i den förordningen fastställer att endast sammanslutningar skall vara berättigade till förskottsbetalning av stödbeloppet. För att förvaltningen skall skötas på ett riktigt sätt bör detta förskott inte överstiga en viss procentuell andel av stödet.
För att stödsystemet skall fungera på rätt sätt, bör medlemsstaterna bestämma vilken kvantitet av olja som är berättigad till stöd i de fall då den verkliga produktionen av olivolja är oklar.
Artikel 1
4. För olivodlare som är medlemmar i en producentorganisation enligt artikel 20c.1 i förordning nr 136/66/EEG och vars normala produktion inte är mindre än 100 kg olivolja per regleringsår, skall stödet beviljas enligt artikel 5.2 första strecksatsen i den förordningen för den kvantitet olja som verkligen framställts vid en godkänd fabrik, om inte annat följer av artikel 7.
6. Före den 31 mars 1986 skall rådet med kvalificerad majoritet på förslag av kommissionen fastställa de kriterier som skall tillämpas från och med regleringsåret 1986/87 vid bestämmande av de olivodlare som normalt framställer minst 100 kg olja per regleringsår.
- närmare uppgifter om de olivträd som odlas och var de finns,
3. Olivodlare som är medlemmar i en producentorganisation skall, på en dag som skall fastställas, till den organisation som de tillhör lämna en ansökan om individuellt stöd med ett bevis på att oliverna är pressade eller bearbetade, eller en faktura för oliverna eller båda dokumenten.
6. För de olivodlare som inte är medlemmar i en producentorganisation skall den inlämnade individuella skördedeklarationen anses som en ansökan om stöd, förutsatt att den före en dag som skall fastställas kompletteras med:
7. Olivodlare som försummar att uppfylla förpliktelserna i denna artikel skall inte beviljas stöd.
a) i fråga om organisationer som producerar och ökar marknadsvärdet av oliver och olivolja, består av minst 700 olivodlare, eller
2. Endast olivodlare med följande kännetecken får tillhöra en organisation: olivodlare som äger en olivodling som de brukar eller olivodlare som har brukat en olivodling under minst tre år.
4. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att uppmuntra inrättandet av de producentgrupper som anges i förordning (EEG) nr 1360/78 () eller andra organisationer för att framställa och öka marknadsvärdet av oliver och olivolja, vilka kan godkännas som producentorganisationer enligt denna förordning.
2. Senast den 15 oktober skall den behöriga myndigheten, efter att ha mottagit ansökan, fatta beslut om denna efter att ha kontrollerat, om organisationen uppfyller kraven enligt artikel 20c.1 i förordning nr 136/66/EEG och enligt artikel 4, och genast anmäla detta till den berörda organisationen och till kommissionen.
Den behöriga myndigheten skall på grundval av denna anmälan och andra lämpliga undersökningar förvissa sig om att villkoren för godkännande fortfarande är uppfyllda.
1. Godkända producentorganisationer skall
- en gång i månaden överlämna medlemmarnas ansökningar om stöd i ett standardformat som kan användas vid den databearbetning som anges i artikel 16. Stöd skall begäras för den kvantitet som framställts av de medlemmar som har avslutat sin oljeproduktion, förutsatt att de kontroller som anges i artikel 8 har utförts och att de skyldigheter som följer av dessa har uppfyllts.
Artikel 7
- har sålt antingen delar av eller hela sin produktion av olja, och
1. Varje producentorganisation skall, före överlämnandet av ansökningan om stöd, kontrollera den kvantitet av olivolja för vilken stöd söks för var och en av dess medlemmar. Organisationen skall särskilt kontrollera:
2. Producentorganisationer skall överlämna sina medlemsregister till de behöriga myndigheterna i den berörda medlemsstaten i följande fall:
- Om upplysningarna i skördedeklarationen inte stämmer med vad som framkommit vid kontrollerna.
De producentorganisationerna som innefattas i en sammanslutning skall dock komma från minst två ekonomiska regioner.
- skall samordna arbetet i de organisationer som de består av och säkerställa att detta arbete är förenligt med bestämmelserna i denna förordning och skall framförallt snarast kontrollera, enligt ett procenttal som skall bestämmas, på vilket sätt de kontroller som anges i artiklarna 6 och 8 har genomförts,
Artikel 11
b) Saldot skall utbetalas till alla producentorganisationer på grundval av
2. De medlemsstater i vilka olivolja framställs skall garantera att de summor som överlämnats till sammanslutningarna och producentorganisationerna vid tillämpningen av punkt 1 endast används av dem för att finansiera den verksamhet som de är ansvariga för enligt denna förordning.
5. De producerande medlemsstaterna skall fastställa bestämmelser om tilldelningen av stödbelopp och tidsbegränsningar för betalning till olivodlare.
2. Under regleringsåren 1984/1985, 1985/1986 samt 1986/1987 skall det förskott som avses i punkt 1 till varje odlare inte överstiga
Artikel 13
b) har samtyckt till att genomgå alla kontroller som föreskrivs enligt stödförfarandet och till att godkänna alla kontroller som anses nödvändiga i sina lokaler samt att tillåta alla kontroller av deras bokföring,
- inte har fått sitt godkännade indraget för en tid som sträcker sig efter den 31 oktober 1984 enligt den förordningen,
3. Under regleringsåren 1984/1985 och 1985/1986 får de berörda medlemsstaterna bevilja tillfälligt godkännande till den berörda fabriken, så snart en ansökan om godkännande innehållande de upplysningar som anges i punkt 1 har överlämnats.
4. I de fall då ett av villkoren för godkännande enligt punkt 1 inte längre är uppfyllt skall godkännandet återkallas för den tid som är beroende av hur allvarlig överträdelsen är.
eller - någon fysisk eller juridisk person som önskar förestå fabriken i fråga, om inte den personen tillfredsställande kan bevisa för den berörda medlemsstaten att ansökan om nytt godkännande inte är ämnad att kringgå den påförda sanktionen.
2. Producerande medlemsstater skall kontrollera verksamheten i varje producentorganisation och sammanslutning och framförallt kontrollera att kontrollförfarandena har genomförts av dessa organ.
4. Om den olivolja som anges i punkt 1 i bilagan till förordning nr 136/66/EEG framställts av odlare som inte är medlemmar i en producentorganisation, skall kontrollen innebära provtagning på plats som skall bekräfta
Kontrollerna skall ske hos en procentuell andel av odlarna och denna andel skall fastställas på grundval av framför allt företagens storlek.
Artikel 15
2. För producenter vars bokföringsuppgifter har överlämnats till medlemsstaten av deras organisationer enligt artikel 8.2 skall medlemsstaten besluta för vilken kvantitet av olja stödet skall ges. 3. Om resultaten av de kontroller som anges i artiklarna 13 och 14 inte överensstämmer med uppgifterna i lagerbokföringen i en godkänd fabrik, skall den ifrågavarande medlemsstaten, med beaktande av alla sanktioner som får åläggas fabriken, fastställa den kvantitet olja för vilken stöd får beviljas för varje producent som är medlem i en organisation som har pressat sin olivskörd i fabriken i fråga.
1. Varje producerande medlemsstat skall upprätta och underhålla permanenta dataregister innehållande uppgifter om produktionen av oliver och olivolja.
- de upplysningar som finns i den skördedeklaration som föreskrivs i artikel 3.
b) För producentorganisationer och sammanslutningar av dessa: all information som behövs för att kontrollera deras verksamhet i samband med det nuvarande stödsystemet samt även resultaten av de kontroller som utförts av medlemsstaterna.
Artikel 17
- De nationella myndigheter som är bemyndigade av medlemsstaten.
2. De dataregister som upprättas och de program som används för att hantera dem skall vara kompatibla med de datasystem som används för registrering av olivodlingen i varje producerande medlemsstat.
Artikel 19
- De skördar som anges i artikel 18.
För att möjliggöra en smidig övergång från den gällande ordningen till den som fastställs enligt denna förordning, får kommissionen besluta om nödvändiga åtgärder för regleringsåret 1984/85, enligt förfarandet i artikel 38 i förordning nr 136/66/EEG.
Artikel 22
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Europaparlamentets yttrande(),
För att skydda människors och djurs hälsa inom gemenskapen har man i direktiv 72/462/EEG(), senast ändrat genom direktiv 83/91/EEG(), fastställt att medlemsstaternas behöriga myndigheter skall utföra hygienundersökningar vid import av färskt kött och att veterinära experter från medlemsstaterna och kommissionen skall genomföra inspektioner inom det exporterande tredje landet.
I samband med dessa hälsoundersökningar och kontroller debiteras avgifter som för närvarande finansieras på olika sätt i de skilda medlemsstaterna. Dessa skillnader kan påverka de konkurrensvillkor som råder för produkter som till största delen omfattas av en gemensam marknadsordning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
P tar ut avgifter för att täcka kostnaderna för hygienundersökningar och kontroller när ett djur enligt punkt 2 slaktas,
1. Rådet skall på förslag av kommissionen och med kvalificerad majoritet före den 1 januari 1986, fatta beslut om den eller de avgiftsbelopp som avses i artikel 1.1 de första två strecksatserna och om principer och tillämpningsföreskrifter för detta direktiv, samt om möjliga undantag. De avgiftsbelopp som skall debiteras för kött som kommer från slakterier som inte har godkänts enligt direktiv 64/433/EEG skall däremot inte fastställas förrän i samband med att rådet före detta datum har antagit bestämmelser om undersökning av detta kött.
Kommissionen skall före den 1 januari 1990 överlämna en rapport om vunna erfarenheter tillsammans med eventuella förslag till ändringar av de ovannämnda artiklarna.
Grekland skall dock ha en ytterligare tidsfrist på två år för att följa det.
med beaktande av kommissionens förslag(),
med beaktande av följande: Enligt fördraget är all särbehandling som grundar sig på nationalitet när det gäller etablering och tillhandahållande av tjänster förbjuden fr.o.m. övergångsperiodens utgång. Principen om sådan behandling som grundar sig på nationalitet förekommer särskilt vid beviljande av de tillstånd som krävs för att utöva vissa former av verksamhet samt inregistrering eller medlemskap i yrkesorganisationer eller motsvarande organ.
Som villkor för att få utöva viss farmaceutisk verksamhet krävs i några medlemsstater förutom utbildnings-, examens- och andra behörighetsbevis en kompletterande yrkeserfarenhet; då det ännu inte föreligger någon överensstämmelse mellan medlemsstaterna inom detta område bör, för att undvika svårigheter, lämplig praktisk yrkeserfarenhet av samma längd som förvärvats i en annan medlemsstat erkännas som tillräcklig.
För att underlätta tillämpningen av detta direktiv för de nationella myndigheterna får en medlemsstat föreskriva att den person som uppfyller utbildningsvillkoren enligt detta direktiv samtidigt med de formella utbildningsbevisen skall förete ett intyg från de behöriga myndigheterna i ursprungslandet eller det senaste hemvistlandet som visar att dessa bevis är de som avses i direktivet.
När det gäller kraven på god vandel och gott anseende bör skillnad göras mellan de krav som ställs för att påbörja verksamhet inom yrket och de krav som ställs för att få utöva yrket.
Artikel 1
2. Medlemsstaterna är emellertid inte skyldiga att låta de utbildnings-, examens- och andra behörighetsbevis som avses i punkt 1 träda i kraft när det gäller att inrätta nya apotek som är öppna för allmänheten. Vid tillämpningen av detta direktiv skall apotek som varit i drift kortare tid än tre år betraktas som nyinrättade.
1. Utan hinder av artikel 2 och utan att det påverkar tillämpningen av artikel 45 i 1979 års anslutningsakt skall Grekland endast åläggas att tillämpa bestämmelserna i artikel 2 om de utbildnings-, examens- och andra behörighetsbevis som utfärdas av de övriga medlemsstaterna, såvida det gäller utövande av de former av verksamhet som avses i artikel 1 som anställd i enlighet med förordning (EEG) nr 1612/68.
Artikel 4
Le diplôme légal de pharmacien/het wettelijk diploma van apoteker (det lagstadgade examensbeviset i farmaci) som utfärdas av universitetens medicinska och farmaceutiska fakulteter, av centrala examensnämnden eller av de statliga examensnämnderna för universitetsutbildningen.
c) I Tyskland:
d) I Grekland:
Statligt examensbevis som utfärdas av universiteten eller statligt examensbevis som farmacie doktor som utfärdas av universiteten.
g) I Italien:
Statligt examensbevis som farmaceut som utfärdas av statens examensnämnd och undertecknas av utbildningsministern.
j) I Storbritannien:
Om det i en medlemsstat inte bara krävs ett utbildnings-, examens- eller annat behörighetsbevis för att påbörja eller utöva någon form av verksamhet som avses i artikel 1 utan även kompletterande yrkeserfarenhet, skall det landet som tillräckligt bevis godta ett intyg utfärdat av de behöriga myndigheterna i ursprungslandet eller det senaste hemvistlandet som visar att personen i fråga har utövat nämnda former av verksamhet under motsvarande period i ursprungslandet eller det senaste hemvistlandet.
De utbildnings-, examens- och andra behörighetsbevis i farmaci som medlemsstaterna utfärdat till medborgare i medlemsstaterna och som inte uppfyller de minimivillkor för utbildningen som fastställts i artikel 2 i direktiv 85/432/EEG skall jämställas med de examensbevis som uppfyller dessa krav,
KAPITEL IV Användning av akademisk titel
2. Om den akademiska titel som används i ursprungslandet eller det senaste hemvistlandet kan förväxlas med en titel som i värdlandet kräver kompletterande utbildning, som personen i fråga inte har genomgått, får värdlandet kräva att denne använder den först nämnda titeln i en lämplig form som värdlandet anger.
2. Om det i ursprungslandet eller det senaste hemvistlandet inte krävs bevis om god vandel eller bevis om gott anseende för att påbörja verksamheten i fråga, får värdlandet kräva att personen i fråga företer utdrag ur kriminalregistret eller eventuellt motsvarande handling utfärdad av en behörig myndighet i ursprungslandet eller det senaste hemvistlandet.
1. Om det i värdlandet finns bestämmelser i lagar och andra författningar om krav på god vandel eller gott anseende samt bestämmelser om disciplinpåföljd i händelse av allvarligt fel i yrkesutövningen eller fällande dom på grund av lagöverträdelser i samband med den yrkesutövning som avses i artikel 1, skall ursprungslandet eller det senaste hemvistlandet till värdlandet överlämna alla upplysningar som behövs om de åtgärder eller disciplinpåföljder av yrkesmässig eller administrativ karaktär som vidtagits mot personen i fråga eller om de straffrättsliga påföljder på grund av lagöverträdelser som ådömts denne under yrkesutövningen i ursprungslandet eller det senaste hemvistlandet.
3. Medlemsstaterna skall garantera de lämnade upplysningarnas konfidentiella natur. Artikel 10
Artikel 11
1. Det förfarande som genomförs enligt artikel 8, 9 och 10 för att personen i fråga skall beviljas tillstånd att utöva sådan verksamhet som avses i artikel 1 avslutas snarast möjligt och senast tre månader efter det att samtliga handlingar som rör denna person inlämnats med beaktande av de förseningar som kan uppstå på grund av eventuella överklaganden efter det att detta förfarande genomförts.
Efter att ha mottagit svaret eller efter tidsfristens utgång skall värdlandet fortsätta det förfarande som avses i punkt 1.
Artikel 14
1. Medlemsstaterna skall vidta nödvändiga åtgärder för att göra det möjligt för personerna i fråga att erhålla upplysningar om hälso- och socialförsäkringslagstiftningen och, där så är tillämpligt, om de yrkesetiska reglerna i värdlandet.
3. Medlemsstaterna skall se till att, där så är lämpligt, personerna i fråga i deras eget och deras patienters intresse förvärvar de språkkunskaper som krävs för att utöva yrket i värdlandet.
Artikel 17
Detta direktiv skall även tillämpas på de medborgare i medlemsstaterna som i enlighet med förordning (EEG) nr 1612/68 i egenskap av anställda utövar eller kommer att utöva sådan verksamhet som avses i artikel 1. Artikel 19
Artikel 20
Artikel 21
med beaktande av kommissionens förslag (1),
med beaktande av följande:Medlemsstaternas författningsregler beträffande företag för kollektiva investeringar varierar avsevärt, särskilt i fråga om de skyldigheter och den övervakning som gäller för sådana företag. Dessa olikheter inverkar negativt på villkoren för konkurrens mellan företagen och ger inte likvärdigt skydd för andelsägarna.
Samordningen av medlemsstaternas lagstiftning skall till en början begränsas till att avse företag för kollektiva investeringar av icke sluten typ som utbjuder sina andelar till allmänheten inom gemenskapen och som har som enda syfte att investera i överlåtbara värdepapper (dvs. väsentligen överlåtbara värdepapper som är officiellt noterade vid fondbörser eller liknande reglerade marknadsplatser). Regleringen av företag för kollektiva investeringar som inte omfattas av direktivet erbjuder en mängd problem som måste lösas med hjälp av andra bestämmelser, och sådana företag kommer följaktligen att bli föremål för samordning i ett senare skede. I avvaktan på sådan samordning får varje enskild medlemsstat bl.a. från direktivets tillämpningsområde undanta kategorier av företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag) som har speciell placerings- och upplåningsinriktning och uppställa särskilda regler för dessa företags verksamhet inom den medlemsstaten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Vid tillämpningen av detta direktiv skall med värdepappersfonder avses även "unit trusts".
6. Med förbehåll för bestämmelserna om kapitalrörelser och bestämmelserna i artiklarna 44, 45 och 52.2 får en medlemsstat, i de avseenden som regleras i detta direktiv, inte tillämpa andra bestämmelser för fondföretag hemmahörande i en annan medlemsstat, eller för andelar som utgivits av sådana företag, i de fall de utbjuder sina andelar inom medlemsstatens territorium.
- Fondföretag vars andelar enligt fondbestämmelserna eller bolagsordningen får säljas endast till allmänheten i icke-medlemsländer.
Artikel 3
Artikel 4
2. En värdepappersfond får auktoriseras endast om de behöriga myndigheterna godkänt förvaltningsbolaget, fondbestämmelserna och valet av förvaringsinstitut. Ett investeringsbolag får auktoriseras endast om de behöriga myndigheterna godkänt både dess bolagsordning och valet av förvaringsinstitut.
4. Utan de behöriga myndigheternas godkännande får varken förvaltningsbolaget eller förvaringsinstitutet bytas ut, eller fondbestämmelserna eller investeringsbolagets bolagsordning ändras.
Ett förvaltningsbolag skall ha finansiella resurser som är tillräckliga för att bolaget skall kunna bedriva sin verksamhet på ett effektivt sätt och uppfylla sina förpliktelser.
Artikel 7
d) tillse att ersättningar för transaktioner som berör en värdepappersfonds tillgångar inbetalas till institutet inom sedvanlig tid,
1. Ett förvaringsinstitut skall antingen ha sitt stadgeenliga säte i samma medlemsstat som förvaltningsbolaget eller vara etablerat där om det har sitt stadgeenliga säte i en annan medlemsstat.
Artikel 9
1. Ett företag får inte samtidigt vara förvaltningsbolag och förvaringsinstitut.
Villkoren för utbyte av förvaltningsbolaget eller förvaringsinstitutet skall, liksom regler till skydd för andelsägare vid sådana utbyten, föreskrivas i lag eller annan författning eller anges i fondbestämmelserna.
Medlemsstaterna skall bestämma vilken rättslig form ett investeringsbolag skall ha. Ett investeringsbolag skall ha ett så stort inbetalt kapital att det kan bedriva verksamheten effektivt och uppfylla sina förpliktelser.
Artikel 14
3. Ett förvaringsinstitut skall vidare
4. En medlemsstat får besluta att investeringsbolag som hör hemma i den staten och som utbjuder sina andelar uteslutande på en eller flera fondbörser där andelarna är officiellt noterade, inte skall vara skyldiga att anlita förvaringsinstitut som avses i detta direktiv.
En medlemsstat får utnyttja den möjlighet som ges i föregående stycke endast om den finner att andelsägarna har ett skydd som är likvärdigt med det som tillkommer andelsägare i fondföretag med förvaringsinstitut som avses i detta direktiv.
Minst två gånger per månad skall en oberoende revisor kontrollera att andelarnas värde beräknas i enlighet med lag eller annan författning och med bolagsordningen. Vid sådana tillfällen skall revisorn kontrollera att bolagets tillgångar är placerade i enlighet med lag eller annan författning och med bolagsordningen.
Artikel 15
3. Medlemsstaterna skall bestämma vilka av de kategorier av institut som avses i punkt 2 som skall kunna utses till förvaringsinstitut.
Artikel 17
Artikel 18
Artikel 19
a) ett fondföretag får placera högst 10% av sina fondtillgångar i andra överlåtbara värdepapper än de som avses i punkt 1,
d) ett fondföretag inte får förvärva ädla metaller eller värdepapper inlösbara i sådana metaller.
Artikel 20
2. Medlemsstaterna får också ge fondföretag tillstånd att vid förvaltningen av sina tillgångar och skulder utnyttja sådan teknik och sådana instrument som syftar till att ge skydd mot valutarisker.
2. Medlemsstaterna får höja den gräns som anges i punkt 1 till högst 10%. I den mån fondföretaget placerar mer än 5% av fondtillgångarna i överlåtbara värdepapper med samme utgivare, får det sammanlagda innehavet av sådana placeringar inte överstiga 40% av fondtillgångarna.
1. Utan hinder av artikel 22, med förbehåll för artikel 68.3 i fördraget, får medlemsstaterna ge fondföretag tillstånd att med tillämpning av principen om riskspridning placera upp till 100% av fondtillgångarna i olika överlåtbara värdepapper utgivna eller garanterade av en medlemsstat, dess lokala myndigheter, en icke-medlemsstat eller offentliga internationella organ i vilka en eller flera medlemsstater är medlemmar.
2. Fondbestämmelserna eller bolagsordningarna för de fondföretag som avses i punkt 1 skall innehålla uttrycklig uppgift om de stater, lokala myndigheter och offentliga internationella organ som utger eller garanterar sådana värdepapper i vilka fondföretaget avser att placera mer än 35% av fondtillgångarna; sådana fondbestämmelser och bolagsordningar måste godkännas av behöriga myndigheter.
1. Ett fondföretag får inte förvärva fondandelar i andra företag för kollektiva investeringar av den öppna typen, såvida dessa inte är företag för kollektiva investeringar i den betydelse som avses i första och andra strecksatserna i artikel 1.2.
Ett förvaltningsbolag får inte debitera några avgifter eller kostnader för transaktioner som hänför sig till en viss värdepappersfonds andelar i fall där några av en värdepappersfonds tillgångar är placerade i andelarna i en annan värdepappersfond som förvaltas av samma förvaltningsbolag eller av ett annat bolag med vilket förvaltningsbolaget är anknutet via gemensam företagsledning eller ägarkontroll eller genom ett betydande direkt eller indirekt ägande.
I avvaktan på vidare samordning skall medlemsstaterna beakta gällande föreskrifter i andra medlemsstaters lagstiftning, som närmare uttrycker den i föregående stycke angivna principen.
De gränsvärden som anges i andra och tredje strecksatserna behöver inte iakttas vid förvärvstillfället, om bruttomängden av skuldebreven eller nettomängden av de värdepapper som är under utgivning då inte kan uppskattas.
Artikel 26
2. Om gränsvärdena enligt punkt 1 överskrids av skäl som ligger utanför ett fondföretags rådighet eller som följd av att teckningsrätter utnyttjas, skall fondföretaget vid sina försäljningstransaktioner prioritera rättelse av detta förhållande under vederbörligt hänsynstagande till andelsägarnas intressen. AVSNITT VI
1. Ett investeringsbolag och ett förvaltningsbolag, det senare för varje värdepappersfond det förvaltar, skall offentliggöra
1. Ett prospekt skall innehålla den information som krävs för att investerare skall kunna göra en välgrundad bedömning av den erbjudna investeringen. Prospektet skall innehålla minst den information som anges i lista A i bilagan till detta direktiv, såvida inte informationen redan framgår av de handlingar som skall bifogas prospektet enligt artikel 29.1.
Artikel 29
Artikel 30
De uppgifter om räkenskaperna som årsrapporten innehåller skall vara granskade av en eller flera personer som enligt lag eller annan författning bemyndigats att granska redovisningar i överensstämmelse med rådets direktiv 84/253/EEG av den 10 april 1984 grundat på artikel 54.3 g i Romfördraget, om godkännande av personer som har ansvar för lagstadgad revision av räkenskaper (4). Revisionsberättelsen, med eventuella anmärkningar, skall i sin helhet återges i årsrapporten.
Artikel 33
3. Årsrapporterna och halvårsrapporterna skall på begäran kostnadsfritt tillställas andelsägarna.
Ett fondföretag skall vid varje tillfälle då det emitterar, säljer, återköper eller löser in andelar, dock minst två gånger per månad, på lämpligt sätt offentliggöra emissions-, försäljnings-, återköps- och inlösenpriserna. De behöriga myndigheterna får dock medge ett fondföretag att offentliggöra sådana uppgifter endast en gång per månad, förutsatt att andelsägarnas intressen inte härigenom åsidosätts.
Fondföretags allmänna förpliktelser
a) upp till 10% - av tillgångarna, i fråga om ett investeringsbolag eller,
Artikel 37
3. I de fall som avses i punkt 2 a, skall ett fondföretag utan dröjsmål underrätta de berörda myndigheterna och myndigheterna i samtliga medlemsstater där företaget utbjuder sina andelar om uppskovsbeslutet.
Artikel 39
Ett fondföretags andelar får emitteras endast om fondtillgångarna inom sedvanlig tid tillförs betalning motsvarande emissionens nettopris. Denna bestämmelse skall inte utgöra hinder för tilldelning av bonusandelar.
- ett förvaltningsbolag eller förvaringsinstitut som handlar för en värdepappersfonds räkning får bevilja lån eller ingå borgen för någon annans räkning.
Artikel 43
AVSNITT VIII Särskilda bestämmelser för fondföretag som utbjuder sina andelar i andra medlemsstater än dem där företagen är hemmahörande
2. Ett fondföretag får marknadsföra sina andelar i de medlemsstater där dessa utbjuds. Det måste därvid följa de bestämmelser om reklam som gäller i det landet.
I det fall som avses i artikel 44 skall fondföretagen, i enlighet med de lagar och andra författningar som gäller i den medlemsstat där andelarna utbjuds, bl.a. vidta erforderliga åtgärder för att där kunna göra utbetalningar till andelsägarna, verkställa återköp och inlösen samt lämna ut den information som fondföretagen är skyldiga att tillhandahålla.
- sitt prospekt,
Artikel 48
Artikel 49
3. Myndigheterna i den stat där ett fondföretag är hemmahörande skall vara behöriga att utöva tillsyn över företaget. Myndigheterna i den stat där ett fondföretag utbjuder sina andelar i enlighet med artikel 44 skall dock vara behöriga att kontrollera att bestämmelserna i avsnitt VIII följs.
1. De medlemsstaters myndigheter som avses i artikel 49 skall fullgöra sina uppgifter i nära samarbete och utbyta nödvändig information.
4. Utöver vad som följer av straffrättsliga föreskrifter får en myndighet som avses i artikel 49 och som erhåller ifrågavarande information använda denna endast för fullgörande av sina uppgifter samt vid överklaganden i administrativ ordning och vid rättsliga förfaranden som har samband med myndighetens verksamhet.
2. Medlemsstaterna skall sörja för att beslut som fattas med avseende på fondföretag med stöd av lag eller annan författning i enlighet med detta direktiv kan prövas av domstol. En möjlighet till domstolsprövning skall finnas också för fall då beslut inte fattats inom sex månader från det att ett fondföretag lämnat in auktorisationsansökan som innehåller all den information som krävs enligt gällande föreskrifter.
2. Myndigheterna i den medlemsstat där ett fondföretags andelar utbjuds får dock vidta åtgärder mot företaget, om det bryter mot de i avsnitt VIII nämnda bestämmelserna.
Artikel 53
b) att underlätta samråd mellan medlemsstater antingen beträffande skärpta eller kompletterande krav som de har rätt att uppställa i enlighet med artikel 1.7, eller beträffande föreskrifter som de får utfärda i enlighet med artiklarna 44 och 45,
3. Kommittén skall vara sammansatt av personer utsedda av medlemsstaterna och av representanter för kommissionen. Ordföranden skall vara en representant för kommissionen. Sekretariatstjänster skall tillhandahållas av kommissionen.
Artikel 54
Trots bestämmelserna i artiklarna 7.1 och 14.1 får de behöriga myndigheterna tillåta sådana fondföretag som i enlighet med nationell lagstiftning hade två eller flera förvaringsinstitut vid tidpunkten för antagandet av detta direktiv att behålla dessa institut, om myndigheterna har garantier för att de uppgifter som föreskrivs i artiklarna 7.3. och 14.3 kommer att fullgöras i praktiken.
2. Medlemsstaterna får bevilja förvaltningsbolag som, vid tidpunkten för antagande av detta direktiv bedriver andra verksamheter än sådana som tillåts enligt artikel 6, att fortsätta med dessa i fem år efter nämnda tidpunkt.
2. Medlemsstaterna får bevilja fondföretag, som var verksamma vid tidpunkten för genomförandet av detta direktiv en frist om högst 12 månader från den tidpunkten att anpassa sig till den nya nationella lagstiftningen.
Kommissionen skall, om så erfordras, föreslå att rådet förlänger uppskovet upp till fyra år.
Artikel 59
med beaktande av kommissionens förslag (1),
med beaktande av följande: En harmonisk utveckling av den ekonomiska verksamheten samt en varaktig och balanserad tillväxt inom gemenskapen som helhet är beroende av att det upprättas en gemensam marknad som fungerar tillfredsställande och erbjuder villkor som motsvarar dem som råder på den nationella marknaden. För att få till stånd denna gemensamma marknad och stärka dess enhet bör rättsliga grundvalar skapas som underlättar för fysiska personer, bolag och andra rättsliga enheter att anpassa sin verksamhet till gemenskapens ekonomiska villkor. Det är därför nödvändigt att dessa fysiska personer, bolag och andra rättsliga enheter kan samarbeta effektivt över gränserna.
En grupperings förmåga att anpassa sig till de ekonomiska villkoren bör garanteras genom en avsevärd handlingsfrihet för grupperingens medlemmar att reglera sina avtalsmässiga förbindelser och grupperingens interna organisation.
Enbart denna förordning ger inte rätt att delta i en gruppering, även om villkoren som föreskrivs i förordningen är uppfyllda.
Skyddet för tredje man kräver en hög grad av offentlighet. Medlemmarna ansvarar obegränsat solidariskt för grupperingens skulder och andra förbindelser, inklusive skulder avseende skatter och sociala avgifter, dock utan att denna princip inverkar på rätten att genom ett särskilt avtal mellan grupperingen och en tredje man bestämma att ansvaret skall uteslutas eller begränsas i fråga om en eller flera medlemmar när det gäller en viss skuld eller någon annan förbindelse.
En gruppering omfattas av bestämmelserna i nationell lagstiftning om obestånd och betalningsinställelse. Dessa bestämmelser kan ange ytterligare grunder för upplösning av grupperingen.
- social- och arbetsrätt,
En gruppering är underkastad medlemsstaternas rättsregler om utövande av verksamheten och kontroll av denna. Om en gruppering eller dess medlemmar missbrukar eller kringgår en medlemsstats lagstiftning får medlemsstaten tillgripa lämpliga sanktioner.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. En gruppering får därför inte
c) ha fler än 500 anställda,
Artikel 4
b) Fysiska personer som utövar industri-, handels-, hant- verks- eller jordbruksverksamhet eller ett fritt yrke eller annan verksamhet inom gemenskapen.
b) två fysiska personer som avses i punkt 1 och som bedriver sin huvudsakliga verksamhet i olika medlemsstater, eller
4. Varje medlemsstat kan med hänsyn till sina allmänna intressen förbjuda eller begränsa rätten för vissa kategorier av fysiska personer, bolag eller andra rättsliga enheter att delta i grupperingar.
a) Grupperingens namn, föregånget eller följt av antingen orden "europeisk ekonomisk intressegruppering" eller förkortningen "EEIG", om inte dessa ord eller denna förkortning redan ingår i namnet.
d) För varje medlem namn, firma, rättslig organisationsform, bostadsadress eller adress för säte samt i förekommande fall registreringsnummer och registreringsort.
I den stat där en gruppering har sitt säte skall den tas in i ett register enligt artikel 39.1.
Följande handlingar och uppgifter skall också ges in till registret: a) Varje ändring i avtalet om att bilda grupperingen, däribland varje ändring i grupperingens sammansättning.
d) Uppgift om vem eller vilka som har utsetts till företagsledare för grupperingen, vederbörandes namn och övriga personuppgifter som krävs enligt lagstiftningen i den medlemsstat där registret förs, uppgift huruvida företagsledarna kan handla var för sig eller om de måste handla i förening samt uppgift om när uppdraget för en företagsledare har upphört.
g) Uppgift om att enligt artikel 35 en eller flera likvidatorer har tillsatts för en gruppering, vederbörandes namn och övriga personuppgifter som krävs enligt lagstiftningen i den medlemsstat där registret förs samt uppgift om när uppdraget för en likvidator har upphört.
j) Avtalsvillkor enligt artikel 26.2 som befriar en ny medlem från ansvar för skulder och andra förpliktelser som har uppkommit innan han antogs som medlem.
a) De obligatoriska uppgifter som enligt artikel 5 skall anges i avtalet om att bilda en gruppering och ändring i dessa uppgifter.
De i a och b angivna uppgifterna skall offentliggöras i sin helhet. I c angivna handlingar och uppgifter skall offentliggöras antingen i sin helhet eller i form av ett utdrag eller ett meddelande om att de har givits in till registret enligt tillämplig nationell lagstiftning.
2. Har handlingar företagits i en grupperings namn innan grupperingen registrerats enligt artikel 6 och åtar sig inte grupperingen efter registreringen att svara för de förbindelser som följer med dessa handlingar, svarar de fysiska personer, bolag eller andra rättsliga enheter som har företagit handlingarna obegränsat solidariskt för dessa.
Artikel 11
Det säte som anges i avtalet om att bilda en gruppering skall finnas inom gemenskapen.
b) i den ort där någon av grupperingens medlemmar har sitt huvudkontor eller, när det är fråga om en fysisk person, utövar sin huvudsakliga verksamhet, förutsatt att grupperingen är verksam där.
Beslut om bytet skall fattas enligt vad som är bestämt i avtalet om att bilda grupperingen, om inte bytet medför att enligt artikel 2 någon annan lagstiftning blir tillämplig.
Beslut om bytet får fattas först två månader efter det att förslaget har offentliggjorts. Beslutet fattas enhälligt av medlemmarna. Det får verkan från den dag då grupperingen enligt artikel 6 tas in i det nya registret. Innan registreringen äger rum måste det visas att förslaget till byte har offentliggjorts.
4. En medlemsstat kan i fråga om grupperingar som enligt artikel 6 är registrerade i den staten föreskriva i sin lagstiftning att ett byte av säte, som skulle medföra att annan lagstiftning blev tillämplig, inte skall få verkan om en behörig myndighet i den nämnda staten motsätter sig bytet inom den i punkt 1 angivna tvåmånadersfristen. En sådan invändning får endast grunda sig på allmänna intressen. Den skall kunna prövas av domstol.
2. En grupperings ogiltighet medför likvidation av grupperingen enligt artikel 35.
Artikel 16
2. Grupperingens medlemmar kan i egenskap av organ för denna fatta alla beslut som syftar till att förverkliga ändamålet med grupperingen.
2. Medlemmarna kan endast enhälligt besluta att
c) ändra förutsättningarna för att fatta beslut,
f) ändra någon annan förpliktelse som åligger en medlem, om inte annat är bestämt i avtalet om att bilda grupperingen,
Varje medlem har rätt att få upplysningar av företagsledarna om grupperingens verksamhet samt att granska grupperingens böcker och affärshandlingar.
Till företagsledare i en gruppering kan inte utses någon som
- enligt ett avgörande av domstol eller annan myndighet som har beslutats eller erkänts inom en medlemsstat
En medlemsstat som begagnar sig av den nu angivna möjligheten skall föreskriva att representanterna skall ha samma ansvar som företagsledarna.
Artikel 20
En begränsning i företagsledarnas rätt att företräda grupperingen i avtalet om att bilda denna eller genom beslut av medlemmarna får inte åberopas mot tredje man, även om begränsningen har offentliggjorts.
1. Vinsten av en grupperings verksamhet skall anses som medlemmarnas egen vinst och delas mellan dem enligt vad som är bestämt i avtalet om att bilda grupperingen eller, om sådana bestämmelser saknas, i lika delar.
1. Varje medlem i en gruppering kan överlåta sin andel i denna eller en del av andelen till någon annan medlem eller till tredje man; överlåtelsen får verkan endast om grupperingens övriga medlemmar enhälligt har tillåtit denna.
En gruppering får inte rikta placeringserbjudanden till allmänheten. Artikel 24
Artikel 25
b) Orten för det register enligt artikel 6 i vilket grupperingen är införd och grupperingens registreringsnummer.
e) I förekommande fall att grupperingen har trätt i likvidation enligt artikel 15, 31, 32 eller 36.
1. Ett beslut att anta en ny medlem skall fattas enhälligt av medlemmarna.
Artikel 27
Artikel 28
2. Om en medlem dör, kan någon annan inträda i grupperingen i den avlidnes ställe endast på de villkor som är bestämda i avtalet om att bilda grupperingen eller efter samtycke av alla övriga medlemmar.
Artikel 30
1. En gruppering får upplösas genom ett beslut av medlemmarna om detta. Ett sådant beslut skall fattas enhälligt om inte något annat är bestämt i avtalet om att bilda grupperingen. 2. En gruppering skall upplösas genom ett beslut av medlemmarna, om
Varje medlem får ansöka om att rätten skall bestämma att upplösning skall ske, om medlemmarna ännu tre månader efter det att en i a eller b angiven omständighet har inträffat inte har beslutat om upplösning.
Artikel 32
3. En medlemsstat kan bestämma att rätten på ansökan av en behörig myndighet inom den staten får förordna att en gruppering med säte inom staten skall upplösas om grupperingen åsidosätter allmänna intressen inom staten, allt under förutsättning att det enligt statens lagstiftning är möjligt att på sådan grund upplösa registrerade bolag eller andra rättsliga enheter.
Värdet av en avgående medlems rättigheter och skyldigheter får inte bestämmas i förväg.
Artikel 35
3. Grupperingen behåller sin rättskapacitet enligt artikel 1.2 till dess likvidationen är avslutad.
En gruppering omfattas av nationell lagstiftning om obestånd och betalningsinställelse. Enbart det förhållandet att ett rättsligt förfarande inleds mot en gruppering på grund av dennas obestånd eller betalningsinställelse får inte medföra att ett sådant förfarande inleds mot medlemmarna.
2. En preskriptionstid på fem år räknat från offentliggörandet enligt artikel 8 av avslutandet av en grupperings likvidation gäller i stället för längre preskriptionstider i nationell lagstiftning i fråga om åtgärder mot en medlem med anledning av förbindelser som har uppkommit genom grupperingens verksamhet.
1. Medlemsstaterna skall inrätta det eller de register som skall svara för registrering enligt artiklarna 6 och 10, samt meddela regler om registreringen. De skall bestämma hur handlingarna som avses i artiklarna 7 och 10 skall ges in. De skall se till att de handlingar och uppgifter som avses i artikel 8 offentliggörs i en lämplig officiell tidning inom den medlemsstat där grupperingen har sitt säte, samt får bestämma hur de handlingar och uppgifter som avses i artikel 8 c skall offentliggöras.
2. Medlemsstaterna skall se till att de upplysningar som enligt artikel 11 skall offentliggöras i Europeiska gemenskapernas officiella tidning sänds till kontoret för de Europeiska gemenskapernas officiella publikationer inom en månad efter offentliggörandet i den officiella tidning som avses i punkt 1.
Endast medlemmarna skall beskattas för resultatet av en grupperings verksamhet.
2. För kännedom skall en medlemsstat underrätta kommissionen om vilka kategorier av fysiska personer, bolag och andra rättsliga enheter som medlemsstaten enligt artikel 4.4 har förbjudit att delta i en gruppering. Kommissionen skall underrätta de övriga medlemsstaterna om förbudet.
a) med förbehåll för artiklarna 169 och 170 i Romfördraget underlätta tillämpningen av förordningen genom regelbundet samråd, särskilt om praktiska problem i samband med tillämpningen,
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: Genom rådets förordning (EEG) nr 3284/83(4) ändras bestämmelserna för beviljande av stöd till frukt- och grönsaksproducenters organisationer.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av rådets förordning (EEG) nr 3117/85 av den 4 november 1985 om allmänna bestämmelser för beviljande av ekonomisk kompensation avseende sardiner(), särskilt artikel 4 i denna, och
De hygienföreskrifter och tekniska bestämmelser som fastställts av de nationella myndigheterna bör säkerställa att produkterna i fråga fullständigt och slutligt beretts i någon av de former som anges i artikel 3.1 i förordning (EEG) nr 3117/85. Det bör kontrolleras att de beredda produkterna överensstämmer med dessa bestämmelser.
För att kunna möjliggöra en fortlöpande kontroll bör bidragsmottagarna hela tiden hålla tillsynsmyndigheten underrättad om sin beredningsverksamhet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. De beredningsprocesser som avses i punkt 1 är
c) filetering eller styckning i förening med en av de beredningsformer som avses i a och b.
Artikel 4
- I fält 41 en beskrivning av varorna i det tillstånd de befann sig vid tidpunkten för avsändandet.
såvida det vid utbetalningstillfället inte finns uppgifter som tyder på att produkterna inte har beretts fullständigt och slutligt.
Artikel 6
- Inspektioner av beredningsföretagen på plats.
- Identifiering genom producentorganisationens försäljningsjournal av de kvantiteter som sålts enligt denna ordning.
2. Medlemsstaterna skall också varje månad till kommissionen anmäla de kvantiteter som sålts under den föregående månaden som berättigar till stöd, fördelade på handelskategorier och beredningsformer, samt kostnaderna för beviljandet av stödet i fråga.
Den omvandlingskurs som skall gälla för bidraget är den på försäljningsdagen gällande representativa kursen.
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), senast ändrad genom förordning (EEG) nr 1298/85(2), särskilt artikel 6.7 i denna, och
Artikel 1
Artikel 2
med beaktande av kommissionens förslag (),
med beaktande av följande: Enligt artikel 2 i fördraget har gemenskapen särskilt till uppgift att främja en harmonisk utveckling av den ekonomiska verksamheten inom gemenskapen som helhet, en fortgående och balanserad tillväxt, en ökad stabilitet, samt närmare förbindelser mellan de stater som gemenskapen förenar. Turism kan bidra till att uppnå dessa mål.
Varje medlemsstat bör låta de andra medlemsstaterna och kommissionen dra fördel av sin erfarenhet inom turistområdet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE
Artikel 2
För de ändamål som anges i artikel 2 skall varje medlemsstat översända en rapport till kommissionen en gång om året om de viktigaste åtgärderna som den har vidtagit och, så långt möjligt, om de åtgärder den avser att vidta i fråga om sådana tjänster för turister som skulle kunna få konsekvenser för resande från andra medlemsstater.
3. Kommittén skall också råda kommissionen i de frågor där kommissionen har begärt ett yttrande.
Kommissionen skall utöva ordförandeskapet i kommittén.
med beaktande av följande: Med anledning av Portugals anslutning är det nödvändigt att göra vissa ytterligare tekniska ändringar av direktiv 85/384/EEG() i dess lydelse enligt direktiv 85/614/EEG() för att säkerställa att det tillämpas på samma sätt av Portugal och de andra medlemsstaterna.
Artikel 1
med beaktande av följande: I artikel 2.1 i förordning (EEG) nr 426/86 föreskrivs ett system för produktionsstöd för vissa produkter. I artikel 6.1 b i samma förordning föreskrivs att stödet endast skall betalas ut för produkter som uppfyller vissa minimikvalitetskrav som skall fastställas.
De kvalitetskrav som fastställs i denna förordning ingår i åtgärderna för genomförandet av systemet med produktionsstöd. Gemenskapen har ännu inte fastställt kvalitetskraven i samband med saluföring av produkterna. Medlemsstaterna får för detta ändamål fortsätta att tillämpa nationella krav under förutsättning att de är förenliga med fördragets bestämmelser om fri rörlighet för varor.
Artikel 1
Artikel 3
Artikel 4
P tomatsaft,
P naturliga kryddor, kryddörter och extrakt av dessa samt naturliga aromämnen.
3. Tillsatt tomatsaft och tomatkoncentrat skall uppfylla de minimikrav som fastställs i avdelning II.
2. Skalade tomater skall vara praktiskt taget fria från skal. Hela skalade tomater skall dessutom vara praktiskt taget fria från skadade delar.
1. Produkterna skall anses uppfylla kraven i artikel 5.2 om följande gränsvärden för skador inte överskrids:
P hela tomater: 300 cm2 sammantagen yta,
2. I punkt 1 avses med
Artikel 7
3. Om skalade konserverade tomater förpackas i glasburkar skall volymen minskas med 20 ml innan de procenttal som avses i punkterna 1 och 2 beräknas.
Artikel 9
P naturliga kryddor, kryddörter och extrakt av dessa samt naturliga aromämnen.
P tomatkoncentrat i pulverform, får kiseldioxid (551) användas. Innehållet av kiseldioxid skall dock inte överstiga 1 % av den färdiga produktens vikt.
b) 3 viktprocent av nettovikten för andra tomatkoncentrat och för tomatsaft.
1. Tomatsaft och tomatkoncentrat skall ha
Produkterna skall vara fria från främmande smaker, särskilt smaken av bränd eller karamelliserad produkt. 2. Tomatsaft och tomatkoncentrat skall vara
3. De krav som fastställs i punkt 2 skall anses vara uppfyllda om
4. Tomatsaft och tomatkoncentrat skall ha
c) en total titrerbar surhet, uttryckt som kristalliserad citronsyremonohydrat, på högst 10 viktprocent av torrsubstansinnehållet minskat med eventuell tillsats av vanligt salt,
5. Mögeltalet för tomatsaft och tomatkoncentrat skall, vid spädning med så mycket vatten att torrsubstanshalten uppgår till 8 %, inte överstiga 70 % positiva fält. För tomatsaft med en torrsubstanshalt på mindre än 8 %, skall procenttalet för positiva fält minskas i proportion till torrsubstanshalten.
Artikel 12
b) ha en god smak som är karakteristisk för en korrekt bearbetad produkt, och
3. Det sammanlagda innehållet av oorganiska och vegetabiliska orenheter får inte överstiga 1 % av produktens vikt. Med "vegetabiliska orenheter" avses här ett material av vegetabiliskt ursprung som kan urskiljas med blotta ögat och som inte är en del av själva tomaten eller som har suttit fast vid den färska tomaten men skulle ha avlägsnats vid bearbetningen, särskilt blad, stjälkar och foderblad från tomatplantan.
1. Behållare med konserverade skalade tomater, hela eller i bitar, och tomatsaft skall märkas med en referens som anger tillverkningsdatum och -år samt bearbetningsföretag. Om tomatsaft som har producerats på olika dagar har lagrats tillsammans innan den förpackas skall märkningen göra det möjligt att fastställa alla tillverkningsdagarna.
Artikel 14
a) torrsubstansinnehållet,
d) sockerinnehållet,
g) innehållet av oorganiska orenheter,
3. De metoder som avses i punkterna 1 och 2 skall användas för att slutgiltigt fastställa om produktionsstöd skall beviljas. Andra metoder får användas för rutinmässiga analyser.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Dessutom utesluter artikel 9.2 i fördraget varje administrativt förfarande som är avsett att skapa olika regler för rörelse av varor, beroende på om varorna har sitt ursprung i gemenskapen eller i tredje land och har övergått till fri omsättning i någon av medlemsstaterna.
Att en gemensam handelspolitik ännu inte helt genomförts innebär att det fortfarande kommer att finnas skillnader mellan medlemsstaterna i fråga om handelspolitiken, vilket kan vålla störning i handeln, något som artikel 115 i fördraget är avsedd att hindra.
Med hänsyn till erfarenheterna och det åtgärdsprogram gemenskapen har fastställt för genomförandet av den enhetliga marknaden bör beslut 80/47/EEG ändras. I synnerhet bör dess räckvidd utsträckas till alla de fall där det kvarstår skillnader inom de handelspolitiska åtgärder som har vidtagits av medlemsstater i enlighet med fördraget, däribland fall där skillnader inom tulltaxebestämmelser fortfarande tillåts, och vissa av de i beslutet angivna kriterierna och förfarandena bör specificeras. För att inarbeta dessa ändringar bör beslutet omarbetas till en enda rättsakt.
De uppgifter och de grunder som medlemsstaterna åberopar till stöd för en begäran om tillstånd för åtgärderna i fråga måste vara av sådan beskaffenhet att kommissionen fullt ut kan bedöma behovet av ett sådant tillstånd.
För att handeln mellan medlemsstaterna inte skall hindras, bör det föreskrivas att medlemsstaterna som regel bara skall begära vissa uppgifter från importören som ett led i uppfyllandet av formaliteterna vid import av en vara från en annan medlemsstat. Vad beträffar kontroll av ursprung skall medlemsstaterna i regel bara begära en enkel ursprungsdeklaration för varan, eftersom importören rimligen kan antas känna till ursprunget.
Räckvidd
Övervakning inom gemenskapen
a) det inte har skett betydande import av den ifrågavarande varan från andra medlemsstater under kalenderåret före det år då ansökan görs,
4. För att erhålla det tillstånd som avses i punkt 1 skall medlemsstaten lämna följande uppgifter i sin ansökan till kommissionen:
c) Den volym eller den mängd av varan som har sitt ursprung
- inom gemenskapen.
5. En medlemsstat som har fått det tillstånd som avses i punkt 1 får av den som ansöker om importhandling bara begära följande uppgifter:
c) En beskrivning av varan med uppgift om
d) Varans värde och kvantitet i de enheter som vanligen används i handeln.
Artikel 3
2. Kommissionen skall bevilja tillståndet bara för en begränsad period och bara när lägets allvar så kräver.
b) Den dag då ansökan om importhandling lämnades in.
- när den har sitt ursprung i andra tredje länder gentemot vilka den ansökande medlemsstaten til lämpar liknande importregler eller regler med motsvarande verkan,
d) Där så är möjligt, den volym eller den mängd av varan med ursprung i tredje landet i fråga som återexporteras till andra medlemsstater och till tredje land.
De uppgifter som begärs enligt punkterna c-e skall omfatta de två närmast föregående åren och det aktuella året.
- Medlemsstaten får avslå ansökan om en importhandling om kommissionens beslut tillåter detta.
Artikel 4
Artikel 5
1. Detta beslut skall tillämpas från och med den 1 oktober 1987.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av kommissionens förslag(1),
För att undanröja risken för missförstånd på grund av ordalydelsen i vissa artiklar i nämnda direktiv, är det nödvändigt att införa mindre rättelser.
För att minska antalet dokument som nu cirkulerar mellan medlemsstaterna bör ett typgodkännandeintyg, antingen i enlighet med det tillämpliga särdirektivet eller med förebilden i direktiv 70/156/EEG, anses uppfylla medlemsstaternas normala informationskrav. Medlemsstaterna har dock rätt att begära utförligare tekniska upplysningar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
I detta direktiv avses med:
- komponent: en anordning för vilken det fastställs krav i ett särdirektiv, som är avsedd att vara en del av ett fordon och som kan vara typgodkänd oberoende av ett fordon.
a) nationellt typgodkännande ett administrativt förfarande som benämns:
- "allgemeine Betriebserlaubnis" i tysk lagstiftning,
- "réception par type" i fransk lagstiftning,
- "agrément" i luxemburgsk lagstiftning,
- "type approval" i brittisk lagstiftning.
"Artikel 4
b) Fordonstypen måste uppfylla de kontrollkrav som anges i den förebild för typgodkännandeintyg som avses i artikel 2 b.
4. Varje medlemsstat skall fylla i alla avsnitt av ett typgodkännandeintyg för varje fordonstyp som den godkänner.
2. Medlemsstater har dock rätt att från en medlemsstat som har utfärdat typgodkännandet, eller från tillverkaren eller dennes representant, begära ytterligare sådana upplysningar som anges i de tekniska dokumenten i typgodkännandeintyget.
"2. Ett sådant intyg får dock inte hindra en medlemsstat från att vidta sådana åtgärder mot fordon som inte överensstämmer med den godkända typen.
"Artikel 8
3. De behöriga myndigheterna i medlemsstaterna skall inom en månad upplysa varandra om varje återkallat EEG-typgodkännande, och orsakerna till en sådan åtgärd.
6. Artikel 9a skall ändras enligt följande:
2. När den särskilda tekniska enheten eller komponenten som skall godkännas fyller sin funktion eller erbjuder en särskild egenskap endast tillsammans med andra fordonskomponenter och dess överensstämmelse med ett eller flera krav av denna anledning endast kan visas när den tekniska enheten eller komponenten som skall godkännas används tillsammans med andra fordonskomponenter, antingen på verkliga eller simulerade, måste omfattningen av EEG-typgodkännandet för den tekniska enheten eller komponenten begränsas i motsvarande grad. EEG-typgodkännandeintyget för en särskild teknisk enhet eller komponent skall i detta fall innehålla uppgifter om begränsning av dess användning och skall utvisa varje villkor för dess montering. Efterlevnaden av dessa begränsningar och villkor skall kontrolleras då fordonet EEG-typgodkänns.
7. Det tredje indraget i artikel 10.1 skall ersättas med följande:
De dokument som anges i bilagan till detta direktiv skall anses likvärdiga med de typgodkännandeintyg, vilka nämns i det tredje indraget i artikel 10.1 i direktiv 70/156/EEG.
2. Medlemsstaterna skall se till att kommissionen tillställs texten till de viktigaste bestämmelser i den nationella lagstiftningen som de antar inom det område som omfattas av detta direktiv.
med beaktande av rådets direktiv 79/117/EEG av den 21 december 1978 om förbud mot att växtskyddsprodukter som innehåller vissa verksamma ämnen släpps ut på marknaden och används(), särskilt artikel 6 i detta, senast ändrat genom direktiv 87/181/EEG(), och
Samtliga medlemsstater har meddelat kommissionen att de inte kommer att eller inte längre avser att utnyttja dessa undantag.
b) under 5, "Alkoxyalkyl- och arylkvicksilverföreningar", skall texten i andra kolumnen ersättas med: "Behandling av utsäde till spannmål och betor".
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: I artikel 13 i förordning (EEG) nr 2261/84(3), senast ändrad genom förordning (EEG) nr 3788/85(4), föreskrivs att tillfälligt godkännande får beviljas för fabriker som lämnar in en ansökan om godkännande under regleringssåren 1984/85 och 1985/86. Erfarenheten har visat att de berörda medlemsstaterna inte är i stånd att genomföra de kontroller som behövs inom den fastställda tiden. Dessa tider bör därför förlängas.
Artikel 1
Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag, och
Lämpliga åtgärder skall vidtas för att genomföra det nya systemet med intyg inom gemenskapen och för att se till att det tillämpas utan att några importörer i gemenskapen missgynnas.
Export från gemenskapen av kaffe och extrakt, essenser eller koncentrat av kaffe enligt undernummer 09.01 A och 21.02 A i Gemensamma tulltaxan skall inte vara beroende av inlämnande av de intyg som föreskrivs i avtalet.
med beaktande av rådets förordning (EEG) nr 3094/86 av den 7 oktober 1986 om vissa tekniska åtgärder för bevarande av fiskeresurserna(), ändrad genom förordning (EEG) nr 4026/86(), särskilt artikel 15 i denna, och med beaktande av följande:
Om en förstärkande nätkasse med mindre maskstorlek användes skulle dessa problem kunna undvikas utan negativ inverkan på fiskebeståndet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 5.5 skall ersättas med följande:
- Punkt 2 skall ersättas med följande:
"3. Maskstorleken skall vara minst dubbelt så stor som lyftets. Om en andra förstärkande nätkasse används skall den ha en maskstorlek på minst 120 mm."
- Punkt 7 skall ersättas med följande:
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 1
Artikel 1 i kommissionens förordning nr 183/66/EEG av den 18 november 1966 om icke-fastställande av en tilläggsavgift för sydafrikanska ägg () skall ersättas med följande: "Artikel 1 I enlighet med artikel 8.2 i förordning (EEG) nr 2771/75 skall de importavgifter som fastställts i enlighet med artikel 3 i samma förordning inte höjas med en tilläggsavgift i samband med import av ägg med skal (undernummer 0407 00 i Kombinerade nomenklaturen) som har sitt ursprung i och kommer från Sydafrika."
Artikel 4
1. Artikel 1 skall ersättas med följande: "Artikel 1 Importavgifter som fastställs i enlighet med artikel 3 i förordning (EEG) nr 2771/75 skall inte höjas med en tilläggsavgift i samband med import av produkter som omfattas av följande nummer i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Österrike: >Plats för tabell>
Artikel 1 i kommissionens förordning (EEG) nr 59/70 av den 14 januari 1970 om ickefastställande av tilläggsavgifter för ägg med skal som importeras från Rumänien () skall ersättas med följande: "Artikel 1 Importavgifter som fastställts i enlighet med artikel 3 i förordning (EEG) nr 2771/75 skall inte höjas med en tilläggsavgift i samband med import av fjäderfäägg med skal, färska eller konserverade, undantaget kläckägg, som omfattas av undernummer 0407 00 30 i Kombinerade nomenklaturen och som har sitt ursprung i och kommer från Rumänien."
Artikel 8
KOMMISSIONENS BESLUT av den 28 oktober 1988 om upprättande av en förteckning över produkter som avses i artikel 3.1 andra stycket i rådets förordning (EEG) nr 1898/87 (88/566/EEG)
Artikel 1 De produkter inom gemenskapens territorium som motsvarar de produkter som avses i artikel 3.1 andra stycket i förordning (EEG) nr 1898/87 upptas i förteckningen i bilagan.
med beaktande av följande: Med hänsyn till vunna erfarenheter och teknikens nuvarande utvecklingsnivå är det nu möjligt att skärpa vissa krav i direktiv 71/127/EEG i syfte att förbättra trafiksäkerheten.
De i detta direktiv fastställda åtgärderna har tillstyrkts av Kommittén för anpassning till teknisk utveckling av direktiv om avskaffande av tekniska handelshinder inom motorfordonssektorn.
Bilagorna 2 och 3 till direktiv 71/127/EEG ändras härigenom i enlighet med bilagan till detta direktiv.
- vare sig vägra att bevilja EEG-typgodkännande eller att utfärda dokumentet enligt artikel 10.1. tredje strecksatsen i rådets direktiv 70/156/EEG(3), eller att bevilja nationellt typgodkännande,
2. Från och med den 1 oktober 1990 gäller följande:
- De får förbjuda att fordon, vars backspeglar inte överensstämmer med bestämmelserna i detta direktiv tas i bruk.
Artikel 4
med beaktande av kommissionens förslag,
För den juridiska klarhetens skull bör ordalydelsen av artikel 11.2 i direktiv 83/181/EEG preciseras.
Direktiv 83/181/EEG ändras på följande sätt:
2. Artikel 22 skall ersättas med följande:
4. Följande kapitel införs efter artikel 38:
Artikel 38 a
"d) Priser, troféer och souvenirer av symbolisk natur och med begränsat värde, avsedda för gratisutdelning till personer som normalt är bosatta i ett annat land än införsellandet vid affärskonferenser eller liknande internationella evenemang, och vars beskaffenhet, värde per styck eller övriga kännetecken inte är sådana att de skulle kunna vara avsedda för kommersiella ändamål."
Med förbehåll för vad som föreskrivs i artikel 63 skall tryckt reklammaterial såsom kataloger, prislistor, bruksanvisningar eller broschyrer vara skattebefriade vid införsel, om de hänför sig till:
c) transport-, handels-, försäkrings- eller banktjänster som erbjuds av en person som är etablerad i ett tredje land.
a) Trycksakerna måste tydligt utvisa namnet på det företag som producerar, säljer eller hyr ut de varor eller som erbjuder de tjänster till vilka de hänför sig.
Villkoren i punkterna b och c skall dock inte tillämpas på trycksaker som avser antingen varor till salu eller uthyrning eller tjänster som erbjuds av en person som är etablerad i en annan medlemsstat, om trycksakerna har införts och kommer att distribueras gratis."
8. Titeln på kapitel VI skall ersättas med följande:
- specialcontainrar,
a) kommersiella motorfordon: motordrivna vägfordon (även traktor med släpvagn) som genom sin konstruktionstyp och utrustning är utformade för och ägnade att transportera, mot eller utan betalning: - mer än nio personer inräknat föraren,
b) privata motorfordon: motorfordon som inte omfattas av definitionen i punkt a.
10. Första punkten i artikel 83 ändras på följande sätt:
"c) till 200 liter per specialcontainer och resa."
Artikel 2
Detta direktiv riktar sig till medlemsstaterna.
Dessa kvalitativa kännetecken bör motsvara de egenskaper som konstateras för sorter som importeras från områden där indicaris traditionellt odlas.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
1. Från och med regleringsåret 1988/89 skall endast de rissorter förtecknas i bilaga B till förordning (EEG) nr 3878/87 som har de morfologiska kännetecken som anges i artikel 2.1 i förordningen och följande kvalitativa kännetecken:
- Ett amylosinnehåll på minst 21 %.
1. Det laboratorium som ansvarar för bearbetningen av riset, skall efter att ha genomfört grobarhetsprov och bearbetat riset, översända prover märkta med en kod till samtliga laboratorier som förtecknas i bilaga 2 samt översända ett förseglat meddelande som möjliggör avkodning av proverna till kommissionens tjänstemän.
1. Kommissionens personal skall bestämma de aktuella sorternas kännetecken på grundval av det aritmetiska medelvärdet av analysresultaten, sedan det högsta och det lägsta värdet uteslutits.
Artikel 5
med beaktande av följande: För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser angående klassificering av de varor som anges i bilagan till den här förordningen.
Nomenklaturkommittén har inte yttrat sig över förslaget inom den tid som ordföranden bestämt.
De varor som beskrivs i kolumn 1 i tabellen i bilagan klassificeras nu inom Kombinerade nomenklaturen enligt de tillämpliga KN-nummer som anges i kolumn 2 i denna tabell.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av följande: Enligt artikel 1.1 i förordning (EEG) nr 2262/84(3), senast ändrad genom förordning (EEG) nr 3462/87(4), skall de producerande medlemsstaterna upprätta organ som skall utföra vissa kontroller och uppgifter i samband med programmet för produktionsstöd för olivolja. Enligt artikel 1.5 i den förordningen skall rådet före den 1 januari 1989 fastställa metoden för finansiering av organens utgifter från och med regleringsåret 1989/90.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"5. Under en tid av fem år från och med den 1 november 1984 skall följande procentsatser av organets faktiska utgifter debiteras de europeiska gemenskapernas allmänna budget:
Under en tid av tre år från och med den 1 november 1989 skall 50 % av de faktiska utgifterna för organen i Italien och Grekland belasta de europeiska gemenskapernas allmänna budget.
Rådet skall med kvalificerad majoritet på förslag från kommissionen senast den 1 januari 1992 fastställa metoden för finansiering av utgifterna i fråga från och med regleringsåret 1992/93."
RÅDETS DIREKTIV av den 12 juni 1989 om åtgärder för att främja förbättringar av arbetstagarnas säkerhet och hälsa i arbetet (89/391/EEG)
med beaktande av kommissionens förslag(1), utarbetat efter samråd med Rådgivande kommittén för arbetarskyddsfrågor,
med beaktande av följande: Enligt artikel 118a i fördraget skall rådet genom direktiv fastställa minimikrav i syfte att främja förbättringar, framför allt på arbetsmiljöområdet, för att trygga en högre skyddsnivå för arbetstagarnas säkerhet och hälsa.
Rådet uppmärksammade i sin resolution av den 21 december 1987 om arbetarskyddsfrågor(5) att kommissionen avsåg att inom en snar framtid föreslå rådet ett direktiv om organisationen av verksamheten för arbetstagarnas säkerhet och hälsa på arbetsplatsen.
Medlemsstaternas arbetarskyddslagstiftning varierar avsevärt och behöver förbättras; nationella bestämmelser, som ofta innehåller tekniska föreskrifter och/eller vägledande normer, kan leda till skilda skyddsnivåer och möjliggöra konkurrens på bekostnad av säkerhet och hälsa.
Information, dialog och avvägd medverkan i frågor som rör säkerhet och hälsa i arbetet måste utvecklas mellan arbetsgivare och arbetstagare och/eller deras representanter med hjälp av ändamålsenliga metoder och medel i överensstämmelse med nationell lagstiftning och/eller praxis.
Utan att det inskränker strängare existerande eller framtida gemenskapsbestämmelser skall detta direktiv tillämpas på alla risker och i synnerhet på dem som härrör från hanteringen av de kemiska, fysiologiska och biologiska agenser, som omfattas av direktiv 80/1107/EEG(6), senast ändrat genom direktiv 88/642/EEG(7).
2. För det ändamålet innehåller direktivet dels allmänna principer för att förebygga yrkesbetingade risker, för arbetarskydd, för att eliminera riskfaktorer och faktorer, som kan förorsaka olycksfall, för information, samråd, avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis samt utbildning av arbetstagarna och deras representanter, dels allmänna riktlinjer för genomförandet av dessa principer.
Räckvidd
I dessa fall skall arbetstagarnas säkerhet och hälsa tryggas så långt möjligt mot bakgrund av direktivets syften.
I detta direktiv avses med
c) arbetstagarrepresentanter med särskilt ansvar för arbetstagarnas säkerhet och hälsa, varje person, som i enlighet med nationell lagstiftning och/eller praxis har utsetts, valts eller utnämnts att representera arbetstagarna i arbetarskyddsfrågor,
1. Medlemsstaterna skall vidta tillräckliga åtgärder för att säkerställa att arbetsgivare, arbetstagare och arbetstagarrepresentanter omfattas av sådana lagar och andra författningar som behövs för att bestämmelserna i detta direktiv skall kunna genomföras i praktiken.
Artikel 5
2. I de fall en arbetsgivare i överensstämmelse med artikel 7.3 anlitar tjänster eller personer utifrån skall han inte fritas från sitt ansvar på detta område.
Arbetsgivarens allmänna skyldigheter
2. Arbetsgivaren skall verkställa de åtgärder som avses i punkt 1 första stycket med utgångspunkt från följande allmänna principer för förebyggande arbete:
Som en följd av denna utvärdering, skall vid behov de förebyggande åtgärder samt de arbets- och produktionsmetoder, som tillämpas av arbetsgivaren
b) Då arbetsgivaren uppdrar åt arbetstagaren att utföra vissa arbetsuppgifter skall han ta hänsyn till dennes kunskaper på arbetarskyddsområdet.
4. Utan att det inskränker övriga bestämmelser i detta direktiv skall arbetsgivare, där flera företag samtidigt driver verksamhet på ett arbetsställe, samverka vid tillämpningen av reglerna om säkerhet, hälsa och arbetshygien samt, med beaktande av verksamhetens art, samordna sina åtgärder i skyddshänseende och i frågor som rör förebyggande av risker i arbetet samt underrätta varandra och sina respektive arbetstagare och/eller arbetstagarrepresentanter om dessa risker.
Skydds- och förebyggande åtgärder
De utsedda arbetstagarna skall ges skälig tid för att kunna fullgöra sina skyldigheter enligt detta direktiv.
- de utsedda arbetstagarna ha tillräckliga kunskaper och resurser,
Arbetstagaren/arbetstagarna och/eller enheten/enheterna skall vid behov samarbeta.
De kan fastställa det erforderliga antal, som åsyftas i punkt 5.
1. Arbetsgivaren skall
Dessa arbetstagare skall vara tillräckligt många, de skall erhålla fullgod utbildning och ha tillgång till ändamålsenlig utrustning med beaktande av företagets och/eller verksamhetens storlek och särskilda risker.
b) vidta åtgärder och ge anvisningar så att alla arbetstagare i händelse av allvarlig, överhängande och oundviklig fara kan avbryta arbetet och/eller omedelbart avlägsna sig från sin arbetsplats och sätta sig i säkerhet,
5. Arbetsgivaren skall säkerställa att alla arbetstagare, i fall då en allvarlig och överhängande fara för arbetstagarnas och/eller andras säkerhet föreligger, och då den närmast ansvariga arbetsledningen inte kan kontaktas, kan vidta lämpliga åtgärder med hänsyn till sin kunskap och de tekniska resurser, som står till deras förfogande, för att avvärja en sådan fara.
Arbetsgivarens skyldigheter i övrigt
b) besluta om de skyddsåtgärder som skall vidtas och den eventuella personliga skyddsutrustning som skall användas,
2. Medlemsstaterna skall fastställa, med hänsyn till verksamhetens art och företagens storlek, de skyldigheter som åvilar skilda grupper av företag i fråga om upprättande av de handlingar som avses i punkt 1 a och b och vid utarbetande av handlingar enligt punkt 1 c och d.
1. I enlighet med nationell lagstiftning och/eller praxis som kan ta hänsyn till bland annat företagets/verksamhetens storlek skall arbetsgivaren vidta lämpliga åtgärder så att arbetstagare och /eller deras representanter i företaget och/eller verksamheten får all den information som behövs om
2. Arbetsgivaren skall vidta lämpliga åtgärder så att arbetsgivare för anställda i utomstående företag och/eller verksamheter, vilka utför arbete i den förstnämndes företag och/eller verksamhet, i enlighet med nationell lagstiftning och/eller praxis, får den information om förhållandena enligt punkterna 1 a och b som skall lämnas arbetstagarna ifråga.
b) det register och de rapporter som åsyftas i artikel 9.1 c och d,
Samråd med och medverkan av arbetstagare
- överläggningar med arbetstagarna,
2. Arbetstagare eller arbetstagarrepresentanter med särskilt ansvar för skyddsfrågor skall ges rätt till avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis, eller rådfrågas i förväg och i god tid beträffande
c) den information som åsyftas i artiklarna 9.1 och 10,
3. Arbetstagarrepresentanter med särskilt ansvar för skyddsfrågor skall ha rätt att anmoda arbetsgivaren att vidta lämpliga åtgärder och lägga fram förslag i syfte att minska riskerna för arbetstagarna och/eller undanröja källan till faran.
Arbetstagarrepresentanter skall ges tillfälle att lägga fram sina iakttagelser i samband med inspektionsbesök av den behöriga myndigheten.
1. Arbetsgivaren skall säkerställa att varje arbetstagare får tillräcklig utbildning i arbetsmiljöfrågor, framför allt i form av information och instruktioner, som har direkt anknytning till platsen där han arbetar eller hans arbetsuppgifter i samband med
- införande av ny arbetsutrustning eller ändring av arbetsutrustning,
- anpassas till nya eller ändrade risksituationer, och
3. Arbetstagarrepresentanter med särskilda uppgifter i skyddsfrågor skall ha rätt till tillräcklig utbildning.
Den utbildning som avses i punkt 3 skall förläggas till arbetstid och i enlighet med nationell praxis äga rum inom eller utanför företaget och/eller verksamheten.
1. Det åligger varje arbetstagare att så långt möjligt sörja för sin egen och andra personers säkerhet och hälsa, i den mån de påverkas av hans handlingar eller förtroendeuppdrag i arbetet, i enlighet med hans utbildning och arbetsgivarens instruktioner.
1. Åtgärder skall vidtas i enlighet med nationell lagstiftning och/eller praxis i syfte att tillförsäkra arbetstagarna hälsokontroller anpassade till de arbetsmiljörisker, som de utsätts för i arbetet.
Artikel 15
Artikel 16
3. Bestämmelserna i detta direktiv skall fullt ut tillämpas på alla områden, som omfattas av särdirektiven utan att hindra tillämpningen av de strängare eller mer specifika bestämmelser som finns i särdirektiven.
1. När rent tekniska justeringar av de särdirektiv som föreskrivs i artikel 16.1 görs för att ta hänsyn till
skall kommissionen biträdas av en kommitté bestående av företrädare för medlemsstaterna och med en företrädare för kommissionen som ordförande.
Beslut om yttrandet skall fattas med tillämpning av de omröstningsregler som enligt fördragets artikel 148.2 gäller för beslut som rådet skall fatta på förslag av kommissionen.
Om förslaget inte har tillstyrkts av kommittén eller om den inte avger något yttrande, skall kommissionen utan dröjsmål föreslå rådet åtgärder. Rådet skall besluta med kvalificerad majoritet.
Slutbestämmelser
Kommissionen skall informera Europaparlamentet, rådet, Ekonomiska och sociala kommittén och Rådgivande kommittén för arbetarskyddsfrågor.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Europaparlamentets yttrande(),
Det är nödvändigt att i möjligaste mån underlätta den fria rörligheten för personer inom gemenskapen.
Artikel 1
"b) som personen i fråga faktiskt har haft i bruk innan bytet av hemvist genomfördes eller andrabostaden inrättades. I fråga om motorfordon (inklusive tillhörande släpvagnar), husvagnar och husbilar, nöjesbåtar och privatflygplan, får medlemsstaterna kräva att den flyttande har haft dem i bruk minst sex månader före bytet av hemvist.
3. Artikel 5.1 skall ersättas med följande:
b) I punkt 1 skall följande stycke tillfogas:
b) Tredje stycket skall utgå.
"1. Utan att det påverkar tillämpningen av artiklarna 2 5, skall var och en vid giftermål vara berättigad till befrielse från de skatter som avses i artikel 1 när han till den medlemsstat dit han avser att flytta inför personlig egendom som han förvärvat eller har haft i bruk, förutsatt att".
7. I artikel 11 görs följande ändringar:
Artikel 3
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(2),
För att samordningen av marknaden med kreatursprodukter och produkter av animaliskt ursprung skall fungera utan störningar krävs att veterinära hinder mot utvecklingen av handeln inom gemenskapen med dessa produkter undanröjs. Den fria rörligheten av jordbruksprodukter är ett grundläggande inslag i samordningen av marknaderna och bör kunna underlätta en rationell utveckling av jordbruksproduktionen och ett optimalt utnyttjande av produktionsmedlen.
Målet är att förverkliga den inre marknaden och i avvaktan på att detta uppnås bör huvudvikten läggas på de kontroller som skall utföras hos avsändaren och på att organisera de kontroller som skulle kunna utföras på destinationsorten. En sådan lösning skulle innebära ett slopande av de veterinära kontrollerna vid gränserna mellan medlemsstaterna.
Det är en uppgift för medlemsstaterna att lägga fram en plan över hur de avser att utföra kontrollerna. Dessa planer bör underställas gemenskapen för godkännande.
För att vara effektiva måste de regler som fastställs i detta direktiv täcka alla varor som är underkastade veterinära krav i samband med handel inom gemenskapen.
Dessa regler bör ses över på nytt före utgången av år 1993.
Artikel 1
I detta direktiv avses med
3. anläggning: varje företag som producerar, lagrar eller bearbetar produkter som avses i artikel 1,
Artikel 3
Utan att påverka de tillsynsskyldigheter som åligger den officiella veterinären i enlighet med gemenskapens lagstiftning skall den behöriga myndigheten utföra regelbunden kontroll vid anläggningarna för att försäkra sig om att de för handel avsedda produkterna uppfyller gemenskapens krav eller, i de fall som avses under punkt 3 i denna artikel och i artikel 14, de krav som gäller i den mottagande medlemsstaten.
När de produkter som åsyftas i artikel 1 är avsedda för export till ett tredje land skall transportproceduren stå under tullövervakning fram till den ort där sändningen lämnar gemenskapens territorium.
De medlemsstater till vilka varorna är destinerade skall förbjuda att de berörda produkterna sänds vidare från deras territorium såvida de inte är avsedda för någon annan medlemsstat som begagnar sig av samma införselmöjlighet.
- de produkter som anskaffats i enlighet med de direktiv som avses i bilaga A kontrolleras på samma sätt ur veterinär synpunkt, oavsett om de är avsedda för handel inom gemenskapen eller för den inhemska marknaden.
1. Mottagande medlemsstater skall vidta följande åtgärder:
b) När de produkter som avses i artikel 1 och som härrör från en annan medlemsstat är avsedda
- för andra mottagare, särskilt när partiet till en del har lossats under transporten, skall förpackningen i enlighet med artikel 3.1 åtföljas av originalet till det intyg som avses i den första strecksatsen.
3. För importörer som får produkter levererade till sig från en annan medlemsstat eller som helt delar upp ett parti av sådana produkter gäller att
c) de skall, om den behöriga myndigheten kräver detta, anmäla ankomsten av sådana produkter från en annan medlemsstat i den mån detta är nödvändigt för att utföra de kontroller som avses under punkt 1,
5. Rådet skall med ledning av en rapport från kommissionen som åtföljs av eventuella ändringsförslag på nytt se över denna artikel inom tre år från det att detta direktiv börjar tillämpas.
a) Kontroller av handlingar skall göras rörande produkternas ursprung.
De produkter som avses i bilaga B och de varor som medlemsstaterna har valt att importera i enlighet med artikel 3.3 och som efter att ha införts till gemenskapens territorium skall vidarebefordras till en annan medlemsstats territorium skall
c) Produkter som härrör från gemenskapen skall inspekteras i enlighet med de besiktningsbestämmelser som fastställs i artikel 5.
1. Om den behöriga myndigheten i en medlemsstat i samband med den inspektion som utförs på destinationsorten eller under transporten konstaterar
De behöriga myndigheterna i den mottagande medlemsstaten skall omedelbart genom telex delge de övriga medlemsstaternas behöriga myndigheter och kommissionen vad som framkommit vid inspektionen, vilka beslut som fattats och på vilka grunder de fattats.
b) att varorna inte uppfyller de villkor som fastställts genom gemenskapens direktiv, eller nationella normer när ett beslut om de gemenskapsnormer som föreskrivits genom direktiven inte fattats, och förutsatt att hänsynen till människors och djurs hälsa tillåter det, låta avsändaren eller hans ombud välja mellan att
Om intyget eller dokumenten befinns innehålla felaktigheter skall dock avsändaren medges en tidsfrist innan den sistnämnda möjligheten tillgrips.
1. I de fall som avses i artikel 7 skall den behöriga myndigheten i den mottagande medlemsstaten utan dröjsmål ta kontakt med de behöriga myndigheterna i den medlemsstat från vilken varorna avsänts. De sistnämnda myndigheterna skall vidta alla nödvändiga åtgärder och meddela den behöriga myndigheten i den förstnämnda medlemsstaten vilka kontroller som utförts, vilka beslut som fattats och motiveringen för dessa.
Kommissionen får på begäran av den behöriga myndigheten i den mottagande medlemsstaten eller på eget initiativ och under hänsynstagande till arten av överträdelsen
- uppmana den behöriga myndigheten att intensifiera provtagningen av den berörda anläggningens produkter.
I avvaktan på vad kommissionen kommit fram till skall den medlemsstat från vilken sändningen härrör, på begäran av den mottagande medlemsstaten, utöka kontrollen av de produkter som kommer från den ifrågavarande anläggningen och tillfälligt dra in tillståndet om det föreligger starka skäl för detta med hänsyn till djurs och människors hälsa.
De allmänna reglerna för tillämpningen av denna artikel skall fastställas i enlighet med förfarandet i artikel 18.
Om avsändaren eller hans ombud begär detta, skall de ifrågavarande besluten tillsammans med motivering vidarebefordras till honom i skriftlig form med uppgifter om den rätt till prövning som står till buds i enlighet med gällande lagstiftning i den mottagande medlemsstaten, tillsammans med uppgift om hur och inom vilken tid detta skall ske.
3. Kostnaderna för att sända tillbaka varorna, lagra dem, överföra dem till annan användning eller förstöra dem skall betalas av mottagaren.
Den mottagande medlemsstaten eller den genom vilken sändningen skall transiteras, som i samband med någon av de kontroller som avses i artikel 5 har konstaterat förekomst av någon av de sjukdomar eller orsaker som avses i första stycket, får om så krävs vidta de försiktighetsmått som fastställs i gemenskapens regler.
2. På begäran av den medlemsstat som avses i första stycket i punkt 1, eller på initiativ av kommissionen, får en eller flera kommissionsledamöter omedelbart bege sig till den berörda platsen för att i samarbete med de behöriga myndigheterna undersöka vilka åtgärder som vidtagits. De skall avge ett yttrande om dessa åtgärder.
5. Utförliga regler för hur denna artikel skall tillämpas och särskilt förteckningen över de zoonoser eller orsaker som kan tänkas utgöra ett allvarlig hot mot människors hälsa skall utarbetas i enlighet med förfarandet i artikel 18.
Artikel 11
- kontrollera att personalen uppfyller de krav som fastställs i de texter som avses i bilaga A,
För detta ändamål skall de inspekterade anläggningarna vara beredda att samarbeta med kontrollanterna i den utsträckning som krävs för att de skall kunna fullgöra sina åligganden.
2. Artikel 5.3 och 5.4 och artiklarna 9, 10 och 11 i direktiv 71/118/EEG(10), senast ändrat genom direktiv 88/657/EEG, utgår.
ii) i artikel 8a skall hänvisningen till artikel 8 ersättas med en hänvisning till artikel 9 i direktiv 89/662/EEG.
i) skall artikel 5.2, 5.3, 5.4 och 5.5 och artiklarna 6 och 7 utgå, och
7. Artikel 10.1 och 10.3 i direktiv 88/657/EEG utgår.
Artikel 13
2. Följande artikel skall läggas till direktiven 72/461/EEG och 80/215/EEG:
"Artikel 24
5. Följande artikel läggs till direktiv 88/437/EEG:
Fram till och med den 31 december 1992 skall, i avvaktan på beslut om att gemenskapsregler skall antas, handeln med de produkter som räknas upp i bilaga B vara underkastade de regler om kontroll som fastställs i detta direktiv, särskilt de som fastställs i artikel 5.2.
Artikel 15
Artikel 16
3. Varje år från och med 1991 skall kommissionen till medlemsstaterna överlämna en rekommendation till program för kontroller att genomföras påföljande år. Den ständiga veterinärkommittén skall i förväg ha avgivit sitt yttrande om rekommendationen som får bli föremål för senare anpassningar.
4. Om förslaget inte är förenligt med yttrandet från kommittén eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas.
Artikel 18
3. Kommissionen skall godkänna de tilltänkta åtgärderna om de är förenliga med kommitténs yttrande.
Artikel 19
2. Före den 31 december 1992 skall rådet se över bestämmelserna i detta direktiv och med ledning av en rapport från kommissionen om de erfarenheter som vunnits, tillsammans med relevanta förslag, fatta beslut om dessa med kvalificerad majoritet.
- upprätthålla kontroller av handlingar under transporten av kött och produkter som härrör från kött för att säkerställa att de speciella krav rörande mul- och klövsjuka och svinpest som fastställs genom gemenskapsregler uppfylls,
Rådet skall före den 1 oktober 1992, med kvalificerad majoritet efter förslag från kommissionen, bestämma vilka arrangemang som skall tillämpas när de övergångsbestämmelser som fastställs i artikel 20 upphör att gälla.
Dock skall Grekland ges en ytterligare ett års respit med att följa det.
RÅDETS DIREKTIV av den 21 december 1989 om samordning av lagar och andra författningar för prövning av offentlig upphandling av varor och bygg- och anläggningsarbeten (89/665/EEG)
med beaktande av kommissionens förslag (1),
med beaktande av följande: Gemenskapens direktiv om offentlig upphandling, särskilt rådets direktiv 71/305/EEG av den 26 juli 1971 för samordning av förfarandena vid tilldelning av bygg- och anläggningsarbeten (4), senast ändrat genom direktiv 89/440/EEG (5) och rådets direktiv 77/62/EEG av den 21 december 1976 om samordningar av förfarandet vid offentlig upphandling av varor (6), senast ändrat genom direktiv 88/295/EEG (7), innehåller ej bestämmelser som säkrar deras effektiva tillämpning.
Eftersom upphandlingsförfarandet för varje särskilt kontrakt är kortvarigt, måste ett sakkunnigt prövningsorgan bl.a. vara behörigt att vidta interimistiska åtgärder i syfte att uppskjuta förfarandet hos myndigheten eller verkställigheten av dess beslut. Med hänsyn till tidsfaktorn måste vidare ges möjlighet att snabbt ingripa mot nämnda överträdelser.
Följaktligen bör kommissionen ges behörighet att föra ärendet inför vederbörande myndigheter i medlemslandet såväl som upphandlingsmyndigheten, så snart den anser, att en klar och konkret överträdelse har begåtts vid upphandlingsförfarandet, så att lämpliga åtgärder vidtas för skyndsam rättelse av en påstådd kränkning.
Artikel 1
3. Medlemsstaterna skall se till att ett prövningsförfarande med detaljerade regler enligt medlemsstaternas bestämmande införs och att det kan åberopas av var och en, som har eller har haft intresse av att få avtal om viss offentlig upphandling av varor eller bygg- och anläggningsarbeten, och som har skadats eller riskerat att skadas av en påstådd överträdelse. Det förutses, att en medlemsstat skall kunna kräva av den person som begär prövning, att han dessförinnan meddelat den avtalsslutande myndigheten att han hävdar förekomsten av diskriminering, och att han ämnar söka prövning.
a) så tidigt som möjligt vidta interimistiska åtgärder för att rätta påstådda överträdelser eller förhindra ytterligare skada för berörda intressen, inklusive åtgärder för att uppskjuta eller garantera uppskjutandet av upphandlingsförfarandet liksom att förhindra verkställighet av den upphandlande myndighetens beslut,
2. Behörighet enligt punkt 1 får ges till separata organ med ansvar för olika sidor av prövningsförfarandet.
6. Verkan av att behörighet har utövats enligt punkt 1 på ett redan slutet avtal om upphandling skall regleras i nationell lag.
8. För de fall prövningsorganen ej utgörs av rättsliga instanser gäller, att skriftliga beslutsmotiveringar alltid skall ges. Dessutom gäller för dessa fall, att det måste finnas en möjlighet att pröva påstådda olagliga åtgärder vidtagna av sådana organ i en rättslig instans eller en domstol som avses i fördragets artikel 177, oberoende av såväl upphandlingsmyndigheten som prövningsorganet.
1. Kommissionen får tillgripa prövningsförfarandet enligt denna artikel, om den innan ett upphandlingskontrakt slutits anser, att en klar och konkret överträdelse av gemenskapsreglerna har ägt rum vid en offentlig upphandling inom områdena för direktiven 71/305/EEG och 77/62/EEG.
a) bekräftelse på att överträdelsen har rättats till,
4. En förklaring enligt punkt 3 b kan bl.a. vila på, att den påstådda överträdelsen redan är föremål för rättslig eller annan undersökning eller prövningsförfarande enligt artikel 2.8. I sådant fall måste medlemsstaten underrätta kommissionen om resultatet av detta, så snart det blir känt.
2. Medlemsstaterna skall årligen före den 1 mars rapportera till kommissionen om sin tillämpning av prövningsbestämmelserna under föregående kalenderår. Anvisningar om rapportens innehåll utarbetas av kommissionen i samråd med Rådgivande kommittén för offentlig upphandling.
Artikel 6
med beaktande av följande: För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser angående klassificering av de varor som anges i bilagan till den här förordningen.
Nomenklaturkommittén har inte yttrat sig över förslaget inom den tid som ordföranden bestämt.
De varor som beskrivs i kolumn 1 i tabellen i bilagan klassificeras nu inom Kombinerade nomenklaturen enligt de till- lämpliga KN-nummer som anges i kolumn 2 i denna tabell.
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom förordning (EEG) nr 20/89(2), särskilt artikel 9 i denna, och
Klädesplagg utan ärmar eller med korta ärmar ger inte detta skydd. Det är därför nödvändigt att ange att anoraker, vindjackor och liknande artiklar, som nämns ovan, måste ha långa ärmar.
Artikel 1
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av kommissionens förslag, som utformats efter yttrande av en grupp experter utsedda av Vetenskapliga och tekniska kommittén(1),
med beaktande av följande: Bilagan till förordning (Euratom) nr 3954/87(4) innehåller rubriker för gränsvärden för livsmedel och djurfoder.
Därför bör det göras tillägg till bilagan till förordningen.
Med hänsyn till det fortsatta arbetet bör det också föreskrivas att förfarandet i artikel 7 i förordning (Euratom) nr 3954/87 också tillämpas för att fastställa gränsvärden för djurfoder. Det bör därför göras lämpliga tillägg till förordningen.
Bilagan till förordning (Euratom) nr 3954/87 skall ersättas med bilagan till denna förordning.
"Artikel 7
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av följande: I enlighet med artikel 13 i direktiv 64/433/EEG och i enlighet med förfarandet i artikel 16 får på begäran undantag från punkt 45 c i bilaga 1 beviljas varje medlemsstat som lämnar liknande garantier. Vid sådana undantag skall hygienkrav som lägst motsvarar kraven i nämnda bilaga fastställas.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
I brev av den 18 januari 1989 har myndigheterna i Frankrike till kommissionen framfört en begäran om undantag från punkt 45 c i bilaga 1 till direktiv 64/433/EEG i fråga om styckning av färskt nötkött, fårkött och griskött. I begäran föreslås hygienkrav. Det är nödvändigt att de alternativa hygienkrav som fastställs i det begärda undantaget i fråga om styckning av färskt kött lägst motsvarar kraven i punkt 45 c i bilaga 1 till direktiv 64/433/EEG.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
I förordning (EEG) nr 2658/87 fastställs allmänna bestämmelser för tolkningen av Kombinerade nomenklaturen och dessa gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna, eller som lägger ytterligare underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser med tanke på tillämpningen av tulltaxebestämmelser eller andra bestämmelser som rör varuhandeln.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Nomenklaturkommittén vad gäller produkterna nr 1, 2, 3, 5 och 6 i tabellen i bilagan.
De varor som beskrivs i kolumn 1 i tabellen i bilagan klassificeras nu inom Kombinerade nomenklaturen enligt de tillämpliga KN-nummer som anges i kolumn 2 i denna tabell.
KOMMISSIONENS BESLUT av den 2 maj 1991 om erkännande av Australien som fritt från Erwinia amylovora (Burr.) Winsl. et al. (91/261/EEG)
med beaktande av rådets direktiv 77/93/EEG av den 21 december om skyddsåtgärder mot att skadegörare på växter eller växtprodukter förs in till medlemsstaterna(1), senast ändrat genom kommissionens direktiv 91/27/EEG(2), särskilt bilaga 3 del B 10 i detta, och med beaktande av följande:
Det kan därför fastslås att det inte finns någon risk för spridning av den ovan nämnda skadegöraren.
De åtgärder som föreskrivs i detta beslut är förenliga medyttrandet från Ständiga kommittén för växtskydd.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
Vissa medlemsstater har redan infört begränsningar i fråga om användning eller utsläppande på marknaden av dessa ämnen eller preparat i vilka de ingår. Åtgärderna inverkar direkt på den inre marknadens upprättande och funktion. En tillnärmning av medlemsstaternas lagstiftning på detta område är således nödvändig. Bilaga 1 till direktiv 76/769/EEG(4), senast ändrat genom direktiv 89/678/EEG(5), bör därför ändras.
RÅDETS DIREKTIV av den 16 december 1991 om det ömsesidiga erkännandet av båtförarcertifikat för transport av gods och passagerare på inre vattenvägar (91/672/EEG)
Vid tillämpningen av detta direktiv skall nationella båtförarcertifikat för transport av gods och passagerare på inre vattenvägar enligt bilaga 1 indelas på följande sätt:
Artikel 3
3. En medlemsstats erkännande av ett båtförarcertifikat enligt grupp A eller grupp B i bilaga 1 får underkastas samma villkor angående minimiålder som de villkor som fastställts i denna medlemsstat för utfärdande av ett båtförarcertifikat i samma grupp.
Artikel 4
Rådet skall senast den 31 december 1994, på grundval av ett förslag från kommissionen som skall inlämnas senast den 31 december 1993, med kvalificerad majoritet besluta om gemensamma bestämmelser för framförande på inre vattenvägar av fartyg som transporterar gods och passagerare.
1. Vid tillämpningen av artikel 4 skall kommissionen biträdas av en kommitté. Den skall bestå av företrädare för medlemsstaterna och ha en företrädare för kommissionen som ordförande.
Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Denna tolerans avser den normala kvantiteten svinn i samband med normal lagring eller bearbetning av jordbruksprodukter i intervention med beaktande av kraven på riktig förvaring av produkten.
Inga lagringsåtgärder har förekommit för griskött under lång tid och denna toleransnivå bör fastställas senare om lagringsåtgärder skulle vidtas på nytt.
Toleranserna har fastställts i sektorsvisa förordningar. De bör av hänsyn till rättslig förenkling fastställas i en enda förordning.
1. För varje jordbruksprodukt som är föremål för offentlig lagring fastställs en toleransnivå för kvantiteten svinn i samband lagringsåtgärder som vidtas i enlighet med godkända regler.
Artikel 2 1. Procentsatserna för normalt tillåtet svinn vid lagring fastställs härmed till följande:
KOMMISSIONENS FÖRORDNING (EEG) nr 1026/91 av den 22 april 1991 om ändring av förordning (EEG) nr 1208/81 om fastställande av en gemenskapsskala för klassificering av slaktkroppar av fullvuxna nötkreatur
med beaktande av rådets förordning (EEG) nr 1358/80 av den 5 juni 1980 om fastställande av orienterings- och interventionspriser för fullvuxna nötkreatur för 1980/1981 års regleringsår och om införande av en gemenskapsskala för klassificering av slaktkroppar av fullvuxna nötkreatur(1), särskilt artikel 4.1 i denna,
Med tanke på de genetiska förbättringar som är ett resultat av avel med nötkreatur bör gemenskapens skala för klassificering av slaktkroppar av vuxna nötkreatur anpassas så att hänsyn tas till förekomsten av djur med dubbelmuskulatur. Det bör därför finnas en möjlighet att frivilligt kunna införa en konformationsklass utöver de existerande klasserna.
1. Artikel 3 skall ersättas med följande:
A. Slaktkroppar av okastrerade ungdjur av hankön under två år.
D. Slaktkroppar av djur av honkön som har kalvat.
Kriterier för att skilja slaktkroppskategorier åt skall fastställas i enlighet med förfarandet i artikel 27 i förordning (EEG) nr 805/68.
b) fettgrupp
Medlemsstater som avser att använda denna möjlighet skall meddela kommissionen och övriga medlemsstater detta.
Artikel 2 Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
För att ta hänsyn till hävdvunnen praxis som fanns när förordning (EEG) nr 1576/89 trädde i kraft bör det vara tillåtet att behålla vissa sammansatta namn på likörer även om inte alkoholen erhållits eller uteslutande erhållits från den spritdryck som angivits. Det är nödvändigt att specificera villkor för beteckningen för sådana likörer för att undvika varje risk för förväxling med de spritdrycker som definieras i artikel 1.4 i förordning (EEG) nr 1576/89.
1. I enlighet med artikel 6.1 andra strecksatsen i förordning (EEG) nr 1576/89, skall användningen av kategoribeteckningar i sammansatta beteckningar vara förbjuden vid presentation av spritdrycker såvida inte alkoholen i drycken uteslutande härrör från den spritdryck som anges.
3. Vad beträffar märkning och presentation av likörer som anges i punkt 2 skall den sammansatta termen finnas på etiketten på en enda rad med samma typsnitt och färg, och ordet "likör" skall finnas i omedelbar närhet med bokstäver som inte är mindre än det typsnittet.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I artikel 8 i kommissionens förordning (EEG) nr 1538/91(2) fastställs tillämpningsföreskrifter för den valfria klassificeringen av fryst och djupfryst fjäderfäkött i viktklasser. Den omedelbara tillämpningen av dessa bestämmelser har visat sig utgöra ett hinder för importen från tredje land av fjäderfäkött som förpackats före nämnda förordnings ikraftträdande. Tillämpningen av artikel 8 bör därför uppskjutas till den 1 mars 1992.
Denna förordning träder i kraft den 20 juni 1991.
EUROPEISKA GEMENSKAPERNAS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Europaparlamentets yttrande(1), och
Behovet för dessa nya bestämmelser är så mycket större eftersom kontroll vid gränserna mellan medlemsstaterna skall slopas.
Man bör därför inom ramen för rådets beslut 90/424/EEG av den 26 juni 1990 om vissa utgifter på veterinärområdet(6) fastställa att gemenskapen skall bidra till finansieringen av genomförandet av de nya åtgärderna i fråga om datorisering av veterinärförfarandena vid import.
- Ett system för att förmedla relevant information när en officiell veterinär vid en gränskontrollstation beslutar att vidaresända en sändning.
2. Den datorisering som avses i punkt 1 skall uppfylla nuvarande internationell standard.
Artikel 3
Artikel 4
Artikel 5
Artikel 6
Beslut 88/192/EEG skall härmed upphöra att gälla.
1. Följande strecksats skall läggas till i artikel 4.1:
3. Följande mening skall läggas till i artikel 9.2 iii:
"- underrätta den officiella veterinären vid kontrollstället på bestämmelseorten om produkternas passage och om trolig ankomstdag via det datoriserade nätverket som länkar samman veterinärmyndigheter (Animo),".
6. I artikel 16.1 a skall första strecksatsen ersättas med följande:
8. Artikel 16.5 skall ersättas med följande:
Direktiv 91/496/EEG ändras på följande sätt:
3. I artikel 6.2 skall följande mening läggas till:
5. I artikel 12.1 c skall första strecksatsen ersättas med följande:
7. Artikel 12.4 skall ersättas med följande:
Artikel 10
Följande artikel skall läggas till i beslut 90/424/EEG:
Artikel 12
1. Kommissionen skall bistås av Ständiga veterinärkommittén som bildats genom beslut 68/361/EEG(8), hädanefter kallad 'kommittén`.
4. a) Kommissionen skall själv anta förslaget och tillämpa det omedelbart om det inte strider mot kommitténs yttrande.
Artikel 14
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
I syfte att säkerställa att systemet Animo fungerar smidigt bör åtgärder vidtas för en harmonisering av samarbetsformerna mellan Animo datacentrum och medlemsländerna.
Artikel 1
Artikel 2
- innehåller en klausul om årlig översyn,
- anger följande taxa:
Artikel 3
Den sammanlagda årliga kostnaden för att delta i systemet som avses i artikel 2a femte strecksatsen och som inte skall överstiga det belopp som är fastställt för det första året, och dess fördelning mellan medlemsstaterna skall tas upp till förnyad prövning före den 1 juli 1993. Det maximala priset för varje medlemsstat under såväl det andra som tredje året skall dock inte öka med mer än 10 % av priset för det första året.
Artikel 6
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
Med hänsyn till de specifikationer som antagits genom Codex Alimentarius och till ny produktionsteknik är det nödvändigt att ändra rådets direktiv 78/663/EEG(2), senast ändrat genom kommissionens direktiv 90/612/EEG(3).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 3
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
i samarbete med Europaparlamentet(2),
Åtgärderna för en tillnärmning av de bestämmelser i medlemsstaterna som hänför sig till den inre marknadens upprättande och funktion skall, vad beträffar hälsan, säkerheten och skyddet för människan och miljön, utgå från en hög skyddsnivå.
Bestämmelser bör fastställas för att införa ett anmälningsförfarande, varigenom en anmälan som gjorts i en medlemsstat gäller i hela gemenskapen. För ämnen som tillverkas utanför gemenskapen kan det vara lämpligt att tillverkaren utser en representant i gemenskapen som ensam svarar för anmälan.
Kommissionen har i enlighet med artikel 13.1 i direktiv 67/548/EEG(6) och enligt riktlinjer fastställda i kommissionens beslut 81/437/EEG gjort upp en förteckning över ämnen som fanns på marknaden i gemenskapen den 18 september 1981 (EINECS), vilken har publicerats i Europeiska gemenskapernas officiella tidning(7).
För att stärka miljöskyddet och arbetarskyddet bör säkerhetsdatablad om farliga ämnen finnas tillgängliga för yrkesmässiga användare.
Enligt artikel 2 i direktiv 67/548/EEG klassificeras ämnen och preparat enligt allmänna definitioner som giftiga, hälsoskadliga, frätande eller irriterande. Erfarenheterna har visat att det är nödvändigt att förbättra denna klassificering. Exakta kriterier för klassificeringen bör anges. Enligt artikel 3 i direktivet skall också en bedömning göras av ämnets miljöfarlighet, vilket gör det nödvändigt att ange vissa kriterier och parametrar för bedömningen och införa ett undersökningsprogram i flera steg.
Medlemsstaterna bör i vissa fall tillåtas att vidta egna skyddsåtgärder.
Artikel 1
b) utbyte av information om anmälda ämnen,
a) Sådana farmaceutiska produkter för användning inom human- eller veterinärmedicin som avses i direktiv 65/65/EEG(1), senast ändrat genom direktiv 87/21/EEG(2).
d) Livsmedel.
g) Radioaktiva ämnen som avses i direktiv 80/836/EEG(7).
Detta direktiv skall inte heller gälla
Definitioner
b) preparat: blandningar eller lösningar som består av två eller flera ämnen.
- för ämnen framställda inom gemenskapen: av den tillverkare som släpper ut ett ämne på marknaden, ensamt eller i ett preparat,
g) processinriktad forskning och utveckling: vidareutvecklandet av ett ämne, varvid användningsområden för ämnet testas genom pilotförsök eller provtillverkning.
a) explosiva ämnen och preparat: fasta och flytande ämnen och ämnen i pasta- eller geléform som även utan närvaro av atmosfäriskt syre kan ge upphov till en exoterm reaktion och därvid snabbt avge gaser, och som under angivna testförhållanden detonerar, snabbt deflagrerar eller delvis inneslutna exploderar vid uppvärmning,
d) Mycket brandfarliga ämnen och preparat:
- flytande ämnen och preparat med mycket låg flampunkt, eller
f) Mycket giftiga ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden i mycket små mängder leder till döden eller ger akuta eller kroniska skador.
i) Frätande ämnen och preparat: ämnen och preparat som vid kontakt med levande vävnader kan förstöra dessa.
l) Cancerogena ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan orsaka eller öka förekomsten av cancer.
o) Miljöfarliga ämnen och preparat: ämnen och preparat som om de kommer ut i miljön utgör eller kan utgöra en omedelbar eller fördröjd fara för en eller flera delar av miljön.
1. Tester på kemikalier som utförs inom ramen för detta direktiv skall som allmän princip utföras enligt de metoder som föreskrivs i bilaga 5. Ämnenas fysikaliskkemiska egenskaper skall bestämmas enligt de metoder som anges i bilaga 5 A. Deras toxicitet skall bestämmas enligt metoderna i bilaga 5 B och deras miljöfarlighet enligt metoderna i bilaga 5 C.
2. De verkliga och potentiella riskerna för människan och miljön skall bedömas enligt de principer som antagits den 30 april 1993 i enlighet med förfarandet i artikel 29.4 b. Dessa principer skall regelbundet ses över och vid behov ändras enligt samma förfarande.
1. Ämnen skall klassificeras på grundval av sina inneboende egenskaper enligt de i artikel 2.2 fastställda kategorierna. Vid klassificering av ämnen skall hänsyn också tas till föroreningar, om dessa förekommer i koncentrationer som överstiger de koncentrationsgränser som anges i punkt 4 i denna artikel och i artikel 3 i direktiv 88/379/EEG.
Artikel 5
- anmälts till den behöriga myndigheten i en av medlemsstaterna enligt detta direktiv,
2. Bestämmelserna i andra strecksatsen i punkt 1 skall gälla tills ämnet upptas i bilaga 1 eller tills ett beslut att inte ta upp ämnet har fattats enligt förfarandet i artikel 29.
Tillverkare, distributörer och importörer av i EINECS upptagna farliga ämnen som ännu inte finns med i bilaga 1 skall vara skyldiga att utföra en undersökning för att utröna vilka relevanta och tillgängliga data som finns om ämnenas egenskaper. Ämnena skall förpackas och provisoriskt märkas på grundval av denna information i enlighet med bestämmelserna i artikel 22-25 och enligt kriterierna i bilaga 6.
1. Om inte annat följer av artikel 1.2, 8.1, 13 och 16.1 skall en anmälare av ett ämne lämna en anmälan till den behöriga myndighet som avses i artikel 16.1 i den medlemsstat där ämnet framställs eller, om tillverkaren befinner sig utanför gemenskapen, i den medlemsstat där anmälaren är verksam. Anmälan skall ha följande innehåll:
- Föreslagen klassificering och märkning av ämnet enligt detta direktiv.
- Anmälaren kan, om han så önskar, bifoga en motiverad begäran om att bestämmelserna i artikel 15.2 inte skall tillämpas i fråga om anmälan under en tidsperiod som inte i något fall får överstiga ett år från tidpunkten för anmälan.
- när den mängd av ämnet som släppts ut på marknaden uppnår 10 ton per år och tillverkare, eller när den totala mängd av ämnet som släppts ut på marknaden uppnår 50 ton per tillverkare, varvid den behöriga myndigheten kan kräva att en del eller samtliga kompletterande tester/undersökningar som föreskrivs i bilaga 8 nivå 1 skall utföras inom den tid som den behöriga myndigheten bestämmer,
3. När kompletterande tester utförs, i enlighet med kraven i punkt 2 eller frivilligt, skall anmälaren meddela resultaten till den behöriga myndigheten.
1. Om inte annat följer av artikel 1.2, 13.1 och 16.1 skall en anmälare som avser att släppa ut ett ämne på marknaden inom gemenskapen i mängder som understiger ett ton per år och tillverkare vara skyldig att till den behöriga myndighet som avses i artikel 16.1 i den medlemsstat där ämnet framställs eller, om tillverkaren befinner sig utanför gemenskapen, i den medlemsstat där anmälaren är verksam, lämna en anmälan med följande innehåll:
2. Om mängden som släpps ut på marknaden understiger 100 kg per år och tillverkare kan anmälaren, om inte annat följer av artikel 16.1, begränsa uppgifterna i den ovannämnda dokumentationen till vad som föreskrivs i bilaga 7 C.
5. De ämnen som anmälts enligt punkt 1 och 2 skall, i den mån anmälaren rimligen kan förväntas känna till deras farliga egenskaper, förpackas och provisoriskt märkas i enlighet med reglerna i artikel 22-25 och enligt kriterierna i bilaga 6. Om det ännu inte är möjligt att märka dem i enlighet med principerna i artikel 23, skall utöver märkningen från de redan utförda testerna på etiketten anges "Varning - ämnet ännu inte fullständigt testat".
Om uppgifter enligt artikel 7 och 8 lämnats minst 10 år tidigare behöver en anmälare inte tillhandahålla sådana uppgifter som krävs för dokumentationen enligt bilaga 7 A 7 D, förutom uppgifterna under punkt 1 och 2 i de nämnda bilagorna.
1. Om inte annat anges av den behöriga myndigheten, får ämnen som anmälts enligt artikel 7.1 släppas ut på marknaden tidigast 60 dagar efter det att myndigheten mottagit en dokumentation som överensstämmer med kraven i detta direktiv.
Om den behöriga myndigheten anser att dokumentationen inte uppfyller kraven i direktivet och meddelar anmälaren detta enligt artikel 16.3, får ämnet släppas ut på marknaden tidigast 30 dagar efter det att myndigheten mottagit de uppgifter som behövs för att anmälan skall överensstämma med direktivets krav. Om anmälaren underrättats enligt artikel 16.3 att dokumentationen har godtagits, gäller dock att ämnet får släppas ut på marknaden tidigast 15 dagar efter det att den behöriga myndigheten mottagit dokumentationen.
Om det i fråga om ämnen som framställs utanför gemenskapen finns mer än en anmälan för ett ämne framställt av samma tillverkare, skall kommissionen och de nationella myndigheterna fastställa den totala årliga mängden som släpps ut på marknaden inom gemenskapen på grundval av de uppgifter som lämnats enligt artikel 7.1, 8.1 och 14. Skyldigheten att utföra kompletterande tester enligt artikel 7.2 åligger samtliga anmälare gemensamt.
I fråga om polymerer skall särskilda bestämmelser fastställas i bilaga 7 i den form som anges i bilaga 7 D och enligt det förfarande som anges i artikel 29.4 b angående den dokumentation som enligt artikel 7.1 och 8.1 skall ingå i anmälan.
1. Bestämmelserna i artikel 7, 8, 14 och 15 tillämpas inte på följande ämnen:
- Ämnen som endast används i livsmedel och omfattas av direktiv 89/107/EEG(2), samt ämnen som endast används som smakämnen i livsmedel och omfattas av direktiv 88/388/EEG.
2. De ämnen som anges nedan skall anses ha anmälts enligt detta direktiv om följande villkor är uppfyllda:
- Ämnen som släpps ut på marknaden i begränsade mängder, inte i något fall över 100 kg per tillverkare och år, och som är avsedda enbart för vetenskaplig forskning och utveckling som utförs under kontrollerade förhållanden.
I undantagsfall får den ovannämnda ettårsperioden förlängas med ytterligare ett år, om anmälaren på ett tillfredsställande sätt kan visa för den behöriga myndigheten att en sådan förlängning är motiverad.
Artikel 14
- förändringar i de årliga eller totala mängder som släpps ut på den gemensamma marknaden av honom eller, om ämnet tillverkas utanför gemenskapen och anmälaren ensam företräder denne, av honom eller någon annan,
- alla ändringar i ämnenas sammansättning som avses i bilaga 7 A, B eller C, avsnitt 1.3,
Artikel 15
2. Innan försök utförs på ryggradsdjur i syfte att upprätta en anmälan i enlighet med artikel 7.1 eller 8.1, och om inte annat följer av punkt 1, skall den som avser att anmäla ett ämne fråga den behöriga myndigheten i den medlemsstat där han ämnar inlämna sin anmälan
a) Den behöriga myndighet som mottar förfrågan finner det styrkt att den nya anmälaren ämnar släppa ut ämnet på marknaden i de uppgivna mängderna.
Den första anmälaren och den nya anmälaren skall vidta alla rimliga åtgärder för att nå en överenskommelse om utbyte av information, så att upprepade tester på ryggradsdjur kan undvikas.
Artikel 16
Om det visar sig nödvändigt för bedömningen av riskerna med ett ämne får de behöriga myndigheterna dessutom begära ytterligare underlag eller kompletterande tester angående ämnen eller nedbrytningsprodukter som har anmälts eller beträffande vilka uppgifter lämnats enligt detta direktiv. Därvid kan begäras att sådana uppgifter som avses i bilaga 8 skall lämnas tidigare än som anges i artikel 7.2.
- begära att anmälaren tillhandahåller ämnet i sådana mängder som anses nödvändiga för att utöva kontrolltester,
2. I fråga om anmälningar som lämnats i enlighet med artikel 7 skall myndigheterna inom 60 dagar efter mottagandet skriftligen underrätta anmälaren om huruvida anmälan anses överensstämma med detta direktiv.
4. Beträffande ämnen som framställts utanför gemenskapen och för vilka fler än en anmälan inkommit som avser ett ämne som framställs av en och samma tillverkare, skall de behöriga myndigheterna tillsammans med kommissionen svara för beräkningen av de årliga och totala mängder som släpps ut på marknaden inom gemenskapen. Om de mängder uppnås som anges i artikel 7.2, skall den behöriga myndighet som mottagit anmälan eller anmälningarna kontakta anmälarna, meddela dem vilka de andra anmälarna är och upplysa dem om deras gemensamma ansvar enligt artikel 11.
Artikel 17
I fråga om de kompletterande uppgifter som avses i artikel 16.1 skall den behöriga myndigheten meddela kommissionen vilka tester som valts, skälen för detta, testresultaten och, i tillämpliga fall, bedömningen av resultaten. I fråga om uppgifter som mottagits i enlighet med artikel 13.2 skall den behöriga myndigheten till kommissionen vidarebefordra sådana som kan vara av allmänt intresse för kommissionen och andra behöriga myndigheter.
Kommissionens skyldigheter
Artikel 19
I fråga om anmälningar och uppgifter som lämnats i enlighet med artikel 7.1, 7.2 och 7.3, samt skall industriell och kommersiell sekretess inte gälla för
c) fysikalisk-kemiska uppgifter om ämnet enligt avsnitt 3 i bilaga 7 A 7 C,
h) informationen som lämnas i säkerhetsdatabladet,
2. Den myndighet som mottagit anmälan eller uppgifterna skall på eget ansvar avgöra vilka uppgifter som omfattas av industriell och kommersiell sekretess i enlighet med punkt 1.
Farliga ämnen kan på begäran från den behöriga myndighet som mottog anmälan upptas endast under sina handelsnamn tills de upptas i bilaga 1.
- får lämnas ut endast till de myndigheter vilkas ansvars områden anges i artikel 16.1,
Utväxling av den sammanfattade dokumentationen
2. Kommissionen skall utforma ett gemensamt system för utväxling av de uppgifter som avses i artikel 17 och 18.1. Detta system skall antas enligt förfarandet i artikel 29.
1. Kommissionen skall upprätta en förteckning över samtliga ämnen som anmälts enligt detta direktiv. Listan skall sammanställas i enlighet med bestämmelserna i kommissionens beslut 85/71/EEG(1).
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att tillse att farliga ämnen endast kan släppas ut på marknaden om förpackningen uppfyller följande krav:
c) Förpackningen och förslutningarna skall genomgående vara starka och stadiga så att de inte kan lossna och så att de tål normal påfrestning under hanteringen.
f) Behållare som innehåller ämnen som säljs till eller tillhandahålls allmänheten och är märkta "hälsoskadligt", "synnerligen brandfarligt" eller "mycket brandfarligt" enligt detta direktiv skall, oberoende av storleken, vara försedda med en varningsmärkning som kan uppfattas vid beröring.
4. Ändringar i de tekniska specifikationerna för de anordningar som avses i punkt 1 e och 1 f skall beslutas enligt förfarandet i artikel 29.4 och återfinns i punkt A och B i bilaga 9 till detta direktiv.
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att säkerställa att farliga ämnen endast släpps ut på marknaden om märkningen på förpackningen uppfyller följande krav.
b) Namn och fullständig adress med telefonnummer för den i gemenskapen verksamma person som är ansvarig för att ämnet släpps ut på marknaden, antingen denne är tillverkare, importör eller distributör.
- Om symbolen T är obligatorisk behöver inte symbolerna X och C anges, om inte annat följer av bilaga 1.
d) Standardfraser (R-fraser) som anger särskilda risker som är förenade med användningen av ämnet. R-fraserna skall överensstämma med vad som anges i bilaga 3. De R-fraser som skall användas för varje ämne anges i bilaga 1. För farliga ämnen som ännu inte finns upptagna i bilaga 1 skall R-fraser tilldelas enligt reglerna i bilaga 6.
För ämnen som finns upptagna i bilaga 1 skall dessutom ordet "EEG-märkning" anges på etiketten.
Artikel 24
2. Etikett krävs inte om uppgifterna är tydligt angivna på själva förpackningen i enlighet med punkt 1.
Särskilda bestämmelser om de upplysningarna som avser utformning och dimensioner förs in i bilaga 6 enligt förfarandet i artikel 29.4 b.
a) När en yttre förpackning innehåller en eller flera inre förpackningar, om den yttre förpackningen är märkt enligt internationella regler för transport av farliga ämnen och den inre förpackningen eller de inre förpackningarna är märkta i enlighet med detta direktiv.
- när det behövs för särskilda typer av förpackningar såsom transportabla gasflaskor, förpackningen är märkt i enlighet med de särskilda krav som anges i bilaga 6.
Undantag från kraven på märkning och förpackning
2. Dessutom får medlemsstaterna
c) om förpackningen är för liten för märkning enligt artikel 23 och 24 och det inte finns någon anledning att anta att de som hanterar ämnet eller andra kan utsättas för fara, trots bestämmelserna i ovanstående artiklar tillåta att förpackningar med explosiva, mycket giftiga eller giftiga ämnen märks på annat lämpligt sätt.
Artikel 26
Artikel 27
Informationen kan lämnas på papper eller elektroniskt. Därefter skall tillverkaren, importören eller distributören till mottagaren av säkerhetsdatabladet sända sådan ny relevant information om ämnet som kommer till hans kännedom.
Anpassning till den tekniska utvecklingen
Förfarandet vid anpassning till den tekniska utvecklingen
3. Kommissionen skall själv anta förslaget om det är förenligt med kommitténs yttrande.
b) I fråga om åtgärder för anpassning till den tekniska utvecklingen som avser bilaga 2, 6, 7 och 8 skall kommissionen om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits själv besluta att de föreslagna åtgärderna skall vidtas, såvida inte rådet med enkel majoritet har avvisat förslaget.
Medlemsstaterna får inte på grunder som rör anmälan, klassificering, förpackning eller märkning i detta direktivs mening förbjuda, begränsa eller hindra att ämnen som uppfyller kraven i detta direktiv släpps ut på marknaden.
1. Om en medlemsstat i ljuset av ny information på goda grunder anser att ett ämne som har bedömts uppfylla kraven i detta direktiv ändå utgör en fara för människan eller miljön på grund av att klassificeringen, förpackningen eller märkningen inte längre är riktig, kan den tillfälligt omklassificera ämnet eller, om så är nödvändigt, förbjuda att ämnet släpps ut på marknaden eller föreskriva att särskilda villkor skall gälla inom det egna territoriet. Den skall omedelbart meddela kommissionen och de andra medlemsstaterna om varje sådan åtgärd och motivera sitt beslut.
Artikel 32
2. Vart tredje år skall kommissionen på grundval av de uppgifter som avses i punkt 1 upprätta en samlad rapport som skall överlämnas till medlemsstaterna."
- Bilaga 2 ändras genom tillägget av en symbol som betecknar miljöfara enligt bilaga 1 i detta direktiv.
- Bilaga 8 ersätts av bilaga 4 till detta direktiv.
- I artikel 6.2 g ersätts "artikel 6" med "artikel 23".
- I det andra och det åttonde stycket i ingressen ersätts hänvisningen till direktiv 79/831/EEG med en hänvisning till föreliggande direktiv.
- Artikel 3.5 o skall ha följande lydelse:
- den koncentration som anges i punkt 6 i bilaga 1 (tabell VI) till detta direktiv, om ämnet inte är upptaget i bilaga 1 till direktiv 67/548/EEG eller förekommer där, men utan angivande av koncentrationsgränser."
- antingen de koncentrationer som anges i bilaga 1 till direktiv 67/548/EEG för ämnet i fråga, eller
"q) Preparat skall anses behöva behandlas som skadliga för fortplantningen och tilldelas minst farosymbolen och faroangivelsen "giftigt" om de innehåller ett ämne som har sådana verkningar och som tilldelas minst en av de R-fraser enligt bilaga 6 till direktiv 67/548/EEG som betecknar ämnen som är skadliga för fortplantningen i kategori 3, i koncentrationer som motsvarar eller överstiger
- I artikel 6.1 a ersätts "artikel 15.1" med "artikel 22.1".
- I artikel 7.1 ersätts "artikel 16.2 c" av "artikel 23.2 c".
Särskilda bestämmelser om upplysningarnas uppställning och format förs in i bilaga 6 till direktiv 67/548/EEG i enlighet med förfarandet i artikel 28.4 b i nämnda direktiv".
- I bilaga 1 tabell 6 ersätts "teratogena ämnen" med "ämnen som är skadliga för fortplantningen".
2. När dessa åtgärder beslutas av medlemsstaterna skall författningarna innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av ekonomiska och sociala kommitténs yttrande(), och
Under övergångstiden bör vissa undantag från reglerna beträffande skatternas antal och nivå vara möjliga.
Direktiv 77/388/EEG ändras på följande sätt:
På grundval av den rapport om hur övergångsbestämmelserna har fungerat och de förslag till slutgiltiga bestämmelser som kommissionen skall lägga fram i överensstämmelse med artikel 281, skall rådet före den 31 december 1995 enhälligt besluta om den lägsta skattesatsnivå som efter den 31 december 1996 skall tillämpas såsom normalskattesats.
c) Regler om vilka skattesatser som skall tillämpas på konstverk, antikviteter och samlarföremål fastställs genom direktivet med specialbestämmelser för begagnade varor, konstverk, antikviteter och samlarföremål. Rådet skall anta detta direktiv före den 31 december 1992.
e) De regler och skattesatser som skall tillämpas på guld skall fastställas genom ett direktiv med specialbestämmelser om guld. Kommissionen skall lägga fram ett förslag härom i sådan tid att det kan enhälligt antagas av rådet före den 31 december 1992.
3. Följande stycke läggs till i artikel 12.4:
"2. Utan hinder av artikel 12.3 skall följande bestämmelser gälla under den övergångsperiod som nämns i artikel 28l:
I händelse av att bestämmelserna i denna punkt för Irlands del skulle skapa snedvridning av konkurrensen när det gäller tillhandahållande av energiprodukter för uppvärmning och belysning, kan kommissionen på särskild begäran ge Irland rätt att tillämpa en reducerade skattesats på sådant tillhandahållande, i enlighet med artikel 12.3. I sådant fall skall Irland inlämna sin begäran till kommissionen tillsammans med alla nödvändiga upplysningar. Om kommissionen inte har fattat något beslut inom tre månader efter mottagandet av denna begäran, skall Irland anses ha fått rätt att tillämpa den föreslagna reducerade skattesatsen.
d) Medlemsstater som den 1 januari 1991 tillämpade en reducerad skattesats på restaurangtjänster, barnkläder, barnskor och bostäder får fortsätta att tillämpa denna på dessa områden.
g) Rådet skall på grundval av en rapport från kommissionen före den 31 december 1994 på nytt granska bestämmelserna i a-f ovan med särskild hänsyn till den inre marknadens riktiga funktion. I den händelse betydande snedvridning av konkurrensen uppstår, skall rådet på kommissionens förslag enhälligt besluta om lämpliga åtgärder."
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 december 1992. De skall genast underrätta kommissionen härom.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
I kommissionens förordning (EEG) nr 410/90(3) fastställs kvalitetsnormer för kiwifrukt.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för frukt och grönsaker.
"Den skall ha sorttypiska egenskaper. Följande smärre fel är dock tillåtna om de inte påverkar produktens allmänna utseende, kvaliteten, hållbarheten och förpackningens presentation:
- Ytliga skador på skalet som täcker en yta av högst 1 cm².
" - Flera mer uttalade "Hayward-märken" med mindre förhöjning."
3. Följande ändringar skall göras i del V. "Bestämmelser angående presentation":
KOMMISSIONENS FÖRORDNING (EEG) nr 762/92 av den 27 mars 1992 om ändring av bilaga V i rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), ändrad genom kommissionens förordning (EEG) nr 675/92(2), särskilt artikel 11, och med beaktande av följande:
Bestämmelserna i denna förordning är förenliga med yttrandet från Kommittén för anpassning till den tekniska utvecklingen av direktiven om avlägsnande av tekniska handelshinder inom den veterinärmedicinska sektorn, inrättad genom artikel 2b i rådets direktiv 81/852/EEG(5), ändrat genom direktiv 87/20/EEG(6).
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Inom den allmänna ramen för den förnyade medelhavspolitiken antog rådet och kommissionen en resolution om handel med icke-medlemsstater i medelhavsområdet på rådets möte den 18 och 19 december 1990, i syfte att stärka banden och öka samarbetet med länderna i regionen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Punkt 1 tillämpas inom ramarna, om sådana finns, för tullkvoter och tidsscheman som fastställts i de protokoll som avses i den punkten och skall beakta de särskilda bestämmelser som där fastställs.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(2),
Branschorganisationer som bildats av enskilda eller grupper och som representerar en betydande del av de olika kategorier som är sysselsatta med produktion, beredning och avsättning inom tobakssektorn skulle sannolikt komma att bidra till att större hänsyn tas till situationen på marknaden liksom till att uppmuntra förändringar i det ekonomiska beteendet i syfte att förbättra kunskapen om och organisationen av produktionen, beredningen och avsättningen. Deras verksamhet skulle i vissa fall kunna bidra till att förbättra balansen på marknaden och därigenom medverka till att målen enligt artikel 39 i fördraget uppfylls. Det bör därför fastställas vilka åtgärder som skulle kunna utgöra ett sådant bidrag från branschorganisationernas sida.
Andra verksamheter som de erkända branschorganisationerna bedriver kan vara av allmänt ekonomiskt eller tekniskt intresse för tobakssektorn och därmed vara värdefulla för alla som är sysselsatta inom branscherna i fråga, vare sig de är medlemmar i organisationen eller inte. I dessa fall förefaller det rimligt att icke medlemmar betalar den medlemsavgift som är avsedd att täcka andra kostnader än de rent administrativa som uppkommer som en direkt följd av verksamheten i fråga.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
b) Utarbetande av standardavtal som är i överensstämmelse med gemenskapens bestämmelser.
e) Omorientering av branschen mot produkter som bättre tillgodoser marknadens behov och hänsynen till folkhälsan.
2. Före erkännandet skall medlemsstaterna anmäla till kommissionen vilka branschorganisationer som ansökt om erkännande och lämna all nödvändig information om vilka näringsgrenar de omfattar, hur representativa de är, vilka verksamheter de bedriver samt den övriga information som behövs för att ta ställning till ansökan.
a) de krav som anges i denna förordning inte längre uppfylls,
Medlemsstaterna skall omedelbart underrätta kommissionen om beslut om återkallande av erkännandet.
a) helt eller delvis bedriver sin verksamhet inom flera medlemsstaters territorier eller inom hela gemenskapen,
2. Kommissionen skall underrätta de medlemsstater inom vilkas territorier branschorganisationen bildats och dess verksamhet bedrivs om inkomna ansökningar om erkännande. De berörda medlemsstaterna skall därefter ha två månader på sig att inkomma med synpunkter.
Artikel 5
Erkännandet av branschorganisationer innebär att de tillåts bedriva de verksamheter som anges i artikel 2.3 på de villkor som föreskrivs i denna förordning.
2. Punkt 1 skall tillämpas endast om
Avtalen och de samordnade förfarandena får inte träda i kraft förrän denna period löpt ut.
- kan medföra att den gemensamma organisationen av marknaden störs,
- kan innebära särbehandling eller sätta konkurrensen ur spel för en betydande del av produkterna i fråga.
1. Branschorganisationerna kan begära att vissa av deras avtal eller samordnade förfaranden inom det område där de är verksamma för en begränsad tid görs bindande för enskilda och grupper inom den berörda ekonomiska sektorn som inte är medlemmar i någon organisation som ingår i branschorganisationen.
a) Kunskap om produktionen och marknaden.
d) Fastställande av minimistandarder för förpackning och presentation.
Artikel 9
2. Vid slutet av denna period och innan beslut fattas, skall medlemsstaterna anmäla till kommissionen vilka bestämmelser de avser att göra bindande och samtidigt lämna all relevant information. I anmälan skall ingå alla de synpunkter som erhållits efter offentliggörandet enligt punkt 1 och en bedömning av ansökan om utvidgad tillämpning.
Om förutsättningarna för att avge ett detaljerat utlåtande enligt artikel 9 i det direktivet är uppfyllda, skall kommissionen, vägra godkänna de bestämmelser för vilka utvidgad tillämpning begärs, utan att detta påverkar tillämpningen av punkt 5.
- förhindrar konkurrensen på en betydande del av den gemensamma marknaden,
6. De bestämmelser för vilka man ansökt om utvidgad tillämpning skall offentliggöras i Europeiska gemenskapernas officiella tidning.
1. När en eller flera av de i punkt 2 angivna verksamheterna bedrivs av en erkänd branschorganisation och är av allmänt ekonomiskt intresse för de personer vilkas verksamhet är knuten till en eller flera av produkterna, får medlemsstaten som beviljat erkännandet eller kommissionen, om erkännandet beviljats i enlighet med artikel 4, besluta att enskilda eller grupper som inte är medlemmar i sammanslutningen men som drar nytta av dess verksamhet skall betala till organisationen hela eller del av medlemsavgiften, i den mån medlemsavgiften är avsedd att täcka kostnader som är en direkt följd av verksamheten med undantag av varje form av administrationskostnad.
- Undersökningar om hur kvaliteten på bladtobak och tobak i balar kan förbättras.
4. Om de verksamheter som en av kommissionen enligt artikel 4 erkänd branschorganisation bedriver är av allmänt ekonomiskt intresse, skall kommissionen anmäla sitt förslag till beslut till de berörda medlemsstaterna, som sedan har två månader på sig att lämna sina synpunkter.
Artikel 12
RÅDETS FÖRORDNING (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel
Med tanke på mångfalden av marknadsförda produkter och överflödet av information om dem måste konsumenterna för att kunna göra ett bra val få klar och koncis information om produkternas ursprung.
Det finns emellertid nationella olikheter i sättet att ordna registrering av ursprungsbeteckning och geografisk beteckning. En gemenskapsmetod bör planeras. Ett gemensamt regelverk för skydd av dessa beteckningar gör det möjligt att utveckla dessa, eftersom ett sådant skydd med enhetlig metod säkerställer konkurrens på lika villkor mellan produkter med sådana beteckningar och höjer produkternas trovärdighet i konsumenternas ögon.
Nuvarande bruk gör det lämpligt att definiera två slags geografiska beskrivningar, nämligen skyddade geografiska beteckningar och skyddade ursprungsbeteckningar.
Registreringsförfarandet bör ge var och en som personligen och direkt berörs i en medlemsstat möjlighet att tillvarata sina rättigheter genom att till kommissionen framställa invändningar.
Föreskrifter bör införas för ett förfarande som innebär nära samverkan mellan medlemsstaterna och kommissionen genom en regleringskommitté som inrättas för ändamålet.
1. Denna förordning fastställer regler för skydd av ursprungsbeteckningar och geografiska beteckningar för sådana jordbruksprodukter som är avsedda att förtäras av människor och som avses i bilaga 2 till fördraget och för sådana livsmedel som avses i bilaga 1 till denna förordning och de jordbruksprodukter som förtecknats i bilaga 2 till denna förordning.
2. Denna förordning skall tillämpas utan att påverka andra särskilda gemenskapsregler.
och - vars kvalitet eller egenskaper helt eller väsentligen beror på viss geografisk omgivning med de naturliga och mänskliga faktorer som därtill hör och vars framställning, bearbetning och beredning äger rum i det ifrågavarande geografiska området.
och - som besitter viss kvalitet, har visst anseende eller äger viss annan egenskap som kan hänföras till detta geografiska ursprung och som framställs, bearbetas och bereds i det ifrågavarande geografiska området.
- det område där råvarorna framställs är begränsat,
5. Vid tolkningen av punkt 4 får endast levande djur, kött och mjölk betraktas som råvaror. Bruk av andra råvaror kan godkännas i enlighet med det förfarande som stadgas i artikel 15.
Artikel 3
När det skall avgöras huruvida ett namn har blivit generiskt, skall hänsyn tas till alla faktorer, i synnerhet
- berörd nationell lagstiftning och gemenskapslagstiftning.
3. Innan denna förordning träder i kraft skall rådet efter beslut med kvalificerad majoritet och på förslag av kommissionen upprätta och i Europeiska gemenskapernas officiella tidning offentliggöra en icke uttömmande vägledande förteckning över namn på jordbruksprodukter och livsmedel som omfattas av denna förordning och enligt punkt 1 skall betraktas som generiska och sålunda såsom icke registrerbara enligt denna förordning.
2. Produktspecifikationen skall omfatta bl. a. följande uppgifter:
c) En definition av det geografiska området och i förekommande fall uppgifter som visar att kraven i artikel 2.4 är uppfyllda.
f) Uppgifter som påvisar sambandet med den lokala omgivningen eller det geografiska ursprunget i den mening som avses i artikel 2.2 a respektive b.
i) De övriga uppgifter som föreskrivits av gemenskapen och/eller nationella stadganden.
3. Ansökan om registrering skall innehålla den produktspecifikation som avses i artikel 4.
Om ansökningen avser ett namn på ett geografiskt område som sträcker sig in i en annan medlemsstat, skall denna senare medlemsstat tillfrågas innan beslut fattas.
2. Om kommissionen med beaktande av vad som har framkommit vid den granskning som avses i punkt 1 finner att namnet är skyddsberättigat, skall den i Europeiska gemenskapernas officiella tidning offentliggöra sökandens namn och adress, produktens benämning, ansökningens huvudsakliga innehåll, hänvisningar till de nationella föreskrifter som kan finnas om produktens framställning och beredning och när så behövs motiveringen för sina slutsatser.
- de namn som införts i registret,
Innan offentliggörande enligt punkt 2 och 4 och registrering enligt punkt 3 sker, får kommissionen inhämta yttrande av den kommitté som föreskrivs i artikel 15.
2. Medlemsstaternas behöriga myndigheter skall se till, att alla personer som kan visa att de har ett lagligen berört ekonomiskt intresse tillåts ta del av ansökningen. Därutöver kan varje medlemsstat i enlighet med vad som eljest gäller i medlemsstaten i fråga bereda även andra parter med ett lagligen berört intresse åtkomst till ansökningen.
- Invändningen visar att överträdelse skett av de villkor som avses i artikel 2.
5. När en invändning enligt punkt 4 är sådan att den skall tas upp till behandling, skall kommissionen uppmana de berörda medlemsstaterna att inom tre månader söka förlikning i enlighet med sina egna förfaranden. Därefter skall förfaras på endera av följande sätt.
Artikel 8
Medlemsstaten i fråga får begära att produktspecifikationen ändras, t. ex. för att ta hänsyn till ny teknik och nya forskningsrön eller för att omdefiniera ett geografiskt område.
Artikel 10
3. Utsedda kontrollmyndigheter och godkända privata organ måste kunna garantera objektivitet och opartiskhet gentemot alla producenter och produktförädlare som underställs deras kontroll och ha ständig tillgång till den kvalificerade personal och de övriga resurser som behövs för att genomföra kontroller av jordbruksprodukter och livsmedel som bär en skyddad beteckning.
4. Om en utsedd kontrollmyndighet respektive ett godkänt privat organ i en medlemsstat konstaterar att en jordbruksprodukt eller ett livsmedel som bär en skyddad ursprungsbeteckning där inte produktspecifikationens kriterier uppfylls, skall kontrollorganet vidta de åtgärder som är nödvändiga för att se till, att denna förordning följs. Kontrollorganet skall underrätta medlemsstaten om de åtgärder som vidtagits i samband med kontrollerna. Berörda parter måste underrättas om alla beslut som fattas.
7. Kostnaderna för de kontroller som föreskrivs i denna förordning skall bäras av de producenter som använder den skyddade beteckningen.
2. Den medlemsstat som avses i punkt 1 skall rikta anmärkningen till den medlemsstat som är berörd. Denna skall granska anmärkningen och underrätta den klagande medlemsstaten om vad som framkommit och i förekommande fall om de åtgärder som har vidtagits.
Artikel 12
2. Om tredje lands skyddade beteckning sammanfaller med en skyddad beteckning i gemenskapen, skall registrering ske med vederbörlig hänsyn till lokalt och traditionellt språkbruk och till risken för förväxling i praktiken.
1. Registrerade beteckningar skall skyddas mot följande.
c) Varje annan osann eller vilseledande uppgift om ursprung, härkomst, beskaffenhet eller väsentliga egenskaper hos produkten på dennas inre eller yttre förpackning, reklammaterial eller handlingar, liksom förpackning av produkten i behållare som är ägnad att inge en oriktig föreställning om produktens verkliga ursprung.
2. Medlemsstaterna får dock låta nationella regler om rätt att bruka sådana beteckningar som avses i punkt 1 b bestå under högst fem år efter den dag denna förordning offentliggörs under förutsättning
Detta undantag får dock inte leda till att produkterna fritt marknadsförs på en medlemsstats territorium där sådana uttryck är förbjudna.
1. När en ursprungsbeteckning eller en geografisk beteckning registrerats i enlighet med denna förordning, skall ansökan om registrering av ett varumärke som svarar mot något av de fall som nämns i artikel 13 och som avser samma slags produkt, avslås om ansökningen ingivits efter dagen för det offentliggörande som avses i artikel 6.2.
Artikel 15
Kommissionen skall själv anta förslaget till åtgärder om detta har tillstyrkts av kommittén.
Artikel 16
1. Inom sex månader efter det att denna förordning har trätt i kraft, skall medlemsstaterna meddela kommissionen vilka hos dem skyddade beteckningarna eller, vad gäller medlemsstater som saknar sådant skyddssystem, vilka inarbetade beteckningar de önskar registrera i enlighet med denna förordning.
Artikel 18
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EEG) nr 1418/76 av den 21 juni 1976 om den gemensamma organisationen av marknaden för ris(3), senast ändrad genom förordning (EEG) nr 674/92(4), särskilt artikel 17.6 i denna, och
Av hänsyn till tydligheten bör förordning (EEG) nr 1124/77 upphöra att gälla och dess bestämmelser bör införas i den här förordningen.
Artikel 1
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
I kommissionens förordning (EEG) nr 1274/91(2), senast ändrad genom förordning (EEG) nr 3540/91(3), fastställs de tillämpningsföreskrifter som krävs för införandet av sådana handelsnormer.
De termer som används för livsmedelsindustrin bör harmoniseras.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fjäderfäkött och ägg.
" - värpdagen skall anges på ägg vilka levereras av en produktionsenhet som är belägen på samma ställe som förpackningsanläggningen och vilka inte förpackas i slutna behållare, i vilket fall de skall klassificeras och förpackas på värpdagen, eller, om värpdagen inte infaller på en arbetsdag, den första därpå följande arbetsdagen."
3. När datum som avses i denna artikel anges på ägg, och i fråga om värpdag även på förpackningen, skall en eller flera av de termer som anges i bilaga 1 användas.
- månaden, från 01 till 12."
- namn och adress avseende de ägglevererande producenterna, som skall registreras efter det att den behöriga myndigheten i medlemsstaten har gjort ett kontrollbesök, och
- insättningsdagen, åldern vid insättning och antalet värphönor uppdelade efter hönshus,
3 Ägg på vilka man avser ange värpdagen skall levereras till förpackningsanläggningar i slutna behållare, om inte produktionsenheten är belägen på samma ställe som förpackningsanläggningen. Leveranser av dessa ägg och av ägg på vilka produktionsföretaget redan har stämplat värpdagen, skall identifieras genom
Dessa uppgifter skall anges på behållaren och på de åtföljande dokumenten, som skall bevaras på förpackningsanläggningen i minst 6 månader.
- stämplas med värpdagen samma dag som de värps medan ägg som värps på annan dag än arbetsdag får stämplas den första därpå följande arbetsdagen tillsammans med de ägg som värps denna dag, varvid den första dagen som inte är arbetsdag skall anges, eller
Om dessa förpackningsanläggningar även får ägg från externa producenter på vilka man inte avser ange värpdagen, skall dessa ägg lagras och hanteras separat. Dagligt register skall föras över uppsamling eller mottagning och klassificering av sådana ägg.
- daglig mängd ägg och äggens viktklass,
4 Artikel 18 skall ändras på följande sätt:
- I punkt 1 skall det andra stycket utgå.
5 Artikel 22.2 c skall ersättas med följande text:
2. Om den banderoll eller etikett som avses i punkt 1 inte kan avlägsnas från förpackningen, skall banderollen eller förpackningen avlägsnas från försäljningsytan senast den sjunde dagen efter förpackningstillfället, varefter äggen skall förpackas på nytt.
Om det kontrollerade partiet omfattar färre ägg än 180, skall ovan angivna procentsatser fördubblas."
Denna förordning träder i kraft den 1 augusti 1992. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Vid en genomgång visade det sig att den tyska utgåvan av förordningen inte återger de bestämmelser som förvaltningskommittén hade fått på remiss. Den tyska utgåvan bör därför ges ut i en helt ny version.
(Berör endast den tyska utgåvan.)
RÅDETS BESLUT av den 8 februari 1993 om ingående av ett avtal om handel och ekonomiskt samarbete mellan Europeiska ekonomiska gemenskapen och Mongoliet (93/101/EEG)
med beaktande av kommissionens förslag,
Artikel 4
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
i samarbete med Europaparlamentet(2),
Det har visat sig önskvärt att samla in uppgifter om de beståndsdelar som används i kosmetiska produkter, så att alla frågor som gäller användningen av dem och de därmed sammanhängande åtgärderna på gemenskapsnivå kan prövas på ett sätt som särskilt syftar till att upprätta en gemensam nomenklatur för beståndsdelar i kosmetiska produkter. Insamlingen av dessa uppgifter kan underlättas om kommissionen genomför en inventering av sådana beståndsdelar. Denna inventering skall vara vägledande och inte syfta till att upprätta en begränsande förteckning över ämnen för användning i kosmetiska produkter.
I förebyggande syfte bör dock den behöriga myndigheten underrättas om tillverkningsplats och ges den information som är nödvändig för en snar och adekvat medicinsk behandling i händelse av betänkligheter.
Artikel 1
"1. Med kosmetisk produkt avses ämnen eller beredningar som är avsedda att appliceras på olika yttre partier av människokroppen (överhud, hår och hårbotten, naglar, läppar och yttre könsorgan) eller på tänder och slemhinnor i munhålan i uteslutande, eller huvudsakligt, syfte att rengöra eller parfymera dem eller förändra deras utseende och/eller korrigera kroppslukt och/eller skydda dem eller bibehålla dem i gott skick."
3. Följande led skall läggas till i artikel 4.1:
Kommissionen skall lämna en årlig rapport till Europaparlamentet och rådet om de framsteg som gjorts i utvecklingen, valideringen och det juridiska godkännandet av alternativa metoder som kan ersätta sådana som förutsätter djurförsök. Denna rapport skall innehålla exakta uppgifter om antal och slag av försök avseende kosmetika som utförts på djur. Medlemsstaterna skall vara skyldiga att samla in sådana uppgifter utöver den statistikinsamling som fastställs i direktiv 86/609/EEG om skydd av djur som används för försök och andra vetenskapliga ändamål. Kommissionen skall särskilt säkerställa att försöksmetoder, i vilka levande djur inte används, utvecklas, valideras och godkänns i lagstiftningen."
1. Senast den 14 december 1994 skall kommissionen, med det förfarande som fastställs i artikel 10, ha sammanställt en inventering av de beståndsdelar som används i kosmetiska produkter, med stöd särskilt av information som lämnats av kosmetikaindustrin.
2. Inventeringen skall innehålla uppgifter om
- då så är tillämpligt, begränsningar och villkor för användningen samt de varningstexter som skall förekomma i märkningen med hänvisning till bilagorna.
"1. Medlemsstaterna skall vidta alla de åtgärder som är nödvändiga för att försäkra sig om att kosmetiska produkter inte kan släppas ut på marknaden utan att följande information finns i outplånlig, lättläst och väl synlig skrift på behållaren och förpackningen. Den information som nämns i g behöver dock endast anges på förpackningen:"
7. Följande led f och g skall läggas till i artikel 6.1:
Följande skall dock inte betraktas som beståndsdelar:
- Material av vilket endast oundgängligen nödvändiga kvantiteter används som lösningsmedel eller som bärare av parfym och aromatiska blandningar.
Beståndsdelar skall identifieras med den generiska benämning som avses i artikel 7.2 eller, om sådan saknas, med någon av de benämningar som avses i artikel 5a.2, första strecksatsen.
"Om det på grund av storlek eller form är ogörligt att uppta de uppgifter som avses i d och g på en bipacksedel skall dessa uppgifter förekomma på en etikett, en tejp eller ett kort som bipackas eller fästs på den kosmetiska produkten.
"Dessutom skall i varje omnämnande av djurförsök klart anges om de utförda försöken gällde slutprodukten och/eller dess beståndsdelar."
11. Artikel 7.3 skall ersättas med följande:
12. Följande artikel skall införas:
a) Produktens kvalitativa och kvantitativa sammansättning. I fråga om parfymsammansättningar och parfymer: sammansättningens namn och kodnummer och uppgift om leverantören.
d) Bedömning av slutproduktens säkerhet för människors hälsa. Tillverkaren skall därvid beakta beståndsdelens allmänna toxikologiska profil, dess kemiska struktur och dess exponeringsgrad.
f) Tillgängliga uppgifter om icke önskvärda verkningar på människors hälsa som orsakas av användning av den kosmetiska produkten.
3. Den information som avses i punkt 1 skall finnas tillgänglig på den berörda medlemsstatens nationella språk eller på ett språk som utan svårighet förstås av de behöriga myndigheterna.
13. Artikel 8.2 skall ersättas med följande:
Artikel 2
Artikel 3
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
RÅDETS DIREKTIV 93/41/EEG av den 14 juni 1993 om upphävande av direktiv 87/22/EEG om tillnärmning av medlemsstaternas åtgärder vad gäller meddelande av försäljningstillstånd för högteknologiska läkemedel på marknaden, särskilt sådana som framställts genom bioteknologi
med beaktande av kommissionens förslag(1),
med beaktande av följande: Bestämmelserna i direktiv 87/22/EEG(4) har nu ersatts med bestämmelserna i rådets förordning (EEG) nr 2309/93 av den 22 juli 1993 om gemenskapsförfaranden för godkännande för försäljning av och tillsyn över humanläkemedel och veterinärmedicinska läkemedel samt om inrättande av en europeisk läkemedelsmyndighet(5) och i rådets direktiv 88/182/EEG av den 22 mars 1988 om ändring av direktiv 83/189/EEG om ett informationsförfarande beträffande tekniska standarder och föreskrifter(6).
Direktiv 87/22/EEG bör därför upphävas.
Artikel 1
Ansökningar om godkännande för försäljning, som före den 1 januari 1995 har förelagts Kommittén för farmaceutiska specialiteter eller Kommittén för veterinärmedicinska läkemedel enligt artikel 2 i direktiv 87/22/EEG och beträffande vilka den berörda kommittén inte har avgivit något yttrande före den 1 januari 1995, skall anses uppfylla bestämmelserna i förordning (EEG) nr 2309/93.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(2),
Den europeiska konventionen om skydd för slaktdjur godkändes på gemenskapens vägnar genom rådets beslut 88/306/EEG(5). Konventionens räckvidd är större än de befintliga gemenskapsbestämmelserna på området.
Vid tidpunkten för slakt eller avlivning bör djur besparas onödig smärta och lidande.
I den förklaring om djurskydd som är knuten till slutakten av Fördraget om Europeiska unionen anmodar konferensen Europaparlamentet, rådet, kommissionen och medlemsstaterna att vid utformning och införande av gemenskapslagstiftning om den gemensamma jordbrukspolitiken fullt ut ta hänsyn till djurens behov av välbefinnande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- djur som avlivas under kultur- eller sportarrangemang,
5. Bedövning: Varje metod som när den används på ett djur omedelbart försätter detta i ett tillstånd av medvetslöshet som varar tills döden inträder.
8. Behörig myndighet: Den centrala myndigheten i en medlemsstat som ansvarar för veterinärkontroller eller annan myndighet till vilken denna befogenhet har delegerats.
Djur skall skonas från all onödig upphetsning, smärta och lidande under förflyttning, uppstallning, fasthållning, bedövning, slakt eller avlivning.
Slakterier, dvs. lokaler och utrustning, skall vara konstruerade på ett sådant sätt att djuren skonas från onödig upphetsning, smärta och lidande.
a) förflyttas och, om nödvändigt, uppstallas i enlighet med bilaga A,
d) avblödas i enlighet med bilaga D.
Artikel 6
Artikel 7
Artikel 8
Artikel 9
Artikel 10
3. Dagsgamla överskottskycklingar enligt definitionen i artikel 2.3 i direktiv 90/539/EEG, och embryon i kläckningsavfall skall avlivas så snabbt som möjligt i enlighet med bilaga G.
Artikel 12
Artikel 13
b) Kommissionen skall vidare senast den 31 december 1995 överlämna en rapport till rådet, som utarbetats på grundval av ett yttrande från Vetenskapliga veterinärmedicinska kommittén, tillsammans med relevanta förslag beträffande användningen av
- varje annan vetenskapligt erkänd metod för bedövning eller avlivning.
i) nödvändig strömstyrka och varaktighet vid bedövning av de olika berörda arterna,
Artikel 14
2. De kontroller som avses i punkt 1 skall utföras i samarbete med den behöriga myndigheten.
Artikel 15
Artikel 16
3. a) Kommissionen skall anta de avsedda åtgärderna när de är förenliga med kommitténs yttrande.
Artikel 17
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar, inklusive sanktionsåtgärder, som är nödvändiga för att följa detta direktiv den 1 januari 1995. De skall genast underrätta kommissionen om detta.
3. Medlemsstaterna skall meddela kommissionen ordalydelsen i de viktigaste nationella bestämmelserna som de antar på det område som omfattas av detta direktiv.
KOMMISSIONENS FÖRORDNING (EEG) nr 752/93 av den 30 mars 1993 om tillämpningsföreskrifter för rådets förordning (EEG) nr 3911/92 om export av kulturföremål
med beaktande av rådets förordning (EEG) nr 3911/92 av den 9 december 1992(1) om export av kulturföremål, särskilt artikel 7 i denna,
För att säkerställa att de exportlicenser som föreskrivs i nämnda förordning är enhetliga är det nödvändigt att fastställa regler för upprättandet, utfärdandet och användningen av formulären. Det bör därför utarbetas en förlaga till en sådan licens.
AVSNITT I Formulär för licens
1. Formuläret skall tryckas på vitt träfritt skrivpapper som väger minst 55 gram per kvadratmeter.
4. Medlemsstaterna skall vara ansvariga
5. Formulären skall företrädesvis fyllas i på mekanisk eller elektronisk väg. Ansökan får emellertid fyllas i läsligt för hand; i det senare fallet skall det fyllas i med bläck och med tryckbokstäver. Oavsett vilken metod som används får formulären inte innehålla raderingar, överskrivna ord eller andra ändringar. AVSNITT II
1. Utan att det påverkar tillämpningen av punkt 3 skall en särskild exportlicens utfärdas för varje sändning av kulturföremål.
Artikel 5
- ett exemplar märkt nr 2 är avsett för innehavaren av licensen,
1. Den sökande skall fylla i fält 1, 3 -19 A och 21 och om nödvändigt 23 på ansökan och de andra exemplaren. Medlemsstaterna får emellertid föreskriva att endast ansökan behöver fyllas i.
3. De behöriga myndigheterna får för att utfärda en exportlicens kräva att de kulturföremål som skall exporteras visas upp.
Artikel 7
- Det exemplar som skall återsändas till den utfärdande myndigheten.
3. Det exemplar av formuläret som skall återsändas till den utfärdande myndigheten skall åtfölja sändningen till kontoret vid platsen för utförsel ur gemenskapen. Tullkontoret skall om nödvändigt fylla i fält 5 i formuläret och stämpla i fält 22 och återsända det till innehavaren av exportlicensen eller dennes representant för att formuläret skall kunna sändas tillbaka till den utfärdande myndigheten.
2. I fråga om ansökan om temporär export får de behöriga myndigheterna specificera den tidsfrist inom vilken kulturföremålen skall återimporteras till den utfärdande medlemsstaten.
Bestämmelserna i avsnitt IX i kommissionens förordning (EEG) nr 1214/92(2) och artikel 22.6 i bilaga 1 till Konventionen om ett gemensamt transiteringsförfarande som slöts den 20 maj 1987(3) mellan gemenskapen och EFTA-länderna skall gälla när varor som omfattas av denna förordning passerar genom ett EFTA-lands territorium vid förflyttning inom gemenskapen.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Enligt kommissionens förordning (EEG) nr 876/75 av den 3 april 1975 om den avgörande faktorn för utbetalning av för lin och hampa samt silkesodling(4), kommissionens förordning (EEG) nr 1426/86 av den 14 maj 1986 om den avgörande faktorn för rätt till stöd för privat lagring av lin- och hampfibrer(5) och artikel 15 i kommissionens förordning (EEG) nr 1201/89 av den 3 maj 1989 om tillämpningsföreskrifter för stödsystemet för bomull(6), senast ändrad genom förordning (EEG) nr 2328/92(7), fastställs de avgörande faktorerna för jordbruksomräkningskursen på grundval av kriterier och rättsliga bestämmelser som genomgående har ändrats i samband med den nya agromonetära ordning som infördes genom förordning (EEG) nr 3813/92. I kommissionens förordning (EEG) nr 1068/93 av den 30 april 1993 om närmare föreskrifter för fastställande och tillämpning av jordbruksomräkningskurserna(8) fastställs på grundval av de nya bestämmelserna de avgörande händelserna för jordbruksomräkningskurserna, bland annat de som gäller ovannämnda belopp.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för lin och hampa.
I artikel 15 i förordning (EEG) nr 1201/89 skall följande stycke läggas till:
Artikel 4
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I kommissionens förordning (EEG) nr 3824/92 av den 28 december 1992 om ändring av priser och belopp fastställda i ecu till följd av centralkursjusteringarna(2), senast ändrad genom förordning (EEG) nr 1663/93(3), fastställs förteckningen över de priser och belopp som från början av regleringsåret 1993/944, skall divideras med koefficienten 1,013088, som fastställs i kommissionens förordning (EEG) nr 537/93(4), ändrad genom förordning (EEG) nr 1331/93(5), som ett led i ordningen för automatisk avveckling av negativa monetära avvikelser. I enlighet med artikel 2 i förordning (EEG) nr 3824/92 skall de sänkta priserna och beloppen fastställas och anges för varje ifrågavarande sektor.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: I förordning (EEG) nr 1907/90(2) föreskrivs vissa handels-normer för ägg.
Det bör klargöras att valfria märkningar på äggförpackningar avsedda som reklam får innehålla symboler och syfta på såväl ägg som andra varor.
Artikel 1
"a) ägg till någon annan än uppsamlare, förpacknings-anläggningar, de marknader som avses i artikel 2.2 a, livsmedelsindustriföretag som godkänts i enlighet med direktiv 89/437/EEG och andra företag än livsmedelsindustrin."
"a) Datum för minsta hållbarhetstid 'bäst-före-datum`".
6. Artikel 10.1 e skall ersättas med följande:
"e) Kommentarer eller symboler avsedda att främja försäljningen av ägg eller andra varor, under förutsättning att dessa kommentarer eller symboler är utformade på ett sådant sätt att det inte är sannolikt att de vilseleder köparen."
9. Artikel 15 b ee skall ersättas med följande:
Denna förordning träder i kraft den 1 december 1993.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(),
Det är bara om de berörda parterna erkänner att systemet är berättigat som det kan ge önskat resultat.
Det krävs att de inblandade parterna inom fiskerinäringen tar på sig ett ökat ansvar för att se till att åtgärderna för bevarande och förvaltning av fiskeresurserna genomförs.
Det är av avgörande betydelse att medlemsstaterna samarbetar under inspektionerna av fiskeverksamheten ute till havs för att dessa skall bli så effektiva och ekonomiskt försvarbara som möjligt, särskilt under de inspektioner som företas i farvattnen utanför en medlemsstats jurisdiktion eller överhöghet.
Förvaltningen av fisket genom fastställande av TAC:er förutsätter en ingående kännedom om fångsternas sammansättning. En sådan kännedom behövs också för övriga förfaranden enligt förordning (EEG) nr 3760/92. Det kräver att befälhavaren på varje fiskefartyg för loggbok.
För att kunna undanta små fiskefartyg från skyldigheten att föra loggbok eller fylla i en landningsdeklaration, för vilka en sådan skyldighet skulle innebära en oproportionerlig börda i förhållande till deras fiskekapacitet, är det nödvändigt att varje medlemsstat kan kontrollera dessa fartygs verksamhet genom att införa en provtagningsplan.
För att säkerställa att alla de utnyttjade resurserna bevaras och förvaltas kan bestämmelserna om loggbok, landnings- och försäljningsdeklarationer samt upplysningar om omlastningar och registrering av fångster utvidgas till att omfatta sådana bestånd som inte omfattas av någon TAC eller kvot.
Om det finns nätredskap med olika maskstorlek ombord kan det inte säkert garanteras att bestämmelserna om hur fiskeredskapen får användas följs om de inte blir föremål för ytterligare kontroll. För vissa former av fiske kan det vara lämpligt att införa speciella regler som till exempel ennätsregeln.
Om de ansvariga för fiskefartygen inte följer bestämmelserna i denna förordning bör dessa fartyg bli föremål för ytterligare kontroll med hänsyn till bevarandet.
Det är nödvändigt att fastställa allmänna regler så att gemenskapens inspektörer som utsetts av kommissionen kan se till att gemenskapsbestämmelserna tillämpas enhetligt och granska de kontroller som gjorts av medlemsstaternas behöriga myndigheter.
Om en landningsmedlemsstat inte effektivt beivrar oegentligheter kommer det att försvaga flaggmedlemsstatens möjligheter att se till att föreskrifterna för bevarande och förvaltning av fiskeresurserna följs. Det är därför nödvändigt att fastställa bestämmelser om att olovliga fångster skrivs av från landningsmedlemsstatens kvot, om denna stat underlåter att vidta effektiva åtgärder.
Det bör säkerställas att de uppgifter som samlas in inom ramen för denna förordning behandlas konfidentiellt.
Det är nödvändigt att fastställa en övergångsperiod för genomförandet av särbestämmelserna i vissa artiklar för att de behöriga myndigheterna i medlemsstaterna skall kunna införa och anpassa sina förfaranden till den nya förordningens krav.
- åtgärderna för bevarande och förvaltning av fiskeresurserna,
samt vissa bestämmelser om hur verkningsfulla de sanktioner bör vara som skall tillämpas om ovan nämnda åtgärder inte genomförs.
1. För att säkerställa att alla gällande föreskrifter om åtgärder för bevarande och kontroll följs skall varje medlemsstat inom sitt territorium och de marina farvatten som lyder under dess överhöghet eller jurisdiktion övervaka fisket och den därmed förbundna verksamheten. Medlemsstaten skall inspektera fiskefartygen och undersöka all verksamhet rörande landning, försäljning, transport och lagring av fisk samt registrering av landningar och försäljning, och kan på så sätt granska tillämpningen av denna förordning.
3. Varje medlemsstat skall kontrollera sina fartygs verksamhet utanför gemenskapens fiskezon, om en sådan kontroll krävs för att säkerställa att de gemenskapsbestämmelser som gäller i dessa farvatten efterlevs.
1. För att åstadkomma större effektivitet i övervakningen av fiskeverksamheten skall rådet före den 1 januari 1996 i enlighet med det förfarande som fastställs i artikel 43 i fördraget besluta om i vilken utsträckning och när ett system bör införas för fortlöpande kontroll av gemenskapens fiskefartygs position från en land- eller satellitbaserad basstation med dataöverföring via satellit.
3. När de pilotprojekt som avses i punkt 2 genomförs skall den medlemsstat vars flagg fartyget för eller i vilken fartyget är registrerat vidta nödvändiga åtgärder för att säkerställa att de data som översänds till eller inhämtas från dess fiskefartyg registreras i maskinläsbar form, oberoende av i vilka vatten fartygen fiskar eller i vilken hamn de befinner sig.
Medlemsstaterna skall när de utför de uppgifter som anförtrotts dem se till att de i artikel 2 angivna bestämmelserna och åtgärderna respekteras. De skall dessutom vid inspektionen undvika att göra onödiga ingrepp i den normala fiskeverksamheten. De skall också se till att ingen diskriminering sker med avseende på de sektorer och fartyg som tas ut för inspektion.
I enlighet med förfarandet i artikel 36 kan tillämpningsföreskrifter antas för artiklarna 2, 3 och 4, speciellt med avseende på
c) det förfarande som inspektörer som har gått ombord på ett fiskefartyg skall följa när de inspekterar fartyget, dess fiskeredskap eller fångster,
f) utfärdande av intyg för fiskefartygens egenskaper avseende fiskeaktiviteter,
Artikel 6
3. Befälhavarna på gemenskapens fiskefartyg skall i loggböckerna skriva in vilka mängder som fångats i havet, datum och plats för dessa fångster samt de i punkt 2 avsedda arterna. De mängder som kastats överbord kan registreras i uppskattningssyfte.
6. Varje medlemmstat skall genom stickprovskontroller kontrollera verksamheten hos de fiskefartyg som är undantagna från de krav som anges i punkterna 4 och 5 för att säkerställa att dessa fartyg följer gällande gemenskapsbestämmelser.
8. Närmare bestämmelser skall antas för tillämpningen av denna artikel enligt det förfarande som anges i artikel 36, i vissa speciella fall med en annan geografisk grundval än den statistiska ICES-rektangeln.
- landningsplatsen eller landningsplatserna och den beräknade ankomsttiden,
3. Kommissionen kan enligt det förfarande som anges i artikel 36 undanta vissa kategorier av fiskefartyg inom gemenskapen från den skyldighet som avses i punkt 1 under en begränsad tid, som kan förnyas, eller fastställa en annan anmälningsfrist, där hänsyn bland annat skall tas till avståndet mellan fiskebankarna, landningsplatserna och de hamnar i vilka fartygen ifråga är registrerade eller förtecknade.
2. Rådet kan med kvalificerad majoritet på förslag av kommissionen besluta om att utsträcka den skyldighet som avses i punkt 1 till sådana fartyg som har en största längd av mindre än 10 m. Rådet kan också med kvalificerad majoritet på förslag av kommissionen besluta om undantag från skyldigheten i punkt 1 för vissa kategorier av fartyg med en största längd av minst 10 m, vilka bedriver viss typ av fiskeverksamhet.
4. Tillämpningsföreskrifter för denna artikel skall antas i enlighet med det förfarande som fastställs i artikel 36.
2. Om den första saluföringen av de fiskeprodukter som landats i en medlemsstat inte sker på det sätt som fastställs i punkt 1 får köparen inte föra bort de landade fiskeprodukterna innan en avräkningsnota lämnats in till de behöriga myndigheterna eller andra godkända organ i den medlemsstat på vars territorium saluföringen ägt rum. Köparen är ansvarig för riktigheten av de uppgifter enligt punkt 3 som avräkningsnotan innehåller.
- Pris och mängd av varje art vid första försäljningstillfället och, i förekommande fall, beroende på de olika arternas storlek eller vikt, kvalitet, produktform och färskhet.
- Dag och plats för försäljningen.
- Namnet på fartygets ägare eller befälhavare.
6. De behöriga myndigheterna skall behålla ett exemplar av varje avräkningsnota under en tid av ett år räknat från början av det år som följer på året för registreringen av den information som översänts till de behöriga myndigheterna.
8. En köpare som köper produkter som inte saluförs vidare utan endast används för privat konsumtion skall undantas från kraven i punkt 2.
1. a) De fiskefartyg som för ett tredje lands flagg eller är registrerade i ett tredje land, och som har tillstånd att bedriva fiske i sådana marina farvatten som lyder under en medlemsstats överhöghet eller jurisdiktion, skall föra loggbok, i vilken den i artikel 6 angivna informationen skall införas.
Befälhavaren får inte landa fångster om medlemsstatens behöriga myndigheter inte bekräftat mottagandet av förhandsanmälan.
3. Punkterna 1 och 2 skall gälla utan att de påverkar tillämpningen av de fiskeavtal som ingåtts mellan gemenskapen och vissa tredje länder.
- omlastar valfria fångstmängder ur ett bestånd eller en grupp av bestånd inom en TAC eller kvot till ett annat fartyg, nedan kallat "mottagarfartyg", oberoende av omlastningsplatsen, eller
2. Senast 24 timmar innan en omlastning eller serie omlastningar som äger rum i en hamn eller i sådana marina farvatten som lyder under en medlemsstats överhöghet eller jurisdiktion inleds, eller när de avslutats, skall mottagarfartygets befälhavare underrätta denna medlemsstats behöriga myndigheter om storleken på de fångster ur ett bestånd eller en grupp av bestånd som omfattas av en TAC eller en kvot, vilka befinner sig ombord på detta fartyg.
Befälhavaren på mottagarfartyget skall också förvara uppgifterna om vilka fångstmängder ur ett bestånd eller en grupp av bestånd inom en TAC eller kvot som mottagarfartyget lastat om till ett tredje fartyg, samt underrätta ovannämnda behöriga myndigheter om denna omlastning minst 24 timmar innan den äger rum. Efter omlastningen skall befälhavaren underrätta nämnda myndigheter om vilka mängder som lastats om.
4. Punkterna 2 och 3 skall även tillämpas på ett mottagarfartyg som för ett tredje lands flagg eller är registrerat i ett tredje land.
Artikel 13
a) försändelsens ursprung (fartygets namn och distriktsbeteckning),
3. Varje transportföretag skall se till att det dokument som avses i punkt 1 innehåller minst alla de uppgifter som anges i punkt 2.
b) Dokumentet enligt punkt 1 ersätts med en kopia av dokumentet T 2 M, som anger de transporterade mängdernas ursprung.
7. Medlemsstaterna skall samordna sin kontrollverksamhet för att kontrollen skall bli så effektiv och ekonomisk som möjligt. Medlemsstaterna skall därför särskilt övervaka de varutransporter som tilldragit sig deras uppmärksamhet och som de misstänker strider mot gemenskapens föreskrifter.
2. Om den första saluföringen av landade fångster inte sker genom offentlig auktion i enlighet med bestämmelserna i artikel 9.2, skall medlemsstaterna se till att auktionsinrättningarna eller de andra organ som de bemyndigat erhåller information om ifrågavarande mängder.
Artikel 15
Varje medlemsstat skall ge kommissionen en prognos över kvotutnyttjandet med angivande av det datum när kvoten beräknas vara uttömd för de arter som tagits från fiskefartyg som för denna medlemsstats flagg eller är registrerade där, när det bedöms att fångsterna av dessa arter uppgår till 70 % av den kvot, tilldelning eller andel som den staten förfogar över.
3. Om kommissionen finner att en medlemsstat inte hållit den frist för överföring av uppgifter om månatliga fångster som fastställs i punkt 1 kan den fastställa ett datum när fångsterna ur ett bestånd eller en grupp av bestånd, som omfattas av en kvot eller någon annan form av mängdbegränsning, och som tas från fiskefartyg som för denna medlemsstats flagg eller är registrerade i denna medlemsstat, skall anses utgöra 70 % av den kvot, tilldelning eller andel som denna medlemsstat förfogar över, samt ett datum för när kvoten, tilldelningen eller andelen skall anses vara uttömd.
1. Utan att det påverkar tillämpningen av artikel 15 skall medlemsstaterna på den berörda medlemsstatens begäran lämna upplysning om de landningar, utbjudningar till försäljning eller omlastningar av fiskeprodukter som äger rum i deras hamnar eller i de farvatten som lyder under deras jurisdiktion från sådana fiskefartyg som för denna medlemsstats flagg eller är registrerade i denna, och som omfattar fisk ur ett bestånd eller en grupp av bestånd från en kvot som tilldelats denna medlemsstat.
Artikel 17
- Fiskefartygen skall ha en loggbok ombord, i vilken befälhavarna registrerar sina fångster.
3. Bestämmelserna i punkterna 1 och 2 skall tillämpas utan att det påverkar tillämpningen av bestämmelserna i de fiskeavtal som slutits mellan gemenskapen och tredje land, samt de internationella konventioner som gemenskapen anslutit sig till.
2. För sådana fångster som tas i ett tredje lands farvatten skall den information som lämnas i enlighet med punkt 1 anges per tredje land och bestånd med hänvisning till det minsta statistiska område som fastställts för ifrågavarande fiskeverksamhet.
Artikel 19
Medlemsstaterna får upprätta decentraliserade databaser på villkor att dessa databaser och de metoder som används för insamling och registrering av data är standardiserade, så att de är kompatibla med varandra på en medlemsstats hela territorium.
5. Inom tolv månader efter det att denna förordning trätt i kraft skall varje medlemsstat lämna in en rapport till kommissionen, i vilken det beskrivs hur uppgifterna samlas in och kontrolleras och hur tillförlitliga de är. Kommissionen skall i samarbete med medlemsstaterna göra en sammanfattning av rapporterna, som den skall delge medlemsstaterna.
1. Alla fångster som bevaras ombord på ett fiskefartyg inom gemenskapen skall vara i överensstämmelse med den artsammansättning som fastställs för nätredskapen ombord på fartyget i fråga i rådets förordning (EEG) nr 3094/86 av den 7 oktober 1986 om vissa tekniska åtgärder för bevarande av fiskeresurserna().
b) Nätredskapen som finns på däck eller ovanför däck skall vara säkert fastgjorda vid någon del av överbyggnaden.
3. Trots bestämmelserna i punkterna 1 och 2 kan rådet på grundval av en rapport utarbetad av kommissionen på dennas förslag med kvalificerad majoritet besluta att
Artikel 21
3. Efter en anmälan i enlighet med punkt 2, eller på eget initiativ, skall kommissionen på grundval av tillgänglig information fastställa ett datum för när de fångster ur ett bestånd eller en grupp av bestånd som omfattas av en TAC, kvot eller någon annan form av mängdbegränsning, som de fiskefartyg tagit som för en medlemsstats flagg eller är registrerade i en medlemsstat, skall anses ha förbrukat den kvot, tilldelning eller andel som står till denna medlemsstats eller, eventuellt, gemenskapens förfogande.
4. När kommissionen i enlighet med punkt 3 första stycket har stoppat fiskeverksamheten på grund av att den TAC, kvot, tilldelning eller andel som står till gemenskapens förfogande antas vara förbrukad, och det visar sig att en medlemsstat i själva verket inte har förbrukat den kvot, tilldelning eller andel som den förfogar över av ifrågavarande bestånd eller grupp av bestånd, skall följande bestämmelser tillämpas.
Artikel 22
Artikel 23
- Överfiskets omfång.
Artikel 24
1. Varje medlemsstat skall anta bestämmelser för att kontrollera att de mål som avses i artikel 24 uppfylls. Den skall därför företa tekniska kontroller, särskilt på följande områden:
c) Begränsning av vissa fiskefartygs verksamhet.
2. Utan att det påverkar tillämpningen av artikel 169 i fördraget kan kommissionen, om den finner att en medlemsstat inte följt bestämmelserna i punkt 1, lägga fram förslag till rådet om att anta lämpliga allmänna åtgärder. Rådet skall fatta beslut med kvalificerad majoritet.
a) fiskefartygens maskinstyrka,
d) fiskeredskapens karakteristika och deras antal per fiskefartyg.
1. För att underlätta den kontroll som avses i artikel 25 skall medlemsstaterna införa ett system för giltighetskontroll, som särskilt skall omfatta en korsvis kontroll av uppgifterna om fiskeflottans kapacitet och verksamhet i bl.a.
- gemenskapens förteckning över fiskefartyg, som avses i kommissionens förordning (EEG) nr 163/89().
4. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som anges i artikel 36.
2. Dessa kontroller skall gälla de tekniska aspekterna av tillämpningen av
- återtagande av produkter från marknaden för andra ändamål än mänsklig konsumtion,
3. Medlemsstaterna skall ge kommissionen upplysningar om utförda kontroller, behöriga kontrollmyndigheter, konstaterade överträdelser och vilka åtgärder som dessa föranlett.
Artikel 29
2. Närhelst kommissionen anser det nödvändigt kan dess inspektörer närvara vid de nationella tillsynsmyndigheternas kontroller och inspektioner. Inom ramen för detta uppdrag skall kommissionen upprätta lämpliga kontakter med medlemsstaterna för att om möjligt utarbeta ett inspektionsprogram som kan godtas av båda parter.
b) Om förhållandena på platsen gör det omöjligt att genomföra den inspektion och kontroll som planerats i det ursprungliga inspektionsprogrammet skall kommissionens inspektörer i samarbete med den behöriga tillsynsmyndigheten, och med dess samtycke, ändra den ursprungligen planerade inspektionen och kontrollen.
3. Kommissionen kan vid behov, särskilt om gemenskapens inspektörer i enlighet med punkt 2 avslöjat att oegentligheter kan ha begåtts vid tillämpningen av denna förordning, anmoda medlemsstaterna att lämna närmare uppgifter om vilket inspektions- och kontrollprogram som de behöriga nationella myndigheterna planerat eller fastställt för en viss period och fiskeverksamhet samt vissa områden. Efter mottagandet av denna information skall kommissionens inspektörer, om denna anser det nödvändigt, göra egna inspektioner för att granska hur en medlemsstats behöriga myndigheter genomfört detta program.
4. Vid inspektioner från luften, till havs eller till lands, får de behöriga inspektörerna inte företa någon kontroll av fysiska personer.
Artikel 30
Den eller de berörda medlemsstaterna skall informera kommissionen om undersökningens förlopp och resultat och lämna kommissionen en kopia av undersökningsrapporten och de centrala bevismaterial som legat till grund för utarbetandet av rapporten.
Om det enligt nationell lagstiftning är förbehållet vissa i lagen angivna tjänstemän att utföra vissa handlingar på det straffrättsliga området skall kommissionens tjänstemän avhålla sig från att medverka i dessa handlingar. De skall särskilt avhålla sig från att delta i husrannsakningar och formella förhör av personer enligt nationell straffrätt. De skall dock ha tillträde till den information som fås på detta sätt.
1. Medlemsstaterna skall se till att lämpliga åtgärder vidtas mot ansvariga fysiska eller juridiska personer, även sådana förvaltnings- eller straffrättsliga åtgärder som överensstämmer med nationell lagstiftning, när det, särskilt efter en kontroll eller inspektion som utförts enligt denna förordning, står klart att den gemensamma fiskeripolitikens bestämmelser inte följts.
- böter,
- tillfällig indragning av licensen,
Artikel 32
Vilken fiskmängd som skall skrivas av från den medlemsstatens kvot skall fastställas på det sätt som anges i artikel 36, när kommissionen har hört de två berörda medlemsstaterna.
1. Medlemsstaternas behöriga myndigheter skall omgående i enlighet med den nationella lagstiftningens förfarande till flagg- eller registreringsmedlemsstaten anmäla alla överträdelser av de gemenskapsbestämmelser som avses i artikel 1, med angivande av det berörda fartygets namn och distriktsbeteckning, befälhavarens och ägarens namn, omständigheterna kring överträdelsen och de förvaltnings- eller straffrättsliga påföljderna, eller andra åtgärder som vidtagits samt alla slutgiltiga avgöranden i samband med sådana överträdelser. I speciella fall skall medlemsstaterna efter anmodan överlämna denna information till kommissionen.
Artikel 34
2. Medlemsstaterna skall regelbundet underrätta kommissionen om resultaten av de inspektioner eller kontroller som görs med stöd av denna förordning, särskilt vilken mängd och typ av överträdelse som konstaterats och vilka åtgärder som vidtagits. Medlemsstaterna skall på kommissionens anmodan till denna anmäla vilka bötesbelopp som tillämpats i de konkreta fallen av överträdelse.
Medlemsstaterna skall före den 1 juni varje år överlämna en rapport till kommissionen om tillämpningen av denna förordning under föregående kalenderår; denna skall innehålla en utvärdering av de tekniska och mänskliga insatserna och ange vilka åtgärder som skulle kunna bidra till att mildra de brister som eventuellt kunnat konstateras. På grundval av medlemsstaternas rapporter och de egna observationerna skall kommissionen sammanställa en årlig rapport och till varje medlemsstat överlämna de delar av rapporten som berör denna. Efter att ha tagit vederbörlig hänsyn till medlemsstaternas svar skall kommissionen offentliggöra hela rapporten med medlemsstaternas svar och eventuella förslag till åtgärder i syfte att avhjälpa de konstaterade bristerna.
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen, varvid medlemsstaternas röster skall vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
Artikel 37
Uppgifterna i punkt 1 skall bara föras vidare om de är så införlivade med andra uppgifter att de berörda fysiska eller juridiska personerna inte direkt eller indirekt kan identifieras.
5. Uppgifterna i punkt 1 får inte användas för något annat ändamål än det som anges i denna förordning, om inte de myndigheter som lämnar dem uttryckligen samtycker till det, och gällande bestämmelser i den medlemsstat vars myndighet tar emot uppgifterna inte förbjuder en sådan användning eller utlämning av uppgifter.
7. Varje gång en medlemsstat meddelar kommissionen att den efter en slutförd undersökning funnit att en fysisk eller juridisk person, vars namn meddelats den i kraft av bestämmelserna i denna förordning, inte varit inblandad i en överträdelse, skall kommissionen omedelbart underrätta alla dem som den lämnat ut den berörda personens namn till om utgången av undersökningen eller de rättsliga åtgärderna. Personen ifråga skall inte längre behandlas som om han eller hon vore inblandad i de oegentligheter som det första meddelandet innehöll uppgift om. De uppgifter som bevaras på ett sådant sätt att den berörda personen kan identifieras skall omgående förstöras.
10. De upplysningar som tas emot inom ramen för denna förordning skall på begäran ställas till de berörda fysiska eller juridiska personernas förfogande.
De nationella åtgärder som avses i första stycket skall anmälas till kommissionen i enlighet med artikel 2.2 i rådets förordning (EEG) nr 101/76 av den 19 januari 1976 om en gemensam strukturpolitik för fiskerisektorn().
2. Hänvisningar till den i punkt 1 upphävda förordningen skall anses som hänvisningar till denna förordning.
Medlemsstaterna skall fram till den 1 januari 1996 undantas från skyldigheten att tillämpa bestämmelserna i artiklarna 9, 15 och 18 i fråga om dataöverföring av avräkningsnotor och registrering av landningar.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas avseende den gemen-samma jordbrukspolitiken(2), särskilt artikel 6 i denna, och
Tillämpningsföreskrifterna bör också omfatta fastställande av ansökningstid för stödet, vilka uppgifter ansökan minst bör innehålla, den behöriga myndighetens tidsgränser för behandling av ansökan och utbetalning av stöd, samt anmälan till kommissionen om utbetalt stöd. Det bör också fastställas bestämmelser om den kontroll som är nödvändig för att säkerställa att stödordningen tillämpas på ett korrekt sätt, och om vilka åtgärder som skall vidtas vid underlåtenhet att uppfylla bestämmelserna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Fram till slutet av 1994 skall stödet dock även betalas ut till alla biodlare som har minst tio fasta producerande bikupor som är registrerade hos den behöriga myndigheten.
- Förbättring av saluföringen genom införande av teknik, mekaniserad slungning, rening och filtrering, samt yrkesutbildning.
2. Sammanslutningarna av honungsproducenter skall förelägga den behöriga myndigheten sina program för god-kännande. Myndigheten skall, senast två månader efter prog-rammets inlämnande, besluta om godkännande eller avslag, efter att i förekommande fall ha anmodat om nödvändiga förändringar.
För år 1993 kan emellertid stödansökningar lämnas in senast den 15 december 1993.
- Antal fasta bikupor i produktion och det registrerings-nummer som den behöriga myndigheten tilldelat dem.
Artikel 4
Artikel 5
- Antal bikupor för vilka producentsammanslutningar och individuella biodlare ansökt om och beviljats stöd.
- Antal oegentligheter som konstaterats och de bikupor som de gäller.
1. Grekland skall, genom kontroller på plats, säkerställa att uppgifterna som lämnats i stödansökan är korrekta, samt att villkoren för utbetalning av stöd uppfylls.
2. Om stöd måste indrivas på grund av oegentligheter som kan tillskrivas sökanden, oavsett om dessa orsakats avsiktligt eller genom grov försumlighet, skall den behöriga myndigheten driva in utbetalda belopp med en höjning på 20 % samt ränta enligt punkt 1. Sökanden skall inte vara berättigad till stöd det följande året.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 84.2 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
Denna förordning inskränker inte tillämpningen av artiklarna 85 och 86 i fördraget.
Huvuddelen av dessa resor är paketresor eller kombinerade produkter, där lufttransport bara utgör en del i hela produkten.
Alla frågor som rör användningen av datoriserade bokningssystem för alla typer av lufttransportprodukter bör behandlas i en och samma förordning, som beslutas av rådet.
De lufttrafikföretag som använder ett datoriserat bokningssystem i sina egna klart markerade kontor eller diskar bör inte omfattas av bestämmelserna om primär textbild.
Att de datoriserade bokningssystemen är konkurrensmässigt neutrala i förhållande till lufttrafikföretag måste säkerställas vad gäller likhet i funktion och datasäkerhet, särskilt genom lika tillträde till funktioner, information/data och gränssnitt samt en klar åtskillnad mellan lufttrafikföretagens egna tjänster och distributionstjänster.
I konsumenternas intresse är det önskvärt att en primär textbild ges för varje transaktion som begärs av en konsument.
I konsumenternas intresse är det önskvärt att klargöra att en flygning eller kombination av flygningar inte skall visas mer än en gång på den primära textbilden, utom i de fall där genom ett konsortium eller någon annan form av uppgörelse varje lufttrafikföretag som bedriver lufttrafik tar på sig separat ansvar för erbjudandet och försäljningen av lufttransportprodukter på de berörda flygningarna.
Artikel 1
P systemleverantörens status eller nationalitet,
Artikel 2
b) kombinerad lufttransportprodukt: en på förhand avtalad kombination av en separat lufttransportprodukt med andra tjänster som inte är bitjänster till lufttransport, och som erbjuds till försäljning och/eller säljs till ett totalpris.
P Den utförs med luftfartyg för befordran av passagerare eller passagerare och gods och/eller post mot vederlag på ett sådant sätt att det på varje flygning finns platser att köpa för enskilda personer (antingen direkt av lufttrafikföretaget eller av dess auktoriserade agenter).
2. med flygningar som är så regelbundna eller täta att de utgör en igenkännlig planmässig serie.
P tidtabeller,
P tjänster i samband med flygbefordran,
P att utställa biljetter
h) systemleverantör: varje företag och dess filialer som har ansvaret för driften eller marknadsföringen av ett datoriserat bokningssystem.
P rättigheten att förfoga över alla eller en del av företagets tillgångar,
l) abonnent: en person eller ett företag som inte är ett deltagande lufttrafikföretag och som enligt avtal eller annan överenskommelse med en systemleverantör använder ett datoriserat bokningssystems distributionstjänster för försäljning av lufttransportprodukter.
o) restid: skillnaden mellan tidtabellsenlig avgångs- och ankomsttid.
knyta oskäliga villkor till ett avtal med ett deltagande lufttrafikföretag,
c) Ett deltagande lufttrafikföretag skall ha rätt att säga upp sitt avtal med en systemleverantör med en uppsägningstid som inte behöver överstiga sex månader, dock att den tidigast får löpa ut vid utgången av det första avtalsåret.
2. Följande artikel skall läggas till:
1. b) Moderföretaget skall inte vara förpliktat att acceptera några kostnader i samband med detta utom för återgivande av den information som skall ges och för accepterade bokningar.
3. Artikel 4 skall ersättas med följande:
3. En systemleverantör skall säkerställa att dess distributionstjänster är avskilda på ett klart och verifierbart sätt från varje lufttrafikföretags privata tjänster rörande platstillgång, företagsledning och avsättning. Åtskillnaden får ske antingen logiskt genom mjukvara eller fysiskt på ett sådant sätt att varje förbindelse mellan distributionstjänsterna och de privata tjänsterna bara uppnås genom ett gränssnitt mellan två tillämpningar. Oavsett metoden för åtskillnad skall ett sådant gränssnitt göras tillgängligt för alla moderföretag och deltagande lufttrafikföretag utan diskriminering samt ge lika behandling avseende procedurer, protokoll, inmatning och utmatning. När relevanta och allmänt accepterade standarder för lufttransportsektorn finns tillgängliga skall systemleverantörerna erbjuda tjänster som är kompatibla med dessa."
2. a) En systemleverantör skall via sitt datoriserade bokningssystem tillhandahålla en eller flera primära textbilder för varje enskild transaktion som visar data som inlevererats av deltagande lufttrafikföretag, om tidtabeller, biljettpriser och tillgången på platser för enskilda köpare på ett klart och tillräckligt omfattande sätt som inte är diskriminerande eller partiskt, i synnerhet vad gäller den ordning i vilken informationen presenteras.
1. d) Ordningsföljden mellan olika flygmöjligheter på den primära textbilden skall vara den som framgår av bilagan.
4. Information om kombinerade produkter avseende bl.a. vem som organiserar resan, platstillgång och priser skall inte visas i den primära textbilden.
1. Följande bestämmelser skall styra tillgängligheten av den information i form av statistik eller av annat slag, som en systemleverantör erbjuder från sitt datoriserade bokningssystem:
i) Att uppgifterna erbjuds med samma skyndsamhet och på ett icke-diskriminerande sätt till alla deltagande lufttrafikföretag, inklusive moderföretag.
2. Personlig information om en passagerare som kommer från ett datoriserat bokningssystem får bara med passagerarens medgivande göras tillgänglig för andra som inte är berörda av transaktionen.
5. Efter att ha mottagit den utförliga beskrivningen av de tekniska och administrativa åtgärder som vidtagits av systemleverantören, skall kommissionen inom tre månader fatta beslut om huruvida åtgärderna är tillräckliga för att uppfylla säkerhetskraven enligt denna artikel. Om så inte är fallet får kommissionen i sitt beslut tillämpa artikel 3a.2. Kommissionen skall genast informera medlemsstaterna om ett sådant beslut. Om rådet, på begäran av en medlemsstat, inte inom två månader efter kommissionens beslut beslutar annorlunda, skall kommissionens beslut träda i kraft."
7. I artikel 7 skall följande punkt läggas till:
1. Ett moderföretag får inte till en abonnents användning av något visst datoriserat bokningssystem direkt eller indirekt knyta någon provision eller annan förmån eller någon avskräckande åtgärd för att sälja företagets lufttransportprodukter som är tillgängliga på dess flygningar.
9. Artikel 9.4, 9.5 och 9.6 skall ersättas med följande:
"4. b) Med förbehåll för punkt 2 skall leverans av teknisk utrustning inte omfattas av villkoren enligt a.
b) att abonnenten inte behandlar det material som levereras av de datoriserade bokningssystemen på ett sätt som skulle leda till att konsumenterna får oriktig, vilseledande eller diskriminerande information.
"1. De avgifter som begärs av en systemleverantör får inte vara diskriminerande och skall vara rimligt strukturerade och stå i ett rimligt förhållande till anskaffningskostnaden för den tjänst som tillhandahålls och utnyttjas och skall i synnerhet vara desamma för samma servicenivå.
P Passagerarens namn.
P Ortkod.
P Resdatum.
P Bokningsnummer (PNR-nummer).
Ett deltagande lufttrafikföretag skall erbjudas möjligheten att bli informerat när det sker en bokning/transaktion för vilken en bokningsavgift kommer att debiteras. Om företaget väljer att bli informerat skall det erbjudas möjligheten att kunna annullera en sådan bokning/transaktion, såvida den inte redan har accepterats.
"Artikel 21
"Artikel 21a
13. Artikel 22 skall ersättas med följande:
2. De som har rättigheter enligt artikel 3.4, 4a, 6 och 21 a får inte avsäga sig dessa rättigheter genom avtal eller på annat sätt."
1. Rådet skall besluta om revidering av denna förordning senast den 31 december 1997 på grundval av ett förslag från kommissionen vilket skall överlämnas senast den 31 mars 1997 tillsammans med en redogörelse för tillämpningen av denna förordning.
Artikel 2
3. Skyldigheten enligt punkt 9 c i bilagan att visa anslutande flygtrafik med en linje per sträcka skall tillämpas från och med den 1 januari 1995.
VERKSTÄLLANDE KOMMITTÉN HAR FATTAT DETTA BESLUT
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av kommissionens förslag, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Texten till tilläggsprotokollet bifogas detta beslut.
Rådets ordförande skall på Europeiska gemenskapens vägnar göra den anmälan som fastställs i artikel 8 i tilläggsprotokollet.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Heartwater, babesios och anaplasmos, som överförs av smittbärande insekter, förekommer i de franska utomeuropeiska departementen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"- Heartwater, som överförs av smittbärande insekter i de franska utomeuropeiska departementen,
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Genom artikel 1 i direktiv 89/556/EEG utesluts från direktivets räckvidd embryon som är resultatet av vissa tekniker. Handel eller import med embryon som skall underkastas tekniker som innebär att zona pellucida genombryts, och med sådana som är resultatet av befruktning in vitro får ske under förutsättning att de uppfyller kraven i direktiv 89/556/EEG samt vissa kompletterande skyddsåtgärder.
Artikel 1
Detta beslut skall tillämpas från och med den 1 mars 1994.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, och
Enligt vad som avses i artikel 209a i fördraget skall medlemsstaterna vidta samma åtgärder för att motarbeta bedrägerier som riktar sig mot gemenskapens finansiella intressen som de vidtar för att motarbeta bedrägerier som riktar sig mot deras egna finansiella intressen. Därför måste de med kommissionens hjälp samordna sina insatser för att skydda gemenskapens finansiella intressen och motarbeta bedrägerier.
De befintliga kommittéernas arbetsuppgifter är begränsade till särskilda områden. Dessa kommittéer ersätts inte. Det finns dock behov av att få en samlad överblick över problematiken när det gäller bedrägerier som riktar sig mot gemenskapens budget. Därför bör en kommitté inrättas som kan behandla hela bedrägeriproblematiken.
Artikel 2
3. Arbetsgrupper kan inrättas för att underlätta kommitténs arbete.
RÅDETS BESLUT av den 19 april 1994 om en av rådet enligt artikel J 3 i Fördraget om den Europeiska unionen beslutad gemensam åtgärd till stöd för fredsprocessen i Mellanöstern (94/276/GUSP)
med beaktande av de allmänna riktlinjer som utfärdades av Europeiska rådet den 29 oktober 1993,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- delta i de internationella arrangemang som parterna kommer överens om för att säkerställa fred inom ramen för den process som startades i Madrid,
b) Europeiska unionen skall
- överväga andra sätt att bidra till regionens utveckling.
- fortsätta att rikta demarscher till de arabiska staterna i syfte att få till stånd ett slut på bojkotten mot Israel,
Rådet skall i enlighet med relevanta gemenskapsförfaranden behandla de förslag som kommissionen lägger fram om
Artikel 3
b) presidiet i nära samverkan med kommissionen underlätta samordningen genom utbyte av information mellan medlemsstaterna om deras bilaterala bistånd,
Europeiska unionen skall på begäran av parterna medverka till att det palestinska folket skyddas genom tillfällig internationell närvaro på de ockuperade områdena i överensstämmelse med säkerhetsrådets resolution 904 (1994).
På begäran av parterna skall Europeiska unionen genomföra ett samordnat program för bistånd till förberedelse och övervakning av de val på de ockuperade områdena som påbjöds i principdeklarationen av den 13 september 1993. De exakta praktiska arrangemangen och finansieringen skall fastställas i ett särskilt rådsbeslut när Israel och PLO har enats om hur valet skall arrangeras. Europaparlamentet kommer att inbjudas att delta i dessa arrangemang.
Artikel 7
Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
För att säkerställa att kontrollerna på bestämmelseorten utförs effektivt, och för att förhindra att det senare uppstår svårigheter i handeln inom gemenskapen, bör det, samtidigt som de berörda parternas intressen skyddas, fastställas vissa närmare bestämmelser om provtagningen.
Artikel 1
RÅDETS BESLUT av den 24 oktober 1994 om utsträckning av det rättsliga skyddet för kretsmönster i halvledarprodukter till personer från Canada (94/700/EG)
med beaktande av rådets direktiv 87/54/EEG av den 16 december 1986 om rättsligt skydd för kretsmönster i halvledarprodukter(1), särskilt artikel 3.7 i detta,
Rätten till skydd kan genom ett rådsbeslut utsträckas till personer som inte åtnjuter skydd genom de nämnda bestämmelserna.
Canada har bestämmelser som ger lämpligt skydd till kretsmönsterskapare och landet har tillkännagett att man planerar att uträcka tillämpningen av dessa bestämmelser från och med den 1 november 1994 till att omfatta gemenskapsmedborgare och fysiska och juridiska personer som bedriver verklig och stadigvarande verksamhet i gemenskapen i syfte att skapa kretsmönster eller tillverka integrerade kretsar.
Med tanke på de kanadensiska myndigheternas åtaganden bör rätten till skydd enligt direktiv 87/54/EEG utsträckas, från och med den 1 november 1994 till dess bestämmelserna i avtalet om handelsrelaterade aspekter på immateriella rättigheter har genomförts, till att omfatta fysiska personer, bolag och andra juridiska personer från Canada.
Medlemsstaterna skall utsträcka det skydd som avses i direktiv 87/54/EEG enligt följande:
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Enligt turkisk lagstiftning ansvarar Ministry of Agriculture and Rural Affairs för hälsokontrollen av levande tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar samt för övervakningen av de hygieniska och sanitära förhållandena vid produktionen. Enligt samma lagstiftning är Ministry of Agriculture and Rural Affairs bemyndigad att tillåta eller förbjuda upptagning av tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar i vissa områden.
De behöriga myndigheterna i Turkiet har officiellt garanterat att de krav som anges i kapitel V i bilagan till direktiv 91/492/EEG och att krav som motsvarar de som föreskrivs i det direktivet vad avser klassificering av upptagnings- och återutläggningsområden, godkännande av leveransanläggningar, hygienkontroll och övervakning av produktionen uppfylls. Kommissionen skall framför allt underrättas om alla eventuella ändringar av upptagningsområdena.
De särskilda importvillkoren påverkar inte tillämpningen av de beslut som fattas enligt rådets direktiv 91/67/EEG av den 28 januari 1991 om djurhälsovillkor för utsläppande på marknaden av djur och produkter från vattenbruk(2).
3. De skall vara förpackade i förseglade förpackningar av en godkänd leveransanläggning som är upptagen i förteckningen i bilaga C.
- Art (gängse och vetenskapligt namn).
Artikel 3
Artikel 4
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Bestämmelserna om kontrollmärkning av produkter från sådana förpackningsanläggningar bör fastställas.
Artikel 1
Artikel 2
Om produkter från olika produktionsföretag plockas samman skall förpackningsanläggningens kontrollmärke åsättas det yttersta emballaget som produkterna paketeras i på förpackningsanläggningen.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 64/433/EEG av den 26 juni 1964 om hälsoproblem som påverkar handeln med färskt kött inom gemenskapen(3), ändrat genom del 1 kapitel 3 punkt 1. d i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 5.4 i detta,
Den 10 oktober och den 13 december 1994 förelade Finland kommissionen sitt operativa program för bekämpning av salmonella i enlighet med artikel 10a.2 i direktiv 64/432/EEG, artiklarna 9a, 9b och 10b i direktiv 90/539/EEG, artikel 5 i direktiv 64/433/EEG, artikel 5 i direktiv 71/118/EEG och första strecksatsen i kapitel 2 i bilaga 2 till direktiv 92/118/EEG.
De salmonellagarantier som gäller för Finland, redan fastställda eller som kommer att fastställas i framtiden, skall specificeras för varje kategori av levande djur och animaliska produkter. Tillämpningen av nämnda garantier är beroende av att de åtgärder som Finland skall vidta inom varje sektor godkänns.
Det finska programmets åtgärder avseende nötkreatur och svin för avel, produktion och slakt godkänns.
Artikel 3
Det finska programmets åtgärder avseende slaktfjäderfä godkänns.
Artikel 6
Det finska programmets åtgärder avseende ägg för direkt konsumtion som livsmedel godkänns.
Artikel 9
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av följande: Enligt rådets förordning (EEG) nr 386/90 av den 12 februari 1990 om kontroll i samband med export av jordbruksprodukter som berättigar till exportbidrag eller andra belopp(3), måste kommissionen för rådet framlägga en rapport om framstegen i tillämpningen av förordningen.
Generellt sett bör kontrollsatsen ligga kvar på 5 %, men ordningen kan göras smidigare, så att kontrollorganen kan koncentrera sina insatser på känsligare produkter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- per tullkontor,
Procentsatsen på 5 % per produktsektor kan dock ersättas med en procentsats på 5 % för samtliga sektorer, förutsatt att medlemsstaten tillämpar ett urvalssystem baserat på riskanalys vilken utförs enligt kriterier som närmare skall fastställas i enlighet med det förfarande som anges i artikel 6. I så fall är en lägsta procentsats på 2 % per produktsektor obligatorisk."
KOMMISSIONENS FÖRORDNING (EG) nr 1966/94 av den 28 juli 1994 om klassificering av vissa varor i Kombinerade nomenklaturen
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom kommissionens förordning (EG) nr 1737/94(2), särskilt artikel 9 i denna, och med beaktande av följande:
Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
Beträffande produkterna nr 1, 2 och 4 i bifogade tabell är de åtgärder som föreskrivs i denna förordning förenliga med yttrandet från Tullkodexkommitténs sektion för tulltaxe- och statistiknomenklatur.
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Sedan förordningen antogs har bilagorna ändrats ett antal gånger. På grund av ändringarnas antal, komplexitet och det faktum att de är spridda i olika nummer av Europeiska gemenskapernas officiella tidning är texterna svåra att använda och saknar den klarhet som bör vara utmärkande för all lagstiftning. De bör därför kodifieras. Samtidigt bör namnen på eller de kemiska beteckningarna för vissa föreningar rättas till eller preciseras och några sakfel korrigeras.
Artikel 1
Denna förordning träder i kraft den sextionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Enligt artikel 2.3 i anslutningsfördraget(4) kan Europeiska unionens institutioner före anslutningen fatta de beslut som avses i artikel 169 i anslutningsakten, varvid dessa beslut träder i kraft om och när detta fördrag träder i kraft.
Förordning (EEG) nr 2273/93 skall ändras på följande sätt: De interventionsorter med tillhörande upplysningar som anges i bilagan till denna förordning skall läggas till i bilagan till förordning (EEG) nr 2273/93.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De rättsliga bestämmelser som gäller i Marocko för hälsobesiktning och -kontroll av fiskeriprodukter kan anses vara likvärdiga med dem som fastställs i direktiv 91/493/EEG.
I enlighet med artikel 11.4 b i direktiv 91/493/EEG är det viktigt att på fiskeriprodukternas förpackningar fästa ett märke som anger namnet på det tredje land som avses och ursprungsanläggningens godkännandenummer.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
2. Intyget bör vara försett med DEMA-ombudets namn, dennes tjänsteställning och underskrift samt med DEMA:s officiella stämpel och allt bör vara i en färg som avviker från de övriga uppgifter som finns på intyget.
Artikel 5
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 2.1 skall ersättas med följande:
KOMMISSIONENS FÖRORDNING (EG) nr 1442/95 av den 26 juni 1995 med ändring av bilagorna I, II, III och IV i rådets förordning (EEG) nr 2377/90 som upprättar ett gemenskapsförfarande för fastställande av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (Text av betydelse för EES)
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 som upprättar ett gemenskapsförfarande för fastställande av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (1), vilket tidigare omformulerats genom kommissionens förordning (EEG) nr 1441/95 (2), särskilt artikel 6, 7 och 8 i denna, och
Det vid fastställandet av gränsvärden för högsta tillåtna restmängder vad gäller restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung är det nödvändigt att klargöra i vilken djurart restmängder förefinnes, såväl den befintliga mängden i samtliga berörda köttvävnader härrörande från det behandlade djuret (målvävnad), som vilken sorts restmängd, vilket är av betydelse vid kontrollen av restmängder (restmängd markör).
Carazolol, diazinon och spiramycin (gäller nöt och kyckling) skulle tillföras bilaga I till förordning (EEG) nr 2377/90.
För att möjliggöra komplettering av vetenskapliga studier, bör giltighetstiden för temporär MRL, tidigare definierad i bilaga III i förordning (EEG) nr 2377/90, förlängas för tylosin och spiramycin (gäller svin).
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för anpassning till tekniska framsteg av direktiven för avskaffande av tekniska handelshinder inom sektorn veterinärmedicinska läkemedel.
Bilaga I, II, III och IV i förordning (EEG) nr 2377/90 skall ändras enligt denna förordning.
KOMMISSIONENS FÖRORDNING (EG) nr 1662/95 av den 7 juli 1995 om fastställande av vissa närmare föreskrifter för genomförandet av gemenskapens beslutförande för att godkänna utsläppandet på marknaden av humanläkemedel och veterinärmedicinska läkemedel
med beaktande av rådets förordning (EEG) nr 2309/93 av den 22 juli 1993 om gemenskapsförfaranden för godkännande för försäljning av och tillsyn över humanläkemedel och veterinärmedicinska läkemedel samt om inrättande av en europeisk läkemedelsmyndighet (1), särskilt artiklarna 10.3 och 32.3 i denna och, med beaktande av följande:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 3
Artikel 4
Artikel 5
Om förslaget till beslut skall behandlas vid ett sammanträde med kommittén skall kallelsen, dagordningen och, i fall enligt artikel 2 andra stycket, det förslag till beslut över vilket kommitténs yttrande begärs, av ordföranden överlämnas till medlemmarna i kommittén i enlighet med bestämmelserna i artikel 7.
Korrespondens till medlemmarna i kommittén skall, då kommittén sammanträder enligt det förfarande som avses i artikel 1, sändas genom skriftlig telekommunikation till de behöriga nationella organ som varje medlemsstat utsett för detta ändamål. En kopia skall sändas till den berörda medlemsstatens ständiga representation.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande, och
Det är väsentligt att den enhetliga modellen för visumhandlingar innehåller alla nödvändiga uppgifter och svarar mot mycket högt ställda tekniska krav, bl.a i fråga om garantier mot efterbildningar och förfalskningar. Den enhetliga modellen måste även vara utformad så att den kan användas i samtliga medlemsstater och innefatta säkerhetsanordningar som är allmänt igenkännliga och kan uppfattas med blotta ögat.
För att uppnå sitt syfte skall denna förordning vara tillämplig på alla typer av visumhandlingar enligt artikel 5. Medlemsstaterna bör ha möjligheten att använda samma modell för att utfärda visumhandlingar för andra ändamål än de som anges i artikel 5, förutsatt att dessa, på grund av ändringar som kan uppfattas med blotta ögat, inte kan förväxlas med den enhetliga visumhandlingen.
Artikel 1
Kompletterande tekniska specifikationer för att förhindra efterbildningar eller förfalskningar av visumhandlingen skall fastställas i enlighet med förfarandet i artikel 6.
2. Varje medlemsstat skall utse endast ett organ som ansvarar för tryckningen av visumhandlingar. Namnet på detta organ meddelas till kommissionen och till de övriga medlemsstaterna. Två eller flera medlemsstater får utse samma organ för detta ändamål. Varje medlemsstat får byta detta organ. I så fall skall kommissionen och de andra medlemsstaterna underrättas.
2. Modellen för visumhandlingen innehåller inga andra maskinellt läsbara upplysningar än de som också finns i de rutor som beskrivs i punkterna 6 till 12 i bilagan eller på motsvarande resehandling.
- en vistelse i denna medlemsstat eller i flera medlemsstater för en period som totalt inte överstiger tre månader,
1. När hänvisning sker till förfarandet enligt denna artikel, gäller följande bestämmelser:
3. a) Kommissionen skall anta förslaget om åtgärder om det är förenligt med kommitténs yttrande.
Artikel 7
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
Den av rådet begärda förnyade granskningen av artiklarna 5, 10 och 11 inför den 1 juli 1994 har visat nödvändigheten av att göra vissa tekniska och redaktionella ändringar i dessa artiklar samt i vissa andra bestämmelser för att kunna garantera en effektiv administrering och tillämpning av förordningen. Utarbetandet av dessa förändrade regler har följaktligen prioriterats och utformningen av regler för animalisk produktion måste därför skjutas upp under en begränsad tid.
Det har dessutom framkommit, att förökningsmaterial bör härröra från ekologiskt odlade växter men att undantagsbestämmelser är nödvändiga för att under en övergångsperiod ge odlarna möjlighet att använda förökningsmaterial som erhållits på konventionellt sätt i fall då det inte finns tillgång till lämpligt material som erhållits enligt ekologiska odlingsmetoder.
Artikel 1
2. Artikel 4.2 ersätts med följande text:
"3. `beredning`: åtgärder för konservering och/eller bearbetning av jordbruksprodukter samt förpackning och/eller ändringar av presentationen av det ekologiska produktionsförfarandet som används vid märkningen av de färska konserverade och/eller bearbetade produkterna."
5. Följande punkter läggs till i artikel 4:
6. I artikel 2, artikel 5.1 b, artikel 9.9 a, artikel 11.1 b, artikel 11.2 a och artikel 11.6 a ersätts orden "artikel 6 och 7" med orden "artikel 6".
8. Artikel 5.2 utgår.
a) minst 95 % av produktens ingredienser av jordbruksursprung är produkter eller är framställda ur produkter som har erhållits i enlighet med de regler som fastställs i artikel 6 eller som har importerats från tredje land inom ramen för den ordning som anges i artikel 11,
d) produkten eller dess ingredienser av jordbruksursprung som anges i punkt a har inte behandlats med andra ämnen än de som anges i bilaga VI punkt b,
g) för produkter som beretts efter den 1 januari 1997 skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som den leverantör som har utfört den sista beredningsåtgärden är underställd. Valet av om namn eller kodnummer skall användas åligger medlemsstaten som skall meddela sitt beslut till kommissionen.
"4. Ingredienser av jordbruksursprung får ej förekomma i bilaga VI punkt C annat än när det visas att dessa ingredienser är av jordbruksursprung, att de inte produceras i tillräcklig mängd inom gemenskapen enligt reglerna i artikel 6 eller att de inte kan importeras från tredje land enligt reglerna i artikel 11."
a) de krav som anges i punkt 1 respektive 3 är helt uppfyllda utom vad gäller längden på den övergångsperiod som avses i punkt 1 i bilaga I,
d) produkten innehåller en enda ingrediens av jordbruksursprung,
"5a. Utan det påverkar tillämpningen av punkt 3 får sådan märkning av och reklam för en produkt som anges i artikel 1.1 b inte vara försedd med uppgifter som hänvisar till den ekologiska produktionsmetoden annat än om följande villkor är uppfyllda:
c) uppgifter som hänvisar till ekologisk produktion nämns i ingrediensförteckningen och hänför sig uppenbarligen endast till de ingredienser som erhållits i enlighet med reglerna i artikel 6 eller som importerats från tredje land inom ramen för den ordning som anges i artikel 11. De skall presenteras i en färg, ett format och en typstil som helt överensstämmer med vad som används för övriga uppgifter som finns på ingrediensförteckningen. Dessa uppgifter skall också nämnas separat inom samma synfält som beskrivningen av den saluförda varan och skall innehålla upplysning om den procentuella andel av ingredienserna som är av jordbruksursprung eller som härrör från ingredienser som är av jordbruksursprung och som har erhållits i enlighet med reglerna i artikel 6 eller som importerats från tredje land inom ramen för den ordning som anges i artikel 11. Det nämnda får inte göras i en färg, ett format eller en typstil som gör den mer framträdande än beskrivningen av den saluförda varan. Omnämnandet skall ges följande utformning: `X % av ingredienserna av jordbruksursprung har erhållits i enlighet med reglerna för ekologisk produktion`,
f) produkten eller dess ingredienser har inte behandlats med joniserande strålning,
13. Artikel 5.6 ersätts med följande:
b) produkten uppfyller kraven i punkt 3 c, d, e och f,
- hänför sig uppenbarligen endast till de ingredienser som erhållits i enlighet med de regler som avses i artikel 6, eller som har importerats inom ramen för den ordning som anges i artikel 11,
14. Inledningen till 5.8 ersätts med följande text:
"9. Beräkningen av de i punkterna 3 och 6 angivna procentandelarna utförs med tillämpning av reglerna i artiklarna 6 och 7 i direktiv 79/112/EEG.
16. Artikel 6 ersätts med följande text:
a) åtminstone de bestämmelser som anges i bilaga I och, i förekommande fall, de tillämpningsförfaranden som hör till dessa skall vara uppfyllda,
2. För utsäde och vegetativt förökningsmaterial innebär den ekologiska produktionsmetoden att både moderplantan - såvitt avser utsäde - och föräldragenerationens planta/plantor - såvitt avser reproduktionsmaterial - har producerats i överensstämmelse med bestämmelserna i punkt 1 a och b under minst en generation eller, när det gäller perenna odlingar, minst två säsonger.
- införande, före den 31 december 2000, av begränsningar gällande den provisoriska åtgärd som anges i a i fråga om vissa arter och/eller typer av förökningsmaterial och/eller avsaknad av kemisk behandling,
4. Före den 31 december 1999, skall kommissionen göra en förnyad granskning av bestämmelserna i denna artikel, särskilt punkt 1 c samt punkt 2 och i förekommande fall presentera lämpliga förslag till ändring av dem."
1. I denna artikel anses med `plantor` hela plantor, avsedda för plantering för produktion av växter.
a) medlemsstatens behöriga myndighet har godkänt användning under förutsättning att användaren eller användarna av sådant material på ett tillfredsställande sätt kunnat visa medlemsstatens kontrollmyndighet eller kontrollorgan att de inte kunnat erhålla lämplig sort av ifrågavarande art på gemenskapsmarknaden,
d) efter plantering skall plantorna ha odlats i enlighet med bestämmelserna i artikel 6.1 a och b under en period av minst sex veckor före skörden,
4. a) När godkännanden som avses i punkt 3 har lämnats skall medlemsstaten omedelbart lämna följande upplysningar till övriga medlemsstater och kommissionen:
- nödvändiga mängder samt skälen för detta,
4. b) Om upplysningar, som av en medlemsstat lämnats till kommissionen och den medlemsstat som har lämnat godkännande, visar att en lämplig sort finns tillgänglig under den tid brist råder, får medlemsstaten återkalla ett godkännande eller förkorta dess giltighetstid. Medlemsstaten skall i sådant fall meddela kommissionen och de andra medlemsstaterna om de åtgärder den vidtagit senast inom tio dagar efter det att den mottagit upplysningarna.
"1a. De villkor som anges i punkt 1 gäller inte för produkter, som före antagandet av denna förordning allmänt användes i enlighet med vedertagna regler för ekologisk odling inom gemenskapen".
21. I artikel 9.6 c ersätts ordet "överträdelser" med orden "avvikelser och/eller överträdelser".
"6a. Medlemsstaterna skall före den 1 januari 1996 tilldela varje kontrollorgan eller kontrollmyndighet som godkänts eller utsetts i enlighet med bestämmelserna i denna förordning ett kodnummer. De skall meddela övriga medlemsstater och kommissionen om detta och kommissionen skall offentliggöra kodnummer i den förteckning som anges i sista stycket i artikel 15."
25. Artikel 10.1 ersätts med följande text:
b) har varit underkastad den kontroll som avses i artikel 9 under hela produktions- och beredningsprocessen,
26. I artikel 10.3 a ersätts orden "artikel 5-7" med orden "artiklarna 5 och 6".
Artikel 10a
28. I artikel 11.3 a ersätts orden "kontrollmyndigheterna" med orden "kontrollorgan och/eller kontrollmyndighet".
"Den upphör från och med den tidpunkt då beslut att föra in ett tredje land i förteckningen som anges i punkt 1 a fattas, förutsatt att den inte rör en produkt som härrör från ett område som inte närmare preciseras i det beslut som anges i punkt 1 a och att den inte har granskats inom ramen för det tredje landets ansökan. Det tredje landet skall vara införstått med den fortsatta tillämpningsregeln av det förfarande för godkännande som anges i denna punkt."
32. I artikel 13 införs följande strecksats före första strecksatsen:
"- de ändringar som skall göras i bilaga V för att fastlägga en logotyp för gemenskapen som kan användas tillsammans med eller i stället för uppgiften om att produkterna omfattas av ett särskilt kontrollsystem."
KOMMISSIONENS FÖRORDNING (EG) nr 2694/95 av den 21 november 1995 om klassificering av vissa varor i Kombinerade nomenklaturen
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 2588/95 (2), särskilt artikel 9 i denna, och med beaktande av följande:
Artikel 1
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
KOMMISSIONENS FÖRORDNING (EG) nr 2802/95 av den 4 december 1995 om klassificering av vissa varor i Kombinerade nomenklaturen
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 2588/95 (2), särskilt artikel 9 i denna, och med beaktande av följande:
Artikel 1
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
KOMMISSIONENS FÖRORDNING (EG) nr 2805/95 av den 5 december 1995 om fastställande av exportbidrag inom vinsektorn och upphävande av förordning (EEG) nr 2137/93
med beaktande av rådets förordning (EEG) nr 822/87 av den 16 mars 1987 om den gemensamma organisationen av marknaden för vin (1), senast ändrad genom förordning (EG) nr 1544/95 (2), särskilt artikel 55.8 i denna, och
Artikel 1
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EEG) nr 2771/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för ägg (3), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94 (4), särskilt artiklarna 3.2, 5.4, 6.4 och 18.13 i denna,
med beaktande av rådets förordning (EEG) nr 715/90 av den 5 mars 1990 om de bestämmelser som gäller för jordbruksprodukter och vissa varor som framställts genom förädling av jordbruksprodukter som har sitt ursprung i AVS-staterna eller i de utomeuropeiska länderna och territorierna (ULT) (7), senast ändrad genom förordning (EG) nr 2484/94 (8), särskilt artikel 27.2 i denna,
med beaktande av rådets förordning (EG) nr 3296/94 av den 19 december 1994 om vissa förfaranden för tillämpning av Europaavtalet om associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Tjeckien, å andra sidan (12), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 774/94 av den 29 mars 1994 om öppnande och förvaltning av vissa gemenskapstullkvoter för nötkött av hög kvalitet, griskött, fjäderfäkött, vete och blandsäd av vete och råg samt kli och andra restprodukter (16), senast ändrad genom kommissionens förordning (EG) nr 2198/95 (17), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 1275/95 av den 29 maj 1995 om vissa förfaranden för tillämpningen av avtalet om frihandel och vissa handelsrelaterade frågor mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Estland, å andra sidan (20), särskilt artikel 1 i denna,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- i artikel 1.1 i förordning (EEG) nr 2777/75,
3. KN-nummer 1602 32 skall införas före KN-nummer 1602 39
4. KN-nummer 0207 23 skall ersättas med KN-nummer 0207 33 i bilaga I till kommissionens förordning (EEG) nr 1729/92 (27).
- kommissionens förordning (EG) nr 1559/94 (30),
- kommissionens förordning (EG) nr 1866/95 (33).
>Plats för tabell>
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
Internationella säkerhetsorganisationskoden för säker drift av fartyg och för förhindrande av förorening (hädanefter kallad "ISM-koden") antogs av Internationella sjöfartsorganisationen (IMO) genom församlingens resolution A.741(18) av den 4 november 1993 i medlemsstaternas närvaro och kommer, genom att den införlivas med 1974 års internationella konvention om säkerheten för människoliv till sjöss, att från och med den 1 juli 1998 tillämpas på ro-ro-passagerarfartyg.
Den mest brådskande angelägenheten för gemenskapen utgörs av säkerhetsorganisationen på ro-ro-passagerarfartyg. Ett enhetligt och sammanhängande genomförande av ISM-koden i alla medlemsstater kan utgöra ett steg i riktning mot en säkerhetsorganisation för ro-ro-passagerarfartyg.
Åtgärder på gemenskapsnivå är det bästa sättet att säkerställa ett påskyndat, tvingande genomförande av bestämmelserna i ISM-koden och en effektiv kontroll av tillämpningen av denna, samtidigt som en snedvridning av konkurrensen mellan olika gemenskapshamnar och ro-ro-passagerarfartyg undviks. Endast en förordning som är direkt tillämplig kan säkerställa ett sådant genomförande. För ett påskyndat genomförande krävs att förordningen tillämpas från och med den 1 juli 1996.
Företag som endast bedriver trafik med ro-ro-passagerarfartyg i skyddade vatten mellan hamnar i samma medlemsstat utgör en mera begränsad risk och kommer att behöva utföra en proportionellt sett större mängd administrativt arbete än andra företag och bör därför beviljas ett temporärt undantag.
En medlemsstat måste under förutsättning av att ett för medlemsstaterna bindande beslut fattas inom ramen för en föreskrivande kommitté ha rätt att tillfälligt dra in rätten att bedriva trafik med vissa ro-ro-passagerarfartyg från dess hamnar när den anser att det föreligger risk för allvarlig fara för säkerheten för liv eller egendom eller för miljön.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- att företagen inrättar och på lämpligt vis upprätthåller ombordbaserade och landbaserade säkerhetsorganisationssystem, och
I denna förordning och för genomförandet av ISM-koden avses med
1. enligt en offentliggjord tidtabell, eller
d) erkänd organisation: ett organ som erkänts i enlighet med bestämmelserna i direktiv 94/57/EG.
g) dokument om godkänd säkerhetsorganisation: det dokument som i enlighet med punkt 13.2 i ISM-koden utfärdas till företag,
Artikel 3
1. Alla företag skall följa samtliga bestämmelser i punkterna 1.2 13.1 och 13.3 i ISM-koden, som om dessa bestämmelser vore tvingande, som ett villkor för att deras fartyg skall få bedriva reguljär trafik till eller från en hamn i en medlemsstat inom den Europeiska gemenskapen.
1. Medlemsstaterna skall, med avseende på företag och ro-ro-passagerarfartyg, följa bestämmelserna i punkterna 13.2, 13.4 och 13.5 i ISM-koden som om dessa bestämmelser vore tvingande.
3. Dokumentet om godkänd säkerhetsorganisation skall endast gälla i fem år från dagen för dess utfärdande, under förutsättning att en kontroll görs en gång om året, för att bekräfta att säkerhetsorganisationssystemet fungerar väl, och att eventuella ändringar som gjorts sedan den senaste kontrollen uppfyller ISM-kodens bestämmelser.
6. En medlemsstat skall erkänna dokument om godkänd säkerhetsorganisation och certifikat om godkänd säkerhetsorganisation som utfärdats av administrationerna i tredje land, eller för dessas räkning, om det kan visas att de följer bestämmelserna i denna förordning.
Medlemsstaterna skall förvissa sig om att bestämmelserna i denna förordning följs av alla företag som bedriver reguljär färjetrafik med ro-ro-passagerarfartyg till eller från deras hamnar.
Under ovannämnda förhållanden skall följande förfarande tillämpas:
Artikel 9
b) Giltighetstiden för dokumentet om godkänd säkerhetsorganisation och/eller certifikatet om godkänd säkerhetsorganisation och intervallen mellan kontrollerna av dem i artikel 5.3 och 5.4.
1. Kommissionen skall biträdas av den kommitté som inrättas enligt artikel 12.1 i rådets direktiv 93/75/EEG (7).
b) Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Utan att det påverkar första stycket skall denna förordning inte tillämpas före den 31 december 1997 på företag som lyder under grekisk lag, har sin huvudsakliga verksamhetsort i Grekland och bedriver färjetrafik med ro-ro-passagerarfartyg som är registrerade i Grekland, för grekisk flagg och bedriver reguljär trafik endast mellan hamnar som är belägna i Grekland.
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Europaparlamentets yttrande (2),
Genom denna övervakningsverksamhet har de viktigaste aspekterna på de förändringar av gemenskapens jordbruksstatistik som krävs fastställts.
a) uppgifterna fortsätter att vara tillräckligt tillförlitliga för varje medlemsstat och jämförbara medlemsstaterna emellan,
d) planeringen av nationella åtgärder tar tillbörlig hänsyn till det kollektiva gemenskapsintresset,
Ett finansiellt bidrag till medlemsstaterna, i förhållande till deras objektiva behov, krävs för att underlätta nödvändiga anpassningar.
Fördelningen av uppgifter mellan kommissionen och medlemsstaterna är helt i överensstämmelse med subsidiaritetsprincipen.
Syfte
Kommissionens uppgift
b) kontrollera uppgifternas kvalitet och jämförbarhet, samt
Tidsplan och förfarande
Tekniska handlingsplaner för jordbruksstatistiken
a) Befintliga åtaganden för åren i fråga, t.ex. en förteckning över de gemenskapsundersökningar som medlemsstaterna skall genomföra och frekvensen av dessa, samt andra uppgifter som skall lämnas till kommissionen.
Artikel 5
a) en kort rapport om genomförandet av de åtgärder som beslutades för det föregående året (år ng 1),
Beskrivningen skall omfatta de ändringar som anges avseende metodologin för genomförandet, arbeten som skall utföras, förutsedda svårigheter och förslag till lösningar på dem, konsekvenser för nationella och gemensamma resurser samt förslag till förbättringar på gemenskapsnivå. De åtgärder för vilka ekonomiskt gemenskapsstöd kommer att begäras skall anges.
Finansiella bestämmelser
3. Bidraget skall ges till medlemsstaterna årsvis efter det att de överlämnat den årliga rapporten om genomförandet av planerade åtgärder under det föregående året och den blivit godkänd av kommissionen. Kommissionen kan i samarbete med behöriga myndigheter i medlemsstaterna utföra alla kontrollåtgärder på plats som den anser nödvändiga.
Då det med hänsyn till syftet med detta beslut är nödvändigt, kan kommissionen för en period som motsvarar en teknisk handlingsplan, i enlighet med förfarandet i artikel 10, godkänna en medlemsstats begäran om att anpassa en eller flera av följande undersökningskarakteristika i bilaga IV: undersökta regioner, territoriella underindelningar, definitioner, undersökningsmetodik, undersökningstidpunkt, variabellista och klassernas storlek.
Kommissionen kan göra ändringar i bilaga I (statistiska områden där möjliga besparingar har fastställts) och i bilaga II (statistiska områden där det finns nya eller växande behov) i enlighet med förfarandet i artikel 10. Den skall informera Europaparlamentet och rådet om de ändringar som gjorts.
Ständiga kommittén för jordbruksstatistik, som inrättades genom rådets beslut 77/279/EEG (5) skall sammanträda minst en gång om året för att diskutera följande:
c) Den tekniska handlingsplanen för det kommande året.
Artikel 10
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittéen skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen, varvid medlemsstaternas röster skall vägas enligt samma artikel. Ordföranden får inte rösta.
Om rådet inte har beslutat inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Senast den 1 november 1997 och efter samråd med Ständiga kommittén för jordbruksstatistik skall kommissionen till Europaparlamentet och rådet överlämna en rapport om genomförandet av detta beslut, vid behov åtföljd av förslag till dess förlängning.
KOMMISSIONENS BESLUT av den 20 maj 1996 om utsläppande på marknaden av en genetiskt modifierad hansteril cikoria med partiell tolerans mot herbiciden glufosinatammonium (Cichorium intybus L.) enligt rådets direktiv 90/220/EEG (Text av betydelse för EES) (96/424/EG)
med beaktande av rådets direktiv 90/220/EEG av den 23 april 1990 om avsiktlig utsättning av genetiskt modifierade organismer i miljön (1), ändrat genom kommissionens direktiv 94/15/EG (2), särskilt artikel 13 i detta, och med beaktande av följande:
Nederländernas behöriga myndighet har överlämnat handlingarna i ärendet till kommissionen med tillstyrkan. De behöriga myndigheterna i andra medlemsstater har rest invändningar mot handlingarna.
- Det finns ingen anledning att tro att det skulle uppstå negativa inverkningar genom en överföring av bar-genen till vilda cikoriapopulationer; eftersom en sådan överföring endast skulle utgöra en konkurrensmässig eller selektiv fördel gentemot vilda populationer om herbiciden glufosinatammonium vore den enda faktorn som begränsade dessa populationer, vilket inte är fallet.
- Eftersom 50 % av det hybrida utsädet är tolerant mot herbiciden i fråga, bör etiketten ange att produkten kan vara tolerant mot herbiciden glufosinatammonium, så att odlarna är medvetna om att det eventuellt inte är möjligt att kontrollera oönskade groddar av produkter med glufosinatammonium.
Detta beslut är förenligt med yttrandet från den kommitté bestående av företrädare för medlemsstaterna som inrättas enligt artikel 21 i direktiv 90/220/EEG.
1. Utan att det påverkar gemenskapslagstiftningen, och i överensstämmelse med de villkor som fastställs i styckena 2, 3 och 4, skall tillstånd för utsläppande på marknaden ges av de nederländska myndigheterna för följande produkt anmäld av Bejo-Zaden BV (ref. C/NL/94/25) i enlighet med artikel 13 i direktiv 90/220/EEG.
ii) Bar-genen från Streptomyces hygroscopicus (fosfinotricinacetyltransferas) med promotorn PSsuAra-tp från Arabidopsis thaliana och TL-DNA-gen-7-promotorn från Agrobacterium tumefaciens.
3. Medgivandet avser användning av produkten för odlingsverksamhet.
- och kan vara tolerant mot herbiciden glufosinatammonium.
KOMMISSIONENS BESLUT av den 28 juni 1996 om särskilda importvillkor för fiskeri- och vattenbruksprodukter med ursprung i Mauretanien (Text av betydelse för EES) (96/425/EG)
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av fiskeriprodukter (1), senast ändrat genom direktiv 95/71/EG (2) uppfylls, särskilt artikel 11 i detta, och med beaktande av följande:
"Ministère des Pêches et de l'Économie Maritime - Centre National de Recherches Océanographiques et des Pêches - Département Valorisation et Inspection Sanitaire (MPEM - CNROP - DVIS)" kan på ett effektivt sätt granska tillämpningen av den gällande lagstiftningen.
I enlighet med artikel 11.4 c i direktiv 91/493/EEG är det viktigt att fastställa en förteckning över godkända anläggningar eller frysfartyg. Denna förteckning bör fastställas på grundval av ett meddelande från MPEM - CNROP - DVIS till kommissionen. Det åligger alltså MPEM - CNROP - DVIS att försäkra sig om att de åtgärder som föreskrivs i detta syfte i artikel 11.4 i direktiv 91/493/EEG efterlevs.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 4
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
En expertdelegation utsänd av kommissionen har kommit tillbaka från Elfenbenskusten efter att ha förvissat sig om villkoren för produktion, lagring och transport av fiskeriprodukter med gemenskapen som destination.
Villkoren för det intyg som avses i artikel 11.4 a i direktiv 91/493/EEG omfattar fastställande av en mall för intyget, vilket eller vilka språk intyget skall vara avfattat på och vilken ställning den som undertecknar intyget skall ha.
MARA-DGRA har officiellt gett försäkringar i fråga om efterlevnaden av de regler som anges i kapitel V i bilagan till direktiv 91/493/EEG och i fråga om krav som är likvärdiga med dem som föreskrivs i det direktivet för godkännande av anläggningar.
1. Det intyg som avses i artikel 2.1 skall utfärdas på minst ett av de officiella språken i den medlemsstat där kontrollen äger rum.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande Ekonomiska och sociala kommitténs yttrande (3), och
3. Vissa substanser med tyreostatisk, östrogen, androgen eller gestagen verkan kan, p.g.a. de restsubstanser de ger i kött och andra livsmedel av animaliskt ursprung, vara farliga för konsumenterna och de kan även påverka kvalitén i livsmedel av animaliskt ursprung.
6. Olämplig användning av â-agonister kan innebära allvarlig fara för människors hälsa. För konsumenternas skull bör innehav av â-agonister liksom tillförsel till alla slags djur samt avyttring för detta syfte förbjudas. Innehav av stilbener och tyreostatiska medel liksom tillförsel till alla slags djur och avyttring bör också förbjudas. Användningen av andra ämnen bör regleras.
9. Det är lämpligt att behålla förbudet mot hormonella ämnen i tillväxtbefrämjande syfte. Om tillförsel av vissa ämnen kan tillåtas i terapeutiskt eller zootekniskt syfte skall den noggrant kontrolleras för att undvika varje form av felaktig användning.
12. Undantag kan tillåtas om tillräckliga garantier ges för att förebygga obalans i handeln. Dessa garantier bör gälla produkter som kan användas, villkor för deras användning och kontroll av dessa villkor, särskilt när det gäller att respektera den nödvändiga karenstiden.
15. För att illegal användning av tillväxtbefrämjande och produktivitetshöjande medel i animalieproduktion skall kunna bekämpas effektivt i alla medlemsstater bör de åtgärder som skall vidtas organiseras på gemenskapsnivå.
Artikel 1
a) husdjur: tama djur av arterna nötkreatur, svin, får getter, hovdjur, fjäderfä och kaniner, samt vilda djur av dessa arter och vilda idisslare, uppfödda i hägn,
i) tillförsel till enstaka husdjur av ett av de ämnen som tillåts enligt artikel 5 i detta direktiv, i syfte att synkronisera östrus och förbereda donatorer och recipienter vid implantation av embryon, efter det att djuret undersökts av veterinär eller enligt artikel 5, stycke 2, på dennes ansvar,
Artikel 3
b) Innehav av djur som avses i a i ett jordbruksföretag, utom under officiell kontroll samt avyttring eller slakt, som livsmedel, av husdjur eller vattenbruksdjur som innehåller ämnen som avses i a eller i vilka förekomsten av sådana ämnen har konstaterats, utom i det fall det kan bevisas att dessa djur har behandlats enligt artikel 4 eller 5.
e) Bearbetning av kött som avses i d.
1. Tillförsel till husdjur i terapeutiskt syfte av östradiol 17 â, testosteron, progesteron eller derivat som efter resorption på platsen för applicering vid hydrolys bildar den ursprungliga komponenten. Veterinärmedicinska läkemedel som används för terapeutisk behandling skall uppfylla föreskrifterna för avyttring enligt direktiv 81/851/EEG och kan tillföras endast av veterinär på husdjur som noggrant identifierats och i form av injektion eller för behandling av äggstocksrubbningar i form av vaginalspiral, men inte i form av implantat. Behandling av identifierade djur skall registreras av den ansvarige veterinären. Denne skall i ett register, som kan vara det som föreskrivs i direktiv 81/851/EEG, anteckna minst följande upplysningar:
- behandlingsdatum,
2. Tillförsel i terapeutiskt syfte av registrerat veterinärmedicinskt läkemedel som innehåller
Tillförseln skall utföras av veterinär eller, vad beträffar veterinärmedicinska läkemedel enligt i, på dennes direkta ansvar; behandlingen skall registreras av den ansvarige veterinären, och minst de upplysningar som anges i punkt 1 skall anges.
Artikel 5
När det gäller vattenbruksdjur kan fiskyngel behandlas med veterinärmedicinska läkemedel med androgen verkan under de tre första månaderna för att erhålla inverterat kön; medicinerna skall vara godkända enligt direktiv 81/851/EEG och 81/852/EEG.
Artikel 6
a) Nedanstående hormonprodukter:
iii) Produkter
- för vilka det inte finns någon reagens eller utrustning som krävs till analysmetoder för att upptäcka förekomst av restsubstanser som överstiger de tillåtna gränserna.
1. I handelssyfte kan medlemsstaterna tillåta avyttring av djur avsedda för avel, eller uttjänta avelsdjur, som under sin aktiva period varit föremål för någon av behandlingarna enligt artikel 4 och 5, samt tillåta anbringande av gemenskapens kontrollmärke på kött från sådana djur, om villkoren i artikel 4 och 5 och om minimal karenstid enligt artikel 6.2 a ii eller b eller karenstiden som avses i avyttringstillståndet respekterats.
Artikel 8
2) Att utöver de kontroller som föreskrivs i direktiv om avyttring av olika produkter i fråga, de officiella kontrollerna enligt artikel 11 i direktiv 96/23/EG (16) genomförs av behöriga nationella myndigheter utan förvarning i syfte att konstatera
c) om karenstider enligt artikel 6 respekteras,
a) förekomst av ämnen som avses under punkt 1 i djur eller djurens dricksvatten, samt på samtliga platser där djuruppfödning eller djurhållning äger rum,
b) visar att kraven under punkt 2 b och 2 c inte iakttagits, skall den behöriga myndigheten vidta lämpliga åtgärder, i proportion till överträdelsens omfattning.
Upplysningarna som avses i första stycket skall på begäran ställas till behörig myndighets förfogande, och om de föreligger i elektronisk form, även som papperskopia.
Artikel 11
a) av husdjur eller vattenbruksdjur
b) av kött eller produkter från djur som enligt punkt a ej får importeras.
Artikel 12
1. Direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG skall upphöra att gälla den 1 juli 1997.
1. Medlemsstaterna skall anta de lagar och andra författningar, i förekommande fall med påföljder, som är nödvändiga för att följa detta direktiv den 1 juli 1997 och vad beträffar â-agonister, senast den 1 juli 1997. De skall genast underrätta kommissionen om detta.
3. Innan bestämmelserna i detta direktiv avseende â-agonister genomförs, skall de nationella reglerna på området vara tillämpliga, varvid allmänna bestämmelser i fördraget skall iakttas.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av följande: I artikel 7a i fördraget föreskrivs ett område utan inre gränser med fri rörlighet för varor, personer, tjänster och kapital.
I meddelande 94/C 138/04 (3) fastställs det förfarande som bör följas av dem (tillverkare eller dennes ombud) som vill att ett gödselmedel skall få betecknas som "EEG-gödselmedel" enligt bilaga II i direktiv 76/116/EEG, genom att lämna i sina tekniska uppgifter till medlemsstatens myndighet. Myndigheten fungerar som rapportör i Europeiska kommissionens arbetsgrupp för gödselmedel.
Artikel 1
Följande produkt och tolerans läggs till under A.1 i bilaga III till direktiv 76/116/EEG:
1. Medlemsstaterna skall anta de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 maj 1997. De skall genast underrätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
Den bästa lösningen består i att tillåta alla medlemsstater att provisoriskt tillämpa en reducerad skattesats för tillhandahållande av jordbruksprodukter från blomster- och trädgårdsodling samt av vedbränsle.
Direktiv 77/388/EEG ändras på följande sätt:
"i) medlemsstaterna får tillämpa en reducerad skattesats för tillhandahållande av levande växter och andra produkter från blomsterodling (inklusive lökar, rötter och liknande produkter, snittblommor och prydnadsbladväxter) liksom för tillhandahållande av vedbränsle."
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100a i detta,
i enlighet med det i artikel 189b i fördraget angivna förfarandet (3), och
3. Den elektricitet som förbrukas av kylskåp och frysar för hushållsbruk utgör en icke obetydlig del av hushållens elförbrukning och därigenom av gemenskapens totala elförbrukning. Elförbrukningen, dvs. energieffektiviteten, varierar kraftigt mellan de olika modeller av kylskåp och frysar med samma volym och egenskaper som erbjuds på gemenskapsmarknaden.
6. Vidtagandet av sådana åtgärder omfattas av gemenskapens befogenheter. Kraven i detta direktiv går inte utöver vad som är nödvändigt för att uppnå direktivets mål och direktivet överensstämmer således med bestämmelserna i artikel 3b i fördraget.
9. I sina slutsatser av den 29 oktober 1990 fastställde rådet målet att till år 2000 stabilisera koldioxidutsläppen (CO2) i gemenskapen på 1990 års nivå. För att nå detta mål krävs kraftigare åtgärder för att stabilisera gemenskapens koldioxidutsläpp.
12. Den energieffektivitetsvinst som automatiskt uppstår till följd av påtryckningar från marknaden och förbättringar av tillverkningsmetoderna och som uppskattas till ungefär 2 % per år, kommer att bidra till ansträngningarna att få till stånd strängare normer för energiförbrukning.
15. Det är viktigt att upprätta ett effektivt verktyg för att säkerställa ett felfritt genomförande av direktivet, rättvisa konkurrensvillkor för tillverkarna och skydd för konsumenternas rättigheter.
18. Kylskåp och frysar för hushållsbruk som överensstämmer med de energieffektivitetskrav som fastställs i detta direktiv skall förses med EG-märkning och tillhörande upplysningar för att möjliggöra deras fria rörlighet.
Artikel 1
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att se till att de kyl- och frysapparater som omfattas av detta direktiv endast får släppas ut på marknaden i gemenskapen om deras elförbrukning är mindre än eller lika med den högsta tillåtna elförbrukningen för denna kategori apparater, vilken skall beräknas enligt de förfaranden som anges i bilaga I.
1. Medlemsstaterna får inte inom sitt respektive territorium förbjuda, begränsa eller hindra att kyl- och frysapparater, försedda med den EG-märkning som intygar att de överensstämmer med samtliga bestämmelser i detta direktiv, släpps ut på marknaden.
b) Om tillverkaren likväl under en övergångsperiod kan välja mellan att tillämpa olika bestämmelser i ett eller flera av dessa direktiv, anger EG-märkningen endast överensstämmelse med bestämmelserna i de direktiv som tillverkaren har tillämpat. I de handlingar, anvisningar och instruktioner som medföljer kyl- och frysapparaterna skall i så fall numren på dessa direktiv anges, enligt den text som offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 5
Artikel 6
Artikel 7
Artikel 8
1. Medlemsstaterna skall anta och offentliggöra de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast inom ett år efter antagandet av detta direktiv. De skall omedelbart underrätta kommissionen om detta.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser de antar inom det område som omfattas av detta direktiv.
KOMMISSIONENS DIREKTIV 96/63/EG av den 30 september 1996 om ändring av rådets direktiv 76/432/EEG om bromsutrustning på jordbruks- eller skogsbrukstraktorer med hjul (Text av betydelse för EES)
med beaktande av rådets direktiv 74/150/EEG av den 4 mars 1974 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av jordbruks- eller skogsbrukstraktorer med hjul (1), senast ändrat genom direktiv 88/297/EEG (2), särskilt artiklarna 12 och 13 i detta, och med beaktande av följande:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
2. Från och med den 1 mars 1998 får medlemsstaterna
för en traktortyp av skäl som hänför sig till bromsutrustningen, om kraven i direktiv 76/432/EEG, ändrat genom detta direktiv, inte är uppfyllda.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 96/73/EG av den 16 december 1996 om vissa metoder för kvantitativ analys av binära textilfiberblandningar
med beaktande av kommissionens förslag (1),
med beaktande av följande: Rådets direktiv 72/276/EEG av den 17 juli 1972 om tillnärmning av medlemsstaternas lagstiftning om vissa metoder för kvantitativ analys av binära textilfiberblandningar (4), har vid ett flertal tillfällen ändrats på väsentliga punkter. Av klarhets- och effektivitetsskäl bör direktivet kodifieras.
Direktivet 96/74/EG föreskriver att den provtagning och de analysmetoder som skall användas i medlemsstaterna för att bestämma fibersammansättningen i varor skall anges i särdirektiv. Följaktligen fastställs i bilaga II till detta direktiv femton enhetliga analysmetoder för de flesta på marknaden förekommande textilvaror som består av binära blandningar.
Bestämmelserna i detta direktiv överensstämmer med det yttrande som avgivits av Kommittén för direktiv om benämningen och märkningen av textilier.
Artikel 1
Analysprov avser ett med hänsyn till analysen lämpligt stort prov, som tas ut från laboratorieprovet, som i sin tur tagits ut från ett varuparti för analys.
Medlemsstaterna skall vidta alla nödvändiga åtgärder för att i enlighet med direktivet 96/74/EG säkerställa att bestämmelserna i bilaga I och II om metoder för den kvantitativa analysen av vissa binära blandningar, inklusive framtagningen av analysprov och provexemplar, tillämpas vid alla officiella provningar för att bestämma sammansättningen av de textilvaror som släpps ut på marknaden.
Artikel 5
3. Anpassning av metoderna för kvantitativ analys till den tekniska utvecklingen enligt bestämmelserna i bilaga II skall ske i enlighet med det förfarande som anges i artikel 6.
2. Kommissionens företrädare skall till kommittén lämna ett förslag om åtgärder som skall beslutas. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande ärendet är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen, varvid medlemsstaternas röster skall vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
Rådet skall besluta med kvalificerad majoritet.
Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Hänvisningar till de upphävda direktiven skall uppfattas som hänvisningar till detta direktiv och läsas enligt jämförelsetabellen i bilaga IV.
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 75 i detta,
i enlighet med det i artikel 189c i fördraget angivna röstningsförfarandet (3), och
För den inre marknadens funktion krävs det i fråga om varutransporter på inre vattenvägar att system med befraktning i turordning anpassas i riktning mot större kommersiell smidighet i syfte att skapa ett system med fri befraktning och fri prissättning för transporter.
Det är viktigt att anta bestämmelser som gör det möjligt att ingripa på den aktuella transportmarknaden om en allvarlig störning skulle inträffa, och för detta ändamål bör kommissionen ges befogenhet att vidta lämpliga åtgärder i enlighet med förfarandet med rådgivande kommitté.
I detta direktiv avses med
c) behörig myndighet: myndighet som av medlemsstaten utsetts att förvalta och organisera systemet med befraktning i turordning,
Inom området nationella och internationella varutransporter på inre vattenvägar inom gemenskapen, skall avtal ingås fritt mellan berörda parter och priser förhandlas fritt.
- att de villkor som räknas upp i artikel 4, 5 och 6 efterlevs, och
Under den övergångsperiod som avses i artikel 3 skall följande undantas från tillämpningsområdet för befraktningssystem i turordning:
- transporter som kräver utrustning för godshantering,
Under den övergångsperiod som avses i artikel 3 skall medlemsstaterna vidta nödvändiga åtgärder för att så långt som möjligt göra systemen med befraktning i turordning mer flexibla, bland annat genom att
Artikel 6
- Tonnageavtal enligt vilket transportören förbinder sig att under en i avtalet fastlagd period transportera ett fastställt antal ton mot betalning av en fraktavgift per ton. Avtalet skall ingås fritt mellan parterna; det måste omfatta betydande godsmängder.
1. Vid allvarlig störning på marknaden får kommissionen, utan att det påverkar tillämpningen av rådets förordning (EEG) nr 1101/89 av den 27 april 1989 om strukturella förbättringar inom inlandssjöfarten (5), på en medlemsstats begäran vidta lämpliga åtgärder, bland annat åtgärder som syftar till att förhindra alla nya ökningar av den transportkapacitet som erbjuds på den ifrågavarande marknaden. Beslutet skall fattas i enlighet med förfarandet i artikel 8.2.
- uppgifter om genomsnittskostnader och priser för olika slags transporter,
Upplysningarna får användas endast i statistiskt syfte. Det är förbjudet att använda dem för beskattningsändamål och att vidarebefordra dem till tredje man.
1. Kommissionen skall biträdas av den kommitté som inrättats genom direktiv 91/672/EEG (6).
Kommissionen skall ta största hänsyn till det yttrande som kommittén avgett. Den skall underrätta kommittén om det sätt på vilket dess yttrande har beaktats.
När en medlemsstat antar dessa bestämmelser, skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras, skall varje medlemsstat själv utfärda.
KOMMISSIONENS FÖRORDNING (EG) nr 242/96 av den 7 februari 1996 om klassificering av vissa varor i Kombinerade nomenklaturen
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 3009/95 (2), särskilt artikel 9 i denna, och med beaktande av följande:
Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapens officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av följande: Rådets förordning (EEG) nr 1014/68 av den 20 juli 1968 om allmänna bestämmelser om offentlig lagring av skummjölkspulver (5), senast ändrad genom förordning (EEG) nr 3577/90 (6), upphörde att gälla från och med den 1 mars 1996 genom rådets förordning (EG) nr 1538/95 (7). Vissa bestämmelser i förordning (EEG) nr 1014/68 har införts i artikel 7 i förordning (EEG) nr 804/68 i dess ändrade lydelse genom förordning (EG) nr 1538/95. Kommissionens förordning (EEG) nr 625/78 av den 30 mars 1978 om tillämpningsföreskrifter för offentlig lagring av skummjölkspulver (8), senast ändrad genom förordning (EG) nr 1802/95 (9), omarbetades när den anpassades till följd av att förordning (EEG) nr 1014/68 upphävdes. Förordning (EEG) nr 625/78 har följaktligen likaså upphört att gälla från och med den 1 mars 1996 genom kommissionens förordning (EG) nr 322/96 av den 22 februari 1996 om tillämpningsföreskrifter för offentlig lagring av skummjölkspulver (10).
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
Förordning (EEG) nr 1362/87 ändras på följande sätt:
b) Punkt e skall ersättas med följande:
Förordning (EEG) nr 1158/91 ändras på följande sätt:
- avseende skummjölkspulver som framställts under de 21 dagarna som omedelbart föregår den sista anbudsdagen; i det fall som avses i bilaga III e andra meningen i förordning (EG) nr 322/96 fastställs denna period till tre veckor,
"c) Det lager dit det skall levereras. Artiklarna 5 och 6 i förordning (EG) nr 322/96 skall tillämpas."
Inom en period som börjar löpa den 120:e dagen efter övertagandet av skummjölkspulvret och som löper ut den 140:e dagen därefter, skall interventionsorganet betala anbudsgivare som tilldelats kontrakt det pris som anges i vederbörandes anbud. Betalning skall ske för varje övertagen kvantitet under förutsättning att kraven i artikel 1 andra stycket är uppfyllda.
- Om proteinhalten i den fettfria torrsubstansen är lägre än 35,6 % men minst 31,4 % skall uppköpspriset vara det pris som anges i anbudet minskat med ett belopp "d" som räknas fram på följande sätt:
Bestämmelserna i artiklarna 2 och 3 i förordning (EG) nr 322/96 skall tillämpas."
>Plats för tabell>
RÅDETS FÖRORDNING (EG) nr 753/96 av den 22 april 1996 om ändring av förordning (EEG) nr 3906/89 i syfte att utvidga det ekonomiska stödet till att omfatta Bosnien-Hercegovina
med beaktande av kommissionens förslag,
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I artikel 39 i förordning (EEG) nr 1785/81 anges att medlemsstaterna och kommissionen skall lämna varandra de uppgifter som behövs för tillämpningen av förordningen. Således fastställdes tillämpningsbestämmelser i kommissionens förordning (EEG) nr 787/83 av den 29 mars 1983 om informationslämnande inom sockersektorn (3), senast ändrad genom förordning (EEG) nr 3819/85 (4). Med tanke på den utveckling som sedan skett av den gemensamma organisationen av marknaden för socker och särskilt gemenskapens åtaganden till följd av det jordbruksavtal som slöts efter Uruguayrundans multilaterala förhandlingar, finns det anledning att se över bestämmelserna i sin helhet och fastställa nya och att upphäva förordning (EEG) nr 787/83 inför regleringsåret 1996/97.
För att det kvoteringssystem som fastställts i avdelning III i förordning (EEG) nr 1785/81 skall fungera effektivt, är det nödvändigt att ha tillgång till all relevant information, särskilt med hänsyn till gemenskapens åtaganden inom ramen för nämnda jordbruksavtal. Detta berör tillämpningen av rådets förordning (EEG) nr 206/68 av den 20 februari 1968 om rambestämmelser för avtal och branschöverenskommelser rörande inköp av betor (19), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige, rådets förordning (EEG) nr 193/82 av den 26 januari 1982 om allmänna bestämmelser för överföring av kvoter inom sockersektorn (20), kommissionens förordning (EEG) nr 2670/81 av den 14 september 1981 om fastställande av tillämpningsföreskrifter för sockerproduktion utöver kvoten (21), senast ändrad genom förordning (EG) nr 158/96 (22), samt kommissionens förordning (EEG) nr 1443/82 av den 8 juni 1982 om tillämpningsföreskrifter för kvotsystemet på sockerområdet (23), senast ändrad genom förordning (EEG) nr 392/94 (24). Ovanstående gäller också för det system för kompensation för lagringskostnader som fastställts i artikel 8 i förordning (EEG) nr 1785/81. Därvid berörs tillämpningen av rådets förordning (EEG) nr 1358/77 av den 20 juni 1977 om allmänna bestämmelser för kompensation för lagringskostnader för socker, samt om upphävande av förordning (EEG) nr 750/68 (25), senast ändrad genom förordning (EEG) nr 3042/78 (26), liksom kommissionens förordning (EEG) nr 1998/78 av den 18 augusti 1978 om tillämpningsföreskrifter för kompensation för lagringskostnader för socker (27), senast ändrad genom förordning (EEG) nr 1758/93 (28).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som erbjudits men ännu inte tagits över av interventionsorganet,
Artikel 2
Vad gäller interventionsåtgärder som vidtagits i enlighet med artikel 9.2 i förordning (EEG) nr 1785/81 skall varje medlemsstat till kommissionen anmäla följande:
Artikel 4
a) en licens om produktionsbidrag har utfärdats,
a) en licens om produktionsbidrag har utfärdats,
Artikel 5
a) de kvantiteter för vilka licens har utfärdats med angivande av motsvarande exportbidrag fastställda i enlighet med artikel 17.5 andra stycket a i förordning (EEG) nr 1785/81, angivna var för sig enligt följande:
- sackarossirap uttryckt som vitsocker KN-nr 1702 60 90, 1702 90 60, 1702 90 71, 1702 90 99 och 2106 90 59,
b) de kvantiteter vitsocker KN-nr 1701 99 10 för vilka licens har utfärdats med angivande av motsvarande exportbidrag fastställda i enlighet med artikel 17.5 andra stycket b i förordning (EEG) nr 1785/81,
2. Senast i slutet av varje kalendermånad, med avseende på närmast föregående kalendermånad, de kvantiteter vitsocker enligt punkt 1 b som exporterats i enlighet med artikel 8.4 och 8.5 i förordning (EEG) nr 3719/88.
b) de kvantiteter socker ur kvoten som exporterats som vitsocker eller som bearbetad produkt uttryckt som vitsocker, för vilka exportlicens har utfärdats med anledning av livsmedelbistånd i gemenskapens eller nationell regi inom ramen för internationella överenskommelser eller andra kompletterande program eller till följd av andra åtgärder inom gemenskapen som avser kostnadsfri livsmedelstilldelning,
e) för export enligt 1 d och d i denna punkt de kvantiteter som exporterats utan bidrag.
Varje medlemsstat skall till kommissionen anmäla följande:
a) importerats från tredje land i form av bearbetade produkter enligt 5.1 d och 5.3 d,
Varje medlemsstat skall till kommissionen anmäla följande:
Artikel 8
2. Att senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, till kommissionen vidarebefordra
c) kopior, i förekommande fall, av den deklaration som avses i artikel 1.3 andra stycket i förordning (EEG) nr 2782/76.
a) den totala kvantiteten vitsocker, angiven i ton,
som importerats i enlighet med förordning (EEG) nr 2782/76 till medlemsstaten under den leveransperiod som löper ut den 30 juni i frågavarande år.
1. Före den 1 mars varje år, med avseende på vart och ett av de sockerproducerande företagen och de företag som framställer inulinsirap, vilka är belägna på dess territorium, anmäla den beräknade socker- och inulinsirapproduktionen under det löpande regleringsåret fastställd i enlighet med artikel 3.1 i förordning (EEG) nr 1443/82. För de franska departementen Guadeloupe och Martinique samt för Spanien skall när det gäller rörsocker emellertid denna dag ersättas med den 1 juli.
Artikel 10
b) de kvantiteter socker som har denaturerats,
Artikel 12
2. Före den 1 mars varje år, med avseende på det löpande regleringsåret och för vart och ett av de sockerproducerande företagen, anmäla de totala kvantiteter B-socker och C-socker som förts över till påföljande regleringsår.
Artikel 13
2. Före den femtonde dagen i varje månad, med avseende på den näst senaste kalendermånaden och på det sätt som framgår av exemplet i bilaga I anmäla
Artikel 14
2. Före den 1 oktober efter varje regleringsår och med avseende på det regleringsåret uppgifter rörande försörjningsbalansen för melass enligt exemplet i bilaga III.
Artikel 16
b) närmast föregående kvartal: den tre månader långa referensperioden juli-september, oktober-december, januari-mars eller april-juni, allt efter vad som är aktuellt,
Kommissionen skall se till att den information som har överlämnats till den i enlighet med denna förordning blir tillgänglig för medlemsstaterna.
Artikel 19
KOMMISSIONENS FÖRORDNING (EG) nr 2214/96 av den 20 november 1996 om harmoniserade konsumentprisindex: överföring och spridning av HIKP:s delindex (Text av betydelse för EES)
med beaktande av rådets förordning (EG) nr 2494/95 av den 23 oktober 1995 om harmoniserade konsumentprisindex (1), och
I artikel 11 i förordning (EG) nr 2494/95 krävs att HIKP och motsvarande delindex skall publiceras av kommissionen (Eurostat). Dessa delindex behöver specifieras.
Enligt artikel 5.3 i förordning (EG) nr 2494/95 har samråd skett med Europeiska monetära institutet som har avgett ett positivt yttrande.
Mål
Definitioner
Framtagande och överföring av delindex
Spridning av delindex
Kvalitetskontroll
Ikraftträdande
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av följande: Identifieringssystemet skall vara frivilligt, åtminstone i ett inledande skede, men det skall genomgå en översyn för att fastställa om det skall införas på obligatorisk grund i ett senare skede.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
- Kompositmaterial betecknar förpackningar gjorda av olika material som inte kan separeras för hand och som inte i något fall överstiger en viss viktprocent som skall fastställas enligt det förfarande som anges i artikel 21 i direktiv 94/62/EG. Eventuella undantag för vissa material får fastställas genom samma förfarande.
Användningen av dessa skall vara frivillig när det gäller de plastmaterial som anges i bilaga I, papper och papp som anges i bilaga II, de metaller som anges i bilaga III, de trämaterial som anges i bilaga IV, de textilmaterial som anges i bilaga V, de glasmaterial som anges i bilaga VI och de kompositmaterial som anges i bilaga VII.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av följande: För att kunna fastställa bruttonationalinkomsten till marknadspris (BNImp) i enlighet med artikel 1 i direktiv 89/130/EEG, Euratom, som enligt artikel 8.1 i rådets förordning (EG) nr 2223/96 av den 25 juni 1996 om det europeiska national- och regionalräkenskapssystemet i gemenskapen (2) skall fortsätta att tillämpas så länge som beslut 94/728/EG, Euratom (3) gäller, är det nödvändigt att klargöra principerna för inkomst från institut för kollektiv investering i enlighet med gällande upplaga av Europasystemet för integrerad ekonomisk redovisning (ENS).
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som inrättas genom artikel 6 i direktiv 89/130/EEG, Euratom,
För tillämpning av direktiv 89/130/EEG, Euratom skall inkomst från institut för kollektiv investering definieras dels som erhållen ränta från inlåning och värdepapper, dels som utdelning på aktier vilka innehas av instituten för kollektiv investering. Denna inkomst kan delas ut till aktieägare eller läggas till kapitalet.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
Kommissionen skall välja det av de två förfaranden enligt artikel 13.3 i direktiv 89/106/EEG för bestyrkande av överensstämmelse av en produkt, som är "minst betungande och samtidigt förenligt med kraven på säkerhet". Detta innebär att det är nödvändigt att besluta huruvida en tillverkningskontroll i fabriken under tillverkarens ansvar är erforderlig och tillräcklig för bestyrkande av överensstämmelse för en bestämd produkt eller produktgrupp, eller om det av orsaker som rör uppfyllandet av de kriterier som avses i artikel 13.4 krävs att ett godkänt certifieringsorgan deltar.
Det förfarande som avses i artikel 13.3 a motsvarar de system som anges i det första alternativet utan fortlöpande övervakning, samt i det andra och det tredje alternativet i punkt 2 ii i bilaga III och det förfarande som avses i artikel 13.3 b motsvarar de system som anges i punkt 2 i i bilaga III samt i det första alternativet med fortlöpande övervakning i punkt 2 ii i bilaga III.
Artikel 1
För de produkter som anges i bilaga II skall överensstämmelsen bestyrkas genom ett förfarande där, förutom ett tillverkningskontrollsystem i fabriken som genomförs av tillverkaren, även ett godkänt certifieringsorgan deltar vid bedömningen och övervakningen av tillverkningskontrollen eller av själva produkten.
Artikel 4
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Den första meningen i artikel 6.1 skall ersättas med följande:
"Efter utgången av treårs- eller tvåårsperioden skall medlemmarna, ordföranden och vice ordföranden sitta kvar tills de ersätts eller deras mandat förnyas."
Medlemmarna skall åta sig att undvika alla intressekonflikter under det att de utövar sina uppdrag."
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Pistaschmandlar som har sitt ursprung i Iran eller som försänds från Iran har i många fall visat sig innehålla alltför höga halter av aflatoxin B1.
De undersökningar som genomförts av de hygieniska förhållandena i Iran har visat att det krävs förbättrad hygienpraxis, och att pistaschmandlarna måste kunna spåras. Undersökningsgruppen lyckades inte kontrollera alla steg i hanteringen av pistaschmandlarna för export. De iranska myndigheterna har dock gjort åtaganden, i synnerhet beträffande förbättringar i fråga om produktion, hantering, sortering, bearbetning, förpackning och transport. Därför är det lämpligt att pistaschmandlar och produkter som är framställda av dessa, som har sitt ursprung i eller försänds från Iran, underkastas vissa särskilda villkor i syfte att säkerställa en hög skyddsnivå för folkhälsan.
De iranska myndigheterna måste tillhandahålla dokumenterade bevis rörande villkoren för produktion, sortering, hantering, bearbetning, förpackning och transport samt resultaten av laboratorieundersökningar av sändningen beträffande halten av aflatoxin B1 och den totala aflatoxinhalten; denna dokumentation måste åtfölja varje sändning av pistaschmandlar som har sitt ursprung i Iran eller som försänds från Iran.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
- rostade pistaschmandlar som omfattas av KN-numren 2008 19 13 och 2008 19 93,
3. Varje sändning skall identifieras med en kod som motsvarar koden på provtagnings- och analysresultaten från den officiella provtagningen och analysen, och på det hälsointyg som avses i punkt 1.
Artikel 3
Medlemsstaterna skall vidta de åtgärder som krävs för att följa detta beslut. De skall underrätta kommissionen om detta.
KOMMISSIONENS DIREKTIV 97/37/EG av den 19 juni 1997 om anpassning av bilaga I och II till Europaparlamentets och rådets direktiv 96/74/EG om benämningar på textilier till den tekniska utvecklingen (Text av betydelse för EES)
med beaktande av Europaparlamentets och rådets direktiv 96/74/EG av den 16 december 1996 om benämningar på textilier (1), särskilt artikel 16.1 i detta, och
Endast textilfibrerna i förteckningen i bilaga I till nämnda direktiv får användas vid sammansättning av textilprodukter som är avsedda för gemenskapens inre marknad. Det är nödvändigt att anpassa bilagornas förteckningar över fibrer till den tekniska utvecklingen genom att tillföra nya fibrer som har införts på marknaden efter den senaste ändringen av direktivet.
Artikel 1
- I kolumnen "beteckning" förs "kashgora" in efter "guanaco".
- Texten i kolumnen "beteckning" skall vara "polyamid eller nylon".
"fiber bildad av syntetiska linjära makromolekyler bestående av aromatiska grupper som binds samman med amid- eller imidbindningar, av vilka minst 85 % binds direkt till två aromatiska ringar och där imidbindningarna, om sådana finns, till antalet inte får överskrida antalet amidbindningar."
6) Ett nytt nr 33 införs enligt följande:
"Med `organiskt lösningsmedel` avses en blandning av organiska ämnen och vatten."
Bilaga II till direktiv 96/74/EEG ändras på följande sätt:
Texten i kolumnerna "benämning" och "procentsatser" skall vara följande:
Texten i kolumnerna "benämning" och "procentsatser" skall vara följande:
Texten i kolumnerna "benämning" och "procentsatser" skall vara följande:
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa direktiv 96/74/EG senast den 1 juni 1998.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 97/52/EG av den 13 oktober 1997 om ändring av direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG om samordning av förfarandena vid tilldelning av kontrakt vid offentlig upphandling av tjänster, varor samt bygg- och anläggningsarbeten
med beaktande av kommissionens förslag (1),
med beaktande av följande: 1. Genom sitt beslut 94/800/EG av den 22 december 1994 om ingående, på Europeiska gemenskapens vägnar - såvitt avser frågor som omfattas av dess behörighet - av de överenskommelser som är resultatet av de multilaterala förhandlingarna inom Uruguayrundan (1986 1994) (4) godkände rådet på Europeiska gemenskapens vägnar bland annat avtalet om offentlig upphandling, nedan kallat "avtalet", vars syfte är att införa ett multilateralt system av väl avvägda rättigheter och skyldigheter när det gäller offentlig upphandling för att liberalisera och utvidga världshandeln. Detta avtal har inte direkt effekt.
4. Med tanke på de internationella rättigheter och åtaganden som ett godtagande av avtalet medför för Europeiska gemenskapen, bör det system som tillämpas på anbudsgivare och varor från tredje land som undertecknat avtalet vara det som anges i avtalet, vars räckvidd när det gäller direktiv 92/50/EEG inte omfattar tjänstekontrakt enligt bilaga I B, kontrakt om forsknings- och utvecklingstjänster enligt kategori 8 i bilaga I A därtill, kontrakt om telekommunikationstjänster enligt kategori 5 i bilaga I A därtill med referensnummer enligt den allmänna klassificeringen av produkter (CPC) 7524, 7525 och 7526 eller kontrakt om finansiella tjänster enligt kategori 6 i bilaga I A därtill i samband med utfärdande, försäljning, förvärv eller överförande av värdepapper eller andra finansiella instrument samt i samband med tjänster som utförs av centralbanker.
7. Det är därför nödvändigt att anpassa och komplettera bestämmelserna i direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG.
10. Upphandlande myndigheter får begära eller ta emot råd som kan användas för att upprätta specifikationer för ett bestämt upphandlingsförfarande under förutsättning att dessa råd inte hindrar konkurrensen.
Artikel 1
- de offentliga kontrakt avseende tjänster som avses i artikel 3.3, de offentliga kontrakt avseende sådana tjänster som avses i bilaga I B, tjänster i kategori 8 i bilaga I A och telekommunikationstjänster i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, förutsatt att det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 200 000 ecu,
ii) som tilldelas av de upphandlande myndigheter som anges i artikel 1 b utom dem som nämns i bilaga I till direktiv 93/36/EEG och vilkas uppskattade värde, exklusive mervärdesskatt, uppgår till minst 200 000 SDR i ecu.
c) De tröskelvärden som framgår av a och deras motvärden uttryckta i ecu och i nationella valutor skall offentliggöras i Europeiska gemenskapernas officiella tidning i början av november månad efter den revision som anges i b i det här stycket.
2. Artikel 12.1 och 12.2 ersätts med följande text:
2. De upphandlande myndigheterna skall så snart som möjligt underrätta de anbudssökande och anbudsgivarna om de beslut som fattas rörande tilldelningen av kontrakt, inklusive skälen till att de har beslutat att avstå från en upphandling för vilken anbud begärts eller att upprepa förfarandet; dessa upplysningar skall på begäran lämnas skriftligen. Myndigheterna skall även underrätta Byrån för Europeiska gemenskapernas officiella publikationer om dessa beslut."
- det tröskelvärde som avses i artikel 7.1 a första strecksatsen för de tjänster som avses i bilaga I B, tjänsterna i kategori 8 i bilaga I A och telekommunikationstjänsterna i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, eller
2. Denna artikel skall tillämpas på alla formgivningstävlingar där det sammanlagda beloppet av tävlingspriserna och ersättningarna till deltagarna uppgår till minst
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen ii för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, utom dem som nämns i bilaga I till direktiv 93/36/EEG."
5. Artikel 19.4 ersätts med följande text:
"2. Anbud skall avges skriftligen, direkt eller per post. Medlemsstaterna får tillåta avgivande av anbud på alla andra sätt som gör det möjligt att säkerställa
- om det är nödvändigt av bevisskäl, att anbud så snart som möjligt bekräftas skriftligen eller genom översändande av en bestyrkt kopia,
"Artikel 38a
a) När det gäller de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG
b) När det gäller övriga upphandlande myndigheter som avses med detta direktiv, antal och värden för kontrakt som av varje kategori av upphandlande myndighet tilldelas över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, tjänstekategori i enlighet med den terminologi som anges i bilaga I och nationalitet för den tjänsteleverantör som tilldelas kontraktet samt, i fråga om förhandlade förfaranden, med uppdelning enligt artikel 11 under angivande av antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
De statistiska rapporter som begärs enligt denna punkt skall inte avse kontrakt som rör tjänster i kategori 8 i bilaga I A, telekommunikationstjänster i kategori 5 i bilaga I A, med CPC-referensnumren 7524, 7525 och 7526, eller tjänster i enlighet med bilaga I B, förutsatt att deras uppskattade värde, exklusive mervärdesskatt, är mindre än 200 000 ecu.
Artikel 2
A) ersätts punkt 1 med följande text:
ii) de upphandlande myndigheterna som anges i bilaga I, om det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 130 000 SDR i ecu. När det gäller upphandlande myndigheter inom försvarssektorn skall detta gälla bara för upphandling av produkter enligt bilaga II.
Den beräkningsmetod som anges i detta stycke skall på förslag av kommissionen ses över av Rådgivande kommittén för offentlig upphandling i princip två år efter det att den tillämpats för första gången.
"7. De upphandlande myndigheterna skall se till att det inte förekommer någon diskriminering mellan olika leverantörer."
De upphandlande myndigheterna får emellertid besluta att viss information som rör tilldelningen av kontrakt och som nämns i första stycket inte skall lämnas ut om det bedöms att detta skulle hindra lagarnas tillämpning eller strida mot allmänintresset eller vara till skada för offentliga eller privata företags legitima kommersiella intressen eller för lojal konkurrens mellan tjänsteleverantörer.
"1 a. Tidsfristen för mottagande av anbud enligt punkt 1 får ersättas av en tidsfrist som är tillräckligt lång för att de berörda parterna skall ha möjlighet att avge giltiga anbud, och som i allmänhet inte skall understiga 36 dagar, men som aldrig skall vara kortare än 22 dagar räknat från dagen för avsändande av meddelandet om upphandling, om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 9.1, utformat enligt förlagan i bilaga IV A (förhandsinformation) till Europeiska gemenskapernas officiella tidning åtminstone 52 dagar och högst tolv månader före insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 9.2, och om förhandsmeddelandet dessutom innehåller åtminstone den information som föreskrivs i förlagan i bilaga IV B (öppet förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
5. I artikel 15 skall följande punkt läggas till:
- att anbudets sekretess består i avvaktan på utvärderingen, och
1. Kommissionen skall i samråd med Rådgivande kommittén för offentlig upphandling granska hur detta direktiv tillämpas, och den skall vid behov lägga fram nya förslag för rådet, särskilt i syfte att samordna medlemsstaternas åtgärder för att följa detta direktiv.
1. För att möjliggöra en bedömning av resultatet av tillämpningen av detta direktiv skall medlemsstaterna till kommissionen översända en statistisk rapport rörande de varukontrakt som under det föregående året tilldelats av de upphandlande myndigheterna, senast den 31 oktober 1996, och när det gäller de upphandlande myndigheter som inte anges i bilaga I, senast den 31 oktober 1997 och därefter senast den 31 oktober varje år.
- det beräknade sammanlagda värdet för kontrakt som av varje upphandlande myndighet tilldelas under tröskelvärdet,
c) När det gäller de upphandlande myndigheter som avses i bilaga I, antal och sammanlagt värde för kontrakt som tilldelas av varje upphandlande myndighet enligt undantagen från avtalet. När det gäller övriga upphandlande myndigheter som omfattas av detta direktiv, det sammanlagda värdet för kontrakt som tilldelas av varje kategori av upphandlande myndighet enligt undantagen från avtalet.
8. Bilaga I ersätts med den text som framgår av bilaga I till det här direktivet, och bilaga IV ersätts med den text som framgår av bilaga III till det här direktivet.
1. I artikel b
a) offentliga bygg- och anläggningsarbeten med ett uppskattat värde, exklusive mervärdesskatt, som uppgår till minst 5 000 000 särskilda dragningsrätter (SDR) i ecu.
Det tröskelvärde som bestäms i punkt 1 och dettas motvärde uttryckt i ecu och i nationella valutor skall offentliggöras i Europeiska gemenskapernas officiella tidning i början av november efter den revision som avses i första stycket.
"6. De upphandlande myndigheterna skall se till att det inte förekommer någon diskriminering mellan olika entreprenörer."
De upphandlande myndigheterna får emellertid besluta att viss information som rör tilldelningen av kontrakt och som nämns i första stycket inte behöver lämnas ut om det bedöms att detta skulle hindra lagarnas tillämpning eller strida mot allmänintresset eller vara till skada för offentliga eller privata företags legitima kommersiella intressen eller för en sund konkurrens mellan entreprenörer.
"2. Tidsfristen för mottagande av anbud enligt punkt 1 får ersättas av en tidsfrist som är tillräckligt lång för att de berörda parterna skall ha möjlighet att avge giltiga anbud, och som i allmänhet inte skall understiga 36 dagar, men som aldrig skall vara kortare än 22 dagar räknat från dagen för avsändandet av meddelandet om upphandling om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 11.1, utformat enligt förlagan i bilaga IV A (förhandsinformation), till Europeiska gemenskapernas officiella tidning åtminstone 52 dagar och högst tolv månader före insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 11.2, och om detta meddelande dessutom innehåller minst den information som föreskrivs i förlagan i bilaga IV B (öppet förfarande), förutsatt att denna information var tillgänglig vid tidpunkten för meddelandets offentliggörande."
5. I artikel 18 blir den befintliga texten punkt 1 och följande punkt läggs till:
- att anbudets sekretess består i avvaktan på utvärderingen, och
6. Följande artikel förs in:
2. Den statistiska rapporten skall åtminstone innehålla följande:
- antal och värden för kontrakt som tilldelats av varje upphandlande myndighet över tröskelvärdet, med uppdelning, så långt som möjligt, efter förfarande, kategori av bygg- och anläggningsarbeten i enlighet med den terminologi som används i bilaga II och nationaliteten hos den entreprenör som tilldelats kontraktet samt, i fråga om förhandlande förfaranden, fördelat enligt artikel 7 med uppgift om antal och värden för de kontrakt som tilldelats varje medlemsstat och tredje land.
d) Alla andra statistiska upplysningar som skall bestämmas i enlighet med förfarandet i artikel 35.3 och som begärs i överensstämmelse med avtalet.
Artikel 4
2. Medlemsstaterna skall till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som regleras av det här direktivet samt en jämförelsetabell över bestämmelserna i detta direktiv och de antagna nationella bestämmelserna.
KOMMISSIONENS FÖRORDNING (EG) nr 142/97 av den 27 januari 1997 om lämnande av uppgifter om vissa existerande ämnen i enlighet med rådets förordning (EEG) nr 793/93 (Text av betydelse för EES)
med beaktande av rådets förordning (EEG) nr 793/93 av den 23 mars 1993 om bedömning och kontroll av risker med existerande ämnen (1), särskilt artikel 12.2 i denna, och med beaktande av följande:
Med beaktande av kommissionens förordning (EEG) nr 1488/94 (2) om principer för bedömning av risker för människor och miljö av existerande ämnen i enlighet med förordning (EEG) nr 793/93.
Artikel 1
- människor avser arbetstagare, konsumenter och andra som kommer i kontakt med ämnet via miljön,
Artikel 2
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EG) nr 1256/96 av den 20 juni 1996 om tillämpningen av en flerårig ordning med allmänna tullförmåner under perioden 1 juli 1996-30 juni 1999 för vissa jordbruksprodukter med ursprung i utvecklingsländerna (2), särskilt artikel 12.3 i denna,
med beaktande av Ekonomiska och sociala kommitténs yttrande (5), och
Den 7 juni 1995 ingav Fria fackföreningsinternationalen (ICFTU) och Europeiska fackliga samorganisationen (ETUC) ett gemensamt klagomål enligt artikel 9 i förordning (EG) nr 3281/94 till kommissionen och begärde ett tillfälligt upphävande av gemenskapens system med allmänna tullförmåner för Myanmar på grund av dess användning av tvångsarbete.
Myanmars myndigheter har officiellt underrättats om att undersökningen har inletts. De bestrider att de metoder som avses i klagomålet utgör tvångsarbete med hänvisning till de undantag som avses i artikel 2.2 i ILO:s konvention nr 29 och hävdar att dessa undantag omfattas av 1907 års Town Act och 1908 års Village Act enligt vilka det är tillåtet att ålägga befolkningen att utföra arbeten och tjänster. ILO bestrider denna tolkning och dess behöriga organ har begärt att lagarna i fråga snarast skall upphävas i syfte att göra dessa lagar förenliga med andan och ordalydelsen i konvention nr 29.
All den bevisning som kommissionen har inhämtat i den undersökning som den har utfört efter ICFTU:s och ETUC:s ursprungliga klagomål samt de slutsatser som den har dragit på grundval av dessa uppgifter är tillräckligt omfattande för att utgöra ett välgrundat underlag för prövningen av det utvidgade klagomål som har inlämnats av dessa organisationer den 2 januari 1997. Detta gör det onödigt med en särskild undersökning för jordbrukssektorn. Kraven i artikel 9.2 i förordning (EG) nr 1256/96 är sålunda uppfyllda och villkoren i artikel 11.5 i den förordningen är uppfyllda.
Det faktum att de fördömda metoderna varit rutinmässiga och omfattande gör att det är befogat att helt upphäva bestämmelserna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Vad gäller produkter bör uttrycken "inte saluförts" och "återtagits från marknaden" likställas och ingå i samma definition. Det är också lämpligt att förtydliga att för produkter som återtas från marknaden behöver förpackningskraven inte vara uppfyllda.
I artikel 28 i förordning (EG) nr 2200/96 förskrivs att medlemsstaterna måste meddela de priser som noteras på de representativa marknaderna för vissa bestämda produkter och för vissa perioder. Följaktligen bör en förteckning upprättas över dessa marknader och över berörda produkter.
Det är lämpligt att fastställa, i enlighet med vad som förskrivs i artikel 25 i förordning (EG) nr 2200/96, de frister för att framlägga de åtgärder som medlemsstaterna vidtar för att skydda miljön vid återtagande.
De bestämmelser som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för frukt och grönsaker samt från Kommittén för den europeiska utvecklings- och garantifonden för jordbruket.
I denna förordning fastställs tillämpningsföreskrifter för interventionsordning som avses i avdelningen IV i förordning (EG) nr 2200/96, och gäller för de produkter som avses i artikel 1.2 i den förordningen.
2. Produkterna som återtagits från marknaden bör överensstämma med gällande normer om sådana normer har fastställts i enlighet med artikel 2 i förordning (EG) nr 2200/96. I detta fall är dock normerna för förpackning inte tillämpliga.
a) medlemmarnas produktion som faktiskt sålts genom eller bearbetats av producentorganisationen,
Den saluförda kvantitet som avses i första stycket omfattar inte den produktion som saluförts av de av producentorganisationens medlemmar som får sälja i enlighet med artikel 11.1 c.3 andra och tredje strecksatsen i förordning (EG) nr 2200/96.
Regleringsåren för produkter som omfattas av gemenskapskompensation för återtagande i enlighet med artikel 23.3 i förordning (EG) nr 2200/96 anges i bilaga I till denna förordning.
2. Ansökan som avses i punkt 1 skall minst gälla en period om en månad. Den skall åtföljas av dokument som intygar kvantiteten av varje saluförd produkt och kvantiteten av varje produkt som inte saluförts genom producentorganisationen samt innehåller detaljerade uppgifter om
c) den produktion som tillförts av var och en av de odlare som inte tillhör någon producentorganisation enligt villkoren i artikel 24 i förordning (EG) nr 2200/96.
Utan att det påverkar tillämpningen av artikel 22 i denna förordning när det gäller utbetalning av kompensation för återtagande av produkter som inte anges i bilaga II till förordning (EG) nr 2200/96 samt utbetalning av det tillägg till gemenskapens ersättning för återtagande som föreskrivs i artikel 15.3 a och 15.3 b i förordning (EG) nr 2200/96, skall bestämmelserna i förordning (EG) nr 411/97 tillämpas.
2. Medlemsstaterna skall en gång i veckan på elektronisk väg meddela kommissionen de på de representativa marknaderna för varje marknadsdag noterade dagspriserna för de produkter och för de perioder som anges i bilaga III till denna förordning. Kommissionen skall vidarebefordra dessa upplysningar till medlemsstaterna.
2. Följande uppgifter skall av producentorganisationerna eller deras sammanslutningar meddelas till medlemsstaterna, vilka i sin tur skall vidarebefordra dem till kommissionen:
Artikel 9
a) senast den 30 juni som följer på varje regleringsår för tomater, auberginer, blomkål, aprikoser, persikor, nektariner, vindruvor, meloner och vattenmeloner samt för produkter utanför bilaga II till förordning (EG) nr 2200/96, och
Artikel 10
2. För att kunna bli godkända skall välgörenhetsorganisationerna förbinda sig att
c) underkasta sig de kontroller som föreskrivs av gemenskapsrätten.
Medlemsstaterna skall till kommissionen lämna in förteckningar över de godkända välgörenhetsorganisationer som avses i första stycket b och c och kommissionen skall i sin tur se till att de offentliggörs i Europeiska gemenskapernas officiella tidning, serie C.
Artikel 13
Artikel 14
Artikel 15
2. Transportkostnaderna skall betalas till den avsändare som faktiskt har burit transportkostnaderna i fråga.
- kvantiteten av aktuella produkter,
Artikel 16
3. Dessa avtal får slutas på villkor att det finns produkter som återtagits från marknaden. Kvantiteterna som anges i avtalen får med hänsyn till situationen på marknaden ökas under regleringsåret.
- de planerade transportmedlen,
- kravet att producentorganisationen tillhandahåller produkter som storlekssorterats på förhand och förpackats i emballage med en vikt på högst 25 kg.
6. Ersättning för sorterings- och förpackningskostnader skall utbetalas till de producentorganisationer som har sorterat och förpackat produkterna och skall utgå på villkor att intyg läggs fram som bekräftar
- de faktiska kostnaderna för förpackning och sortering,
1. Medlemsstaterna skall vidta alla nödvändiga åtgärder för att säkerställa att bestämmelserna i avdelning IV i förordning 2200/96 efterlevs, särskilt de som föreskrivs i punkterna 2, 3 och 4.
Vid tillämpning av artikel 30.2 i förordning (EG) nr 2200/96, skall medlemsstaterna kontrollera alla återtagna kvantiteter.
4. Om kontrollerna visar på väsentliga oriktigheter skall de behöriga myndigheterna genomföra ytterligare kontroller det pågående regleringsåret och öka antalet kontroller det påföljande regleringsåret.
b) välgörenhetsorganisationernas slutliga användning av produkterna, särskilt genom att kräva av dessa ett övertagandeintyg som intygar användningen av produkterna, och
3. Beträffande utdelning inom gemenskapen och utan att det påverkar bestämmelserna i artikel 39 i förordning (EG) nr 2200/96 skall de behöriga nationella myndigheterna genomföra kontroller av produkternas användning och slutliga bestämmelse på det territorium där gratisutdelningen sker.
1. Den som mottar gemenskapernas kompensation för återtagande eller finansiering genom driftsfonden är skyldig att återbetala dubbelt så mycket som de belopp som felaktigt betalats ut plus ränta för den tid som förflutit mellan utbetalningen och mottagarens återbetalning om det vid kontroll enligt artikel 17 visar sig att
c) avsättningen av produkter som inte saluförts medför allvarliga skador för miljön.
Artikel 20
3. De institutioner som anges i artikel 12 har inte rätt till gratis utdelning under nästa regleringsår.
6. Räntesatsen för denna ränta skall vara den som tillämpas av Europeiska monetära institutet för dess transaktioner i ecu som offentliggörs i Europeiska gemenskapernas officiella tidning C-serien, och som gäller den dag den felaktiga utbetalningen gjordes, ökad med tre procentenheter.
Artikel 22
Förordningarna (EEG) nr 3587/86, (EEG) nr 827/90, (EEG) nr 2103/90, (EEG) nr 2276/92 samt (EG) nr 113/97 upphör att gälla.
KOMMISSIONENS FÖRORDNING (EG) nr 888/97 av den 16 maj 1997 om ändring av vissa bestämmelser i de normer som fastställts för färsk frukt och färska grönsaker
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker (1), särskilt artiklarna 2.2 och 10 i denna, och
I Ekonomiska kommissionens för Europa internationella normer för färsk frukt och färska grönsaker fastställs tydligt hur packaren och avsändaren skall anges på förpackningen. Dessa internationella bestämmelser bör, i synnerhet för den juridiska tydlighetens skull, införlivas i gemenskapens alla normer för färsk frukt och färska grönsaker.
I rådets förordning nr 211/66/EEG av den 14 december 1966 om utökning av de gemensamma kvalitetsnormerna för vissa frukt och grönsaksslag med en kompletterande kvalitetsklass (2), senast ändrad genom kommissionens förordning (EEG) nr 3596/90 (3), fastställs också en kategori III för blomkål. Av samma skäl som ovan bör förordning nr 211/66/EEG upphävas.
a) i de förordningar som anges i bilaga I skall ändras på följande sätt:
b) i de förordningar som anges i bilaga II skall ändras på följande sätt:
2. I de förordningar som anges i bilaga III skall all hänvisning till kategori III utgå.
Denna förordning träder i kraft den 1 juli 1997.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
För att åstadkomma en enhetlig tillämpning av den Kombinerade nomenklatur som intagits i bilagan till ovannämnda förordning bör bestämmelser antas avseende klassificering av de varor som intagits i bilagan till den här förordningen.
Om inte annat följer av gällande bestämmelser i gemenskapen avseende systemet för dubbelkontroll samt övervakning på gemenskapsnivå, i förväg eller i efterhand, av textilvaror som importeras till gemenskapen, är det lämpligt att bindande tulltaxeupplysningar i fråga om klassificering av varor i Kombinerade nomenklaturen som lämnats av tullmyndigheterna i medlemsstaterna och som inte överensstämmer med den här förordningen får fortsätta att åberopas av innehavaren under en period av 60 dagar, i enlighet med bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen (3), senast ändrad genom förordning (EG) nr 82/97 (4).
Artikel 1
Om inte annat följer av gällande bestämmelser i gemenskapen avseende systemen för dubbelkontroll samt övervakning på gemenskapsnivå, i förväg eller i efterhand, av textilvaror som importeras till gemenskapen får bindande tulltaxeupplysningar i fråga om klassificering av varor i Kombinerade nomenklaturen, som lämnats av tullmyndigheterna i medlemsstaterna och som inte överensstämmer med den här förordningen, fortsätta att åberopas, i enlighet med bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 under en period av 60 dagar.
KOMMISSIONENS FÖRORDNING (EG) nr 1059/97 av den 11 juni 1997 om anpassning av den årliga maximala fiskeansträngningsnivån för vissa fiskevatten
med beaktande av rådets förordning (EG) nr 2027/95 av den 15 juni 1995 om en förvaltningsordning för fiskeansträngningen för vissa fiskezoner och fisketillgångar inom gemenskapen (1), särskilt artikel 4 andra strecksatsen i denna, och
Med beaktande av rådets förordning, skall följande träda i kraft omedelbart så att Nederländerna kan använda sin tilldelade kvot.
Artikel 1
Denna förordning träder i kraft dagen efter det att den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Förvaltningskommittén för nötkött har inte yttrat sig inom den tid som dess ordförande har bestämt.
1. Det pris som den behöriga myndigheten i Förenade kungariket skall betala till producenterna eller deras ombud enligt artikel 1.1 skall vara:
Ingen betalning utgår för djur vars levande vikt överskrider 560 kg, i förekommande fall beräknad genom tillämpning av koefficienterna i punkt 2.
- 1,70 när det gäller alla andra djur.
4. Om det köp som avses i artikel 1.1 avser ett kastrerat nötkreatur av hankön, skall utbetalningen av hela det pris som avses i punkt 1 endast göras om det sålda djuret inte omfattas av den ansökan om säsongsutjämningsbidrag som avses i artikel 4c i förordning (EEG) nr 805/68.
5. Den omräkningskurs som skall tillämpas är den jordbruksomräkningskurs som gäller den första dagen i den månad då djuret i fråga köps."
RÅDETS FÖRORDNING (EG) nr 2046/97 av den 13 oktober 1997 om samarbete mellan nordliga och sydliga länder i kampen mot narkotika och narkotikamissbruk
med beaktande av kommissionens förslag (1),
Snedvridningen av de sociala strukturerna i utvecklingsländerna på grund av narkotikamissbruk och den industri som är knuten till detta, skadar den hållbara sociala utvecklingen och hindrar uppnåendet av målen för gemenskapens politik inom området för utvecklingssamarbete enligt artikel 130 u i fördraget.
I sitt meddelande av den 23 juni 1994 till Europaparlamentet och rådet, lade kommissionen fram sina riktlinjer för en åtgärdsplan för Europeiska unionen som rör kampen mot narkotika (1995-1999), särskilt på internationell nivå.
Den allmänna anslutningen till konventionen ersättande äldre konventioner rörande narkotika från 1961, till samma konvention ändrad enligt protokollet från 1972, till konventionen från 1971 om psykotropa ämnen och till konventionen 1988 mot olaglig hantering av narkotika och psykotropa ämnen, liksom en systematisk tillämpning på nationell och internationell nivå av bestämmelserna i dessa fördrag, utgör hörnstenen i en internationell strategi för att bekämpa missbruk och illegal handel med narkotika.
De mänskliga rättigheterna måste respekteras när åtgärder genomförs i enlighet med denna förordning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Gemenskapen skall prioritera begäran från ett samarbetsland om att stödja utarbetandet av en nationell övergripande plan för narkotikakontroll, i nära samarbete med Förenta nationernas program för narkotikakontroll (UNDCP). Dessa planer skall fastställa mål, strategier och prioriteringar i kampen mot narkotika och därtill knutna krav på resurser (inklusive finansiella krav), för att kunna skapa ett integrerat, tvärvetenskapligt angreppssätt som spänner över flera områden och kan ge bästa möjliga effektivitet i nationella program för narkotikakontroll och internationellt bistånd.
Artikel 4
- utvecklingsländerna skall kunna genomföra "National Drug Control Master Plans", och
- Främja pilotprojekt för alternativ utveckling; genom denna process kan på lång sikt odling av illegal narkotika såväl bekämpas som elimineras genom lämpliga åtgärder för landsbygdsutveckling inom ramen för en hållbar ekonomisk tillväxt nationellt. Dessa projekt skall innefatta ekonomiska och sociala åtgärder som tar hänsyn till de faktorer som bidrar till den illegala framställningen och samtidigt åtgärder som kan underlätta ett bättre utnyttjande av handelsförmånerna. I detta sammanhang skall systematiska undersökningar genomföras om det är möjligt att ytterligare utnyttja andra finansiella gemenskapsinstrument (till exempel ALA) och Europeiska utvecklingsfonden för projekt för alternativ utveckling.
Gemenskapen ger endast stöd till projekt i vilka respekten för de mänskliga rättigheterna garanteras.
Artikel 6
3. Ekonomiska bidrag från de parter som anges i artikel 5 skall sökas för alla samarbetsåtgärder. Bidrag skall begäras inom ramen för de berörda parternas möjligheter och med hänsyn till varje åtgärds art.
6. Kommissionen skall säkerställa att gemenskapskaraktären på det bistånd som ges i enlighet med denna förordning framhävs.
b) samordning på plats av genomförandet av åtgärderna med hjälp av regelbundna möten och utbyte av information mellan kommissionens och medlemsstaternas företrädare i mottagarlandet.
Det ekonomiska stöd som ges enligt denna förordning skall vara i form av gåvobistånd.
Årliga anslag skall beviljas av budgetmyndigheten inom budgetramarna.
2. Vid bedömningen av projekt och program skall följande faktorer beaktas:
- Vilken institutionell utveckling som är nödvändig för att projektmålen skall kunna uppnås.
Kommissionen skall kortfattat informera den kommitté som avses i artikel 10 om de finansieringsbeslut som den ämnar fatta avseende projekt och program vars kostnad understiger 2 miljoner ecu. Sådan information skall lämnas senast en vecka innan beslutet fattas.
6. Om åtgärderna är föremål för finansieringsöverenskommelser mellan gemenskapen och mottagarlandet, skall i dessa föreskrivas att betalning av skatter, tullar och andra avgifter inte skall erläggas av gemenskapen.
9. Särskild uppmärksamhet skall ägnas
Artikel 10
Kommissionen skall själv anta de planerade åtgärderna om de är förenliga med kommitténs yttrande.
3. En gång om året skall en diskussion hållas på grundval av en framställning av kommissionens företrädare om de allmänna riktlinjerna för de åtgärder som skall vidtas under det kommande året inom de kommittéer som avses i punkt 1.
Sammanfattningen skall i synnerhet innehålla upplysningar om dem med vilka avtal eller kontrakt har slutits.
Artikel 12
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA BESLUT
med beaktande av rådets direktiv 94/67/EG om förbränning av farligt avfall (2), och
Den första rapporten kommer att omfatta åren från och med 1998 till och med 2000.
Artikel 1
Medlemsstaterna skall använda frågeformuläret som underlag när de utarbetar den rapport som de skall lämna till kommissionen i enlighet med artikel 5 i direktiv 91/692/EEG och artikel 17 i direktiv 94/67/EG.
KOMMISSIONENS BESLUT av den 29 juli 1998 om ändring av rådets beslut 96/411/EG om förbättring av gemenskapens jordbruksstatistik [delgivet med nr K(1998) 2135] (Text av betydelse för EES) (98/514/EG)
med beaktande av rådets beslut 96/411/EG av den 25 juni 1996 om förbättring av gemenskapens jordbruksstatistik (1), ändrat genom beslut 98/3/EG (2), särskilt artikel 8 i detta, och av följande skäl:
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för jordbruksstatistik.
Bilaga II till beslut 96/411/EG skall ersättas med bilagan till detta beslut.
RÅDETS BESLUT av den 20 juli 1998 om ingående av ett avtal om ömsesidigt erkännande mellan Europeiska gemenskapen och Kanada (98/566/EG)
med beaktande av kommissionens förslag, och
För att säkerställa att avtalet fungerar korrekt bör lämpliga interna förfaranden fastställas och det är nödvändigt att bemyndiga kommissionen att göra vissa ändringar av teknisk natur i avtalet och att fatta vissa beslut för dess genomförande.
Avtalet om ömsesidigt erkännande mellan Europeiska gemenskapen och Kanada, inbegripet dess bilagor, godkänns härmed på Europeiska gemenskapens vägnar.
Rådets ordförande skall på gemenskapens vägnar överlämna den skrivelse som avses i artikel XIX i avtalet.
2. Gemenskapens ståndpunkt vad gäller beslut som skall fattas av den gemensamma kommittén eller i förekommande fall av de gemensamma sektoriella grupperna skall, såvitt gäller ändringar i de sektoriella bilagorna (artikel XI.3 a och XI.4 i avtalet) och kontroll enligt artiklarna VIII och XI.4 c i avtalet av att gällande krav är uppfyllda, fastställas av kommissionen efter samråd med den särskilda kommitté som avses i punkt 1 i den här artikeln.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av följande: (1) Kreditförsäkringar för medellånga och långa exportaffärer spelar en viktig roll i internationell handel och utgör ett viktigt handelspolitiskt instrument.
(4) De åtgärder som föreskrivs i detta direktiv bör inte gå utöver vad som är nödvändigt för att uppnå det mål, som består i att åstadkomma den harmonisering som är nödvändig för att säkerställa att exportpolitiken grundas på enhetliga principer och att konkurrensen mellan företagen inom gemenskapen inte snedvrids.
(7) Den premie som kreditförsäkraren tar ut bör motsvara den risk som försäkras.
(10) I kommissionens vitbok om den inre marknadens fullbordande som antogs av Europeiska rådet i juni 1985 betonas vikten av ett samarbetsvänligt klimat hos gemenskapens företag.
(13) Genom beslut 93/112/EEG (3) genomförde rådet OECD-överenskommelsen om riktlinjer för exportkrediter med offentligt stöd i gemenskapsrätten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Detta direktiv är tillämpligt på försäkringsskydd för affärer avseende export av varor och/eller tjänster med ursprung i en medlemsstat, under förutsättning att detta stöd ges, direkt eller indirekt, för en eller flera medlemsstaters räkning eller med stöd av en eller flera medlemsstater och omfattar en total riskperiod på minst två år, dvs. återbetalningsperioden inklusive tillverkningsperioden.
Medlemsstaternas skyldigheter
Genomförandebeslut
Kommitté
Kommissionen skall besluta med omedelbar verkan. Om beslutet inte är förenligt med kommitténs yttrande skall kommissionen emellertid genast underrätta rådet. I sådana fall:
Artikel 5
Artikel 6
Artikel 7
Artikel 8
Ikraftträdande
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 51 och 235 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
(3) Den lagstiftning som rådet redan har antagit för att skydda rättigheterna på den sociala trygghetens område för de arbetstagare och deras familjemedlemmar som flyttar inom gemenskapen, det vill säga rådets förordningar (EEG) nr 1408/71 av den 14 juli 1971 om tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen (4) och (EEG) nr 574/72 av den 21 mars 1972 om tillämpning av förordning (EEG) nr 1408/71 om tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen (5), avser endast lagstadgade pensionssystem; det samordningssystem som föreskrivs i dessa förordningar omfattar inte kompletterande pensionssystem med undantag för system som täcks av begreppet "lagstiftning" enligt definitionen i artikel 1 j första stycket i förordning (EEG) nr 1408/71 eller med avseende på vilka en medlemsstat avger en förklaring enligt den artikeln.
(6) I sin rekommendation 92/442/EEG av den 27 juli 1992 om samstämmighet mellan mål och politik på det sociala skyddets område (6) rekommenderar rådet medlemsstaterna att "vid behov främja ändringar av villkoren för förvärv av rätt till pension, särskilt kompletterande pensionsrättigheter, för att avskaffa hindren för anställdas rörlighet".
(9) Fördraget innehåller inga andra befogenheter än de som finns i artikel 235 för att vidta lämpliga åtgärder på området social trygghet för egenföretagare.
(12) För att underlätta utövandet av rätten till fri rörlighet bör, när så behövs, nationella bestämmelser i enlighet med avdelning II i förordning (EEG) nr 1408/71 anpassas så att det blir möjligt att fortsätta att betala in avgifter till ett kompletterande pensionssystem i en medlemsstat från eller för arbetstagare som är utsända till en annan medlemsstat.
(15) Detta direktiv påverkar inte medlemsstaternas lagar ifråga om kollektiva åtgärder för att försvara yrkesintressen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Detta direktiv skall tillämpas på försäkringstagare som omfattas av kompletterande pensionssystem och andra personer som är berättigade enligt sådana system och som har förvärvat eller håller på att förvärva rättigheter i en eller flera medlemsstater.
Artikel 3
b) kompletterande pensionssystem: alla i enlighet med nationell lagstiftning och praxis inrättade tjänstepensionssystem, såsom gruppförsäkringsavtal eller system med löpande inbetalning ("pay as you go") om vilka en eller flera branscher eller sektorer kommit överens, premiereservsystem eller utfästelser om pension som garanteras av bokförda reserver, eller alla kollektiva eller andra jämförbara system vilka är avsedda som en kompletterande pension för anställda eller egenföretagare,
e) utsänd arbetstagare: en person som är utsänd till en annan medlemsstat för att arbeta och som enligt villkoren i avdelning II i förordning (EEG) nr 1408/71 fortsätter att omfattas av ursprungsmedlemsstatens lagstiftning; utsändning skall tolkas i enlighet härmed,
ÅTGÄRDER FÖR ATT SKYDDA KOMPLETTERANDE PENSIONSRÄTTIGHETER FÖR ARBETSTAGARE SOM FLYTTAR INOM GEMENSKAPEN
Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa bevarande av intjänade pensionsrättigheter för de personer, som är försäkringstagare enligt ett kompletterande pensionssystem och för vilka avgifter inte längre betalas därför att de har flyttat från en medlemsstat till en annan medlemsstat, i samma utsträckning som för de försäkringstagare för vilka avgifter inte längre betalas men som bor kvar i samma medlemsstat. Denna artikel skall också tillämpas på andra personer som är berättigade enligt bestämmelserna för det kompletterande pensionssystemet i fråga.
Medlemsstaterna skall se till att de kompletterande pensionssystemen till försäkringstagare och andra personer som är berättigade enligt dessa system i andra medlemsstater betalar ut alla förmåner som utfaller enligt dessa system, efter avdrag för de skatter och transaktionskostnader som kan vara tillämpliga.
1. Medlemsstaterna skall besluta om sådana åtgärder som behövs för att göra det möjligt att fortsätta att betala avgifter från eller för en utsänd arbetstagare som är försäkringstagare i ett kompletterande pensionssystem i en medlemsstat, under den tid som arbetstagaren är utsänd till en annan medlemsstat.
Information till försäkringstagarna
SLUTBESTÄMMELSER
Artikel 9
1. Medlemsstaterna skall sätta i kraft de lagar och författningar som är nödvändiga för att följa detta direktiv senast 36 månader efter det att direktivet har trätt i kraft eller skall säkerställa att arbetsgivare och arbetstagare senast den dagen avtalar om de bestämmelser som krävs. Medlemsstaterna är skyldiga att vidta alla de åtgärder som krävs för att de alltid skall kunna garantera de resultat som föreskrivs i detta direktiv. De skall genast underrätta kommissionen om detta.
2. Medlemsstaterna skall senast 25 januari 2002 till kommissionen överlämna texten till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 11
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
Om odlingen av potatis och tomater skyddas mot sådana skadegörare skulle produktionskapaciteten upprätthållas och dessutom skulle jordbruksproduktionen öka.
Det föreligger en avsevärd risk för odlingen av potatis och tomater i hela gemenskapen om effektiva åtgärder inte vidtas med avseende på dessa grödor för att lokalisera denna skadegörare och avgöra dess utbredning, för att förhindra dess förekomst och spridning samt, om den påträffas, för att förhindra dess spridning och bekämpa den i syfte att utrota den.
Spridningen av den sjukdomsalstrande organismen kan minskas eller förhindras genom desinfektion av sådana föremål. Varje angrepp på utsädespotatis innebär en stor risk för att den sjukdomsalstrande organismen sprids. Utsädespotatisens latenta smitta utgör på liknande sätt en stor risk för att den sjukdomsalstrande organismen sprids, och detta kan förhindras genom användning av utsädespotatis som har producerats i ett officiellt godkänt program, där utsädespotatis har testats och konstaterats vara fri från smitta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) lokalisera skadegöraren och kartlägga dess utbredning,
Artikel 2
a) på det förtecknade växtmaterialet i enlighet med de uppgifter som anges i punkt 1 i avsnitt II i bilaga I,
Ytterligare uppgifter om besiktningarna och om stickprovernas antal, ursprung och inledning samt om tidpunkten för deras insamling skall för dessa undersökningar beslutas av de ansvariga officiella organen enligt direktiv 77/93/EEG, på grundval av sunda vetenskapliga och statistiska principer och skadegörarens biologiska egenskaper samt med beaktande av de berörda medlemsstaternas särskilda produktionssystem för det förtecknade växtmaterialet och, i förekommande fall, för skadegörarens andra värdväxter.
- De lämpliga metoderna för de undersökningar och laboratorietest som avses i punkt 2 första stycket under b.
- Närmare uppgifter om de undersökningar som avses i punkt 2 andra stycket, för att säkerställa jämförbara nivåer på medlemsstaternas garantier.
Artikel 4
i) de sjukdomssymptom som orsakas av skadegöraren har diagnostiserats och ett eller flera snabbscreeningtest har genomförts med positivt resultat på sätt som anges i avsnitt I punkt 1 och avsnitt II i bilaga II, eller
c) införa lämpliga ytterligare försiktighetsåtgärder på grundval av hur stor risken bedöms vara, särskilt i förhållande till produktionen av det förtecknade växtmaterialet och flyttning av andra partier av utsädespotatis än sådana som avses under a, som har producerats på den odlingsplats där de stickprov, som avses under a, har tagits, för att hindra att skadegöraren på något sätt sprids.
- De åtgärder som anges i punkt 2 c.
a) i fråga om det förtecknade växtmaterialet vidta följande åtgärder:
iii) I enlighet med bestämmelserna i punkt 1 i bilaga V fastställa omfattningen av troliga angrepp genom kontakt före eller efter skörd, genom produktionsmässig anknytning, bevattning eller duschning eller genom klonsläktskap med det angivna angreppet.
i) Genomföra en utredning i enlighet med punkt a i.
c) I fråga om ytvatten (även flytande avfall från anläggningar för industriell bearbetning eller förpackning där det förtecknade växtmaterialet hanteras) och besläktade vilda värdväxter av familjen Solanaceae, då det har konstaterats att produktionen av det förtecknade växtmaterialet utgör en risk genom bevattning, duschning eller översvämning med ytvattnet vidta följande åtgärder:
iii) Fastställa det troliga angreppet och avgränsa ett område på grundval av förklaringen om angreppet enligt punkt ii och skadegörarens möjliga spridning med beaktande av bestämmelserna i punkt 1 och 2 ii i bilaga V.
3. Till följd av den anmälan som avses i punkt 2 och dess beståndsdelar, skall de andra medlemsstater som anges i anmälan genomföra en utredning i enlighet med punkt 1 a i och, där så är tillämpligt, punkt 1 c i och om så är lämpligt vidta ytterligare åtgärder i enlighet med punkterna 1 och 2.
2. Medlemsstaterna skall föreskriva att det förtecknade växtmaterial som förklarats troligen angripet enligt artikel 5.1 a iii och 5.1 c iii inbegripet det förtecknade växtmaterial för vilket en risk har konstaterats föreligga, och som producerats på produktionsplatser som förklarats troligen angripna enligt artikel 5.1 a iii inte får planteras och att det, under övervakning av deras ansvariga officiella organ, skall användas på lämpligt sätt eller bortförskaffas enligt punkt 2 i bilaga VI, så att det kan fastställas att det inte finns någon identifierbar risk för att skadegöraren sprids.
Artikel 7
a) i de fall då bekräftade fynd av skadegöraren har gjorts i dess egen produktion av utsädespotatis
b) i andra fall, antingen av varje planta i det ursprungliga klonurvalet eller av representativa stickprov av basutsädespotatis eller tidigare generationer.
- De bestämmelser om representativa stickprov som föreskrivs i punkt 1, andra stycket, punkt b.
Artikel 9
Artikel 11
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 21 augusti 1999. De skall genast underrätta kommissionen om detta.
Artikel 13
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 103 a.1 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
(3) Genom direktiv 73/238/EEG (5) fattade rådet beslut om lämpliga åtgärder - däribland uttag ur oljelager - som skall vidtas om det uppstår svårigheter i fråga om försörjningen av råolja och petroleumprodukter till gemenskapen. Medlemsstaterna har åtagit sig liknande skyldigheter i avtalet om ett "Internationellt energiprogram".
(6) Bestämmelserna i detta direktiv påverkar inte den fullständiga tillämpningen av fördraget, särskilt bestämmelserna om den inre marknaden och konkurrens.
(9) Lagerhållningen bör vara så organiserad att lagrens tillgänglighet och förbrukarnas tillgång till lagren säkerställs.
(12) En inhemsk utvinning bidrar i sig till försörjningssäkerhet. För medlemsstater med inhemsk oljeutvinning kan utvecklingen på oljemarknaden motivera ett lämpligt undantag från skyldigheten att hålla oljelager. I enlighet med subsidiaritetsprincipen får medlemsstaterna befria företag från skyldigheten att hålla lager i en omfattning som inte överstiger den kvantitet produkter som dessa företag framställer från råolja som utvunnits i medlemsstaten.
(15) Oljelager kan i princip hållas var som helst i gemenskapen och därför är det lämpligt att göra det enklare att upprätta lager utanför det nationella territoriets gränser. Det är nödvändigt att beslut om att hålla lager utanför det nationella territoriets gränser fattas av den berörda medlemsstatens regering i enlighet med dess behov och med hänsyn till försörjningssäkerheten. För lager som hålls tillgängliga för andra företag eller organ/enheter behövs utförligare bestämmelser för att garantera att de är tillgängliga och åtkomliga vid händelse av oljeförsörjningssvårigheter.
(18) Genom direktiv 72/425/EEG ökades den referenstid som anges i artikel 1 första stycket i direktiv 68/414/EEG från 65 till 90 dagar och villkor för genomförandet av denna utökning fastlades. Det direktivet har gjorts obsolet genom det här direktivet. Direktiv 72/425/EEG bör därför upphävas.
Artikel 1
2. Den del av den inhemska förbrukningen som täcks av petroleumprodukter baserade på utvinning inom den berörda medlemsstaten får dras av upp till högst 25 % från nämnda förbrukning. Fördelningen inom medlemsstaterna av resultatet av ett sådant avdrag skall beslutas av den berörda medlemsstaten." 2. Artikel 2 skall utgå.
"Artikel 4
I det statistiska sammandraget skall lager av jetbränsle av fotogentyp särredovisas under kategori II." 6. Artikel 5 skall ersättas med följande:
I det statistiska sammandraget av lagren som föreskrivs i artikel 4, skall färdiga produkter redovisas efter sin verkliga vikt. Råolja och halvfabrikat skall redovisas
- på grundval av förhållandet mellan den totala kvantitet som tillverkats under föregående kalenderår i den berörda staten av de produkter som omfattas av lagringsskyldigheten och den totala mängd råolja som använts under det året. Det föregående skall gälla högst 40 % av den totala lagringsskyldigheten för de första och andra kategorierna (motorbensin och tunn eldningsolja) och högst 50 % för den tredje kategorin (tjocka eldningsoljor).
"1. Vid beräkning av nivån på de minimilager som föreskrivs i artikel 1 skall endast de kvantiteter räknas in i det statistiska sammandraget som hålls i enlighet med artikel 3.1". b) Punkt 2 skall ersättas med följande:
I dessa fall skall varje medlemsstat, tillsammans med det statistiska sammandrag som föreskrivs i artikel 4, överlämna en rapport till kommissionen om de lager som hålls på medlemsstatens eget territorium till förmån för en annan medlemsstat, liksom om de lager som hålls i andra medlemsstater till dess egen förmån. I båda fallen skall rapporten innehålla uppgift om var lagren är belägna och/eller om de företag som håller lagren, lagrade kvantiteter och produktkategorier - eller uppgift om att det rör sig om råolja.
- De skall avse råolja samt alla petroleumprodukter som omfattas av detta direktiv.
- De skall normalt gälla under obegränsad tid.
- Det företag, organ eller den enhet som har rätt till lagren skall ha kontraktsenlig rätt att förvärva dessa lager under avtalsperioden. Sättet att fastställa priset för detta förvärv skall överenskommas mellan de berörda parterna.
- Den faktiska tillgången till lagren för det företag, organ/enhet som har rätt till dem måste, när som helst under avtalsperioden, garanteras av det företag, organ/enhet som håller lagren tillgängliga för det företag, organ eller den enhet som har rätt till dem.
"Artikel 6a
"Artikel 6b
Direktiv 72/425/EEG skall upphävas med verkan från och med den 31 december 1999.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 5
KOMMISSIONENS FÖRORDNING (EG) nr 121/98 av den 16 januari 1998 om ändring av bilagorna I, II och III i rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(Text av betydelse för EES)
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (1), senast ändrad genom kommissionens förordning (EG) nr 1850/97 (2), särskilt artikel 6, 7 och 8 i denna, och med beaktande av följande:
Vid fastställandet av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung är det nödvändigt att ange de djurarter i vilka restmängder kan förekomma, vilka mängder som kan förekomma i var och en av de relevanta vävnaderna från det behandlade djuret (målvävnad) samt vilket slag av restmängd som är relevant vid övervakningen av restmängder (restmarkör).
Danofloxacin, cefazolin och trimetoprim skall införas i bilaga I till förordning (EEG) nr 2377/90.
En tidsfrist på 60 dagar bör tillåtas innan denna förordning träder i kraft så att medlemsstaterna kan göra de nödvändiga anpassningarna till bestämmelserna i denna förordning av tillstånden att släppa ut de berörda veterinärmedicinska läkemedlen på marknaden, vilka beviljats enligt rådets direktiv 81/851/EEG (3), senast ändrat genom direktiv 93/40/EEG (4).
Artikel 1
Denna förordning träder i kraft den kraft den sextionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
För att säkerställa ett enhetligt genomförande av Internationella säkerhetsorganisationskoden (ISM), antog IMO genom resolution A.788 (19) av den 23 november 1995 riktlinjer om myndigheters genomförande av Internationella säkerhetsorganisationskoden (ISM-koden).
Förordning (EG) nr 3051/95 bör ändras till följd av detta.
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
Artikel 1
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
KOMMISSIONENS FÖRORDNING (EG) nr 539/98 av den 9 mars 1998 medförande ändring av förordning (EEG) nr 3077/78 om godkännande av intyg för humle som importeras från tredje land som likvärdiga med gemenskapsintyg
med beaktande av rådets förordning (EEG) nr 1696/71 av den 26 juli 1971 om den gemensamma organisationen av marknaden för humle (1), senast ändrad genom förordning (EG) nr 1554/97 (2), särskilt artikel 5.2 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I kommissionens förordning (EG) nr 2543/95 (3), ändrad genom förordning (EG) nr 2126/96 (4), föreskrivs särskilda tillämpningsföreskrifter för ordningen med exportlicenser inom olivoljesektorn. För att förbättra det sätt på vilket ordningen fungerar bör vissa särskilda tillämpningsföreskrifter fastställas för licenser utan förutfastställelse av bidraget, bl.a. vad gäller säkerhetsbeloppet och ordningen för inlämnande av ansökningar och utfärdande av licenser. Erfarenheten visar att det också är lämpligt att anpassa beloppet för säkerheten liksom tidsfristen både för inlämnandet av licensansökningar och för utfärdandet av dessa. Det är lämpligt att föreskriva att de åtgärder som vidtas när det finns risk för att de normala avsättningskvantiteterna överskrida endast får gälla exportlicenser med förutfastställelse av bidraget. För att på ett bättre sätt kunna följa exportförloppet måste de upplysningar medlemsstaterna skall lämna in preciseras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 2.2 skall "elva" ersättas med "tolv".
"3. Beloppet för säkerheten för exportlicenserna skall fastställas till
2. Följande punkt skall läggas till:
1. Punkt 1 skall ersättas med följande:
"2. Exportlicenserna med förutfastställelse av bidraget skall utfärdas första arbetsdagen från och med tisdagen den vecka som följer efter den period som avses i punkt 1, såvida inte kommissionen under tiden har vidtagit någon av de särskilda åtgärder som avses i punkt 3."
4. I artikel 3.5 sista strecksatsen skall "måndagen" ersättas med "tisdagen" och följande mening läggas till:
"6. Ansökningarna om exportlicenser utan förutfastställelse av bidraget skall lämnas in till de behöriga myndigheterna från måndag till fredag varje vecka. Licenserna skall utfärdas omedelbart."
2. Punkt 1 a skall ersättas med följande:
4. I punkt 2 skall den del av meningen som föregår den första strecksatsen ersättas med följande:
6. I punkt 2 skall följande stycke läggas till:
". . . ., och ange det regleringsår under vilket licensen utfärdades."
KOMMISSIONENS FÖRORDNING (EG) nr 1011/98 av den 14 maj 1998 om ändring av förordning (EEG) nr 1722/93 om tillämpningsföreskrifter för rådets förordningar (EEG) nr 1766/92 och (EEG) nr 1418/76 om produktionsbidrag inom spannmåls- respektive rissektorn
med beaktande av rådets förordning (EEG) nr 1766/92 av den 30 juni 1992 om den gemensamma organisationen av marknaden för spannmål (1), senast ändrad genom kommissionens förordning (EG) nr 923/96 (2), särskilt artikel 7.3 i denna,
Särskilda åtgärder kan förväntas när regleringsåret ändras, vilket innebär att såväl bidragslicensernas giltighetstid som beloppet för det enhetliga bidraget förändras.
Förvaltningskommittén för spannmål har inte yttrat sig inom den tid som dess ordförande har bestämt.
1. När ett bidrag beviljas skall det fastställas en gång i månaden. Om marknadspriserna för majs och/eller vete i gemenskapen eller på världsmarknaden varierar betydligt, får det bidrag som beräknas i enlighet med punkt 2 ändras så att hänsyn tas till sådana svängningar.
ii) genomsnittet av de representativa cif-importpriser för Rotterdam, vilket används för att beräkna importavgiften för majs och som konstaterats under de fem dagar som föregår den första tillämpningsdagen,
4. De beslut som föreskrivs i denna artikel skall fattas av kommissionen enligt förfarandet i artikel 23 i förordning (EEG) nr 1766/92."
De licenser som utfärdats efter en ansökan inlämnad under juli, augusti och fram till och med den 24 september skall dock endast vara giltiga under 30 dagar från och med den dag de utfärdas, och får inte löpa längre än till och med den 30 september.
3) I artikel 9.2 skall följande stycke läggas till:
"De köpare som per kvartal använder en kvantitet på mindre än 1 000 kg av produkterna enligt detta KN-nummer får emellertid undantas från denna bestämmelse."
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING,
För vissa beteckningar som medlemsstaterna har meddelat i enlighet med artikel 17 i förordning (EEG) nr 2018/92 har det begärts kompletterande uppgifter för att säkerställa att dessa beteckningar uppfyller kraven i artiklarna 2 och 4 i nämnda förordning. Efter granskning av dessa kompletterande uppgifter har det visat sig att dessa beteckningar stämmer överens med artiklarna i nämnda förordning. De bör därför registreras och läggas till i bilagan till kommissionens förordning (EG) nr 1107/96 (3), senast ändrad genom förordning (EG) nr 644/98 (4).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl: Bestämmelser om egenskaperna hos substrat till svampproduktion bör införas i bilaga I så att det blir möjligt att tillåta ekologisk svampproduktion i medlemsstaterna enligt samma produktionsvillkor.
I artikel 7.2 tredje strecksatsen ges möjligheten att fastställa särskilda krav på märkning av produkter som framställts med hjälp av vissa produkter som anges i bilaga II till förordning (EEG) nr 2092/91. För just denna produktionstyp är det lämpligt att för en övergångsperiod föreskriva en märkning med upplysningar om det icke-ekologiska ursprunget hos komponenterna i substratet.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som avses i artikel 14 i förordning (EEG) nr 2092/91.
Bilaga I till förordning (EEG) nr 2092/91 skall ändras i enlighet med bilagan till den här förordningen.
2. Trots vad som sägs i bestämmelserna i punkt 5.1 och 5.2 i bilaga I får medlemsstaterna under en övergångsperiod som löper ut den 1 december 2001 använda
om de produkter som anges i punkt 5.1 a och 5.2 inte kan erhållas från jordbruksföretag där en ekologisk produktionsmetod används och behovet godkänts av kontrollmyndigheten eller kontrollorganet.
RÅDETS FÖRORDNING (EG, EKSG, EURATOM) nr 2460/98 av den 12 november 1998 om ändring av förordning nr 7/66/Euratom, 122/66/EEG om fastställande av en lista över de orter för vilka transportbidrag kan beviljas, detta bidrags maximala belopp samt reglerna för dess beviljande
med beaktande av kommissionens förslag, och
Artikel 1
Artikel 2
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl: I artikel 2.1 i kommissionens förordning (EG) nr 577/97 av den 1 april 1997 om vissa tillämpningsföreskrifter för rådets förordning (EG) nr 2991/94 om regler för bredbara fetter och rådets förordning (EEG) nr 1898/87 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter (3), senast ändrad genom förordning (EG) nr 1298/98 (4), föreskrivs regler för uppgifter om totala fetthalter i bredbara fetter med undantag för de produkter som avses i förordning (EG) nr 2991/94 med en lägsta fetthalt på 80 %. I artikel 2.3 i förordning (EG) nr 577/97 och i bilaga II till den förordningen fastställs en metod för kontroll av att dessa regler iakttas. Den dag då metoden skall börja tillämpas har skjutits fram till den 1 januari 1999 för att användarna skall ha tid att inhämta erfarenheter från användningen av metoden och för att möjliggöra grundliga studier av metodens genomförbarhet med hjälp av de resultat som kommissionen fått ta del av.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
c) I alla dessa fall skall den genomsnittliga fetthalten ligga inom de gränser som fastställs i bilagan till förordning (EG) nr 2991/94."
RÅDETS FÖRORDNING (EG) nr 2531/98 av den 23 november 1998 om Europeiska centralbankens tillämpning av minimireserver
med beaktande av Europeiska centralbankens (nedan kallad ECB) rekommendation (1),
i enlighet med det förfarande som anges i artikel 106.6 i Fördraget om upprättandet av Europeiska gemenskapen (nedan kallat fördraget) samt i artikel 42 i stadgan, och på de villkor som anges i artikel 43.1 i stadgan och punkt 8 i protokoll nr 11 om vissa bestämmelser angående Förenade konungariket Storbritannien och Nordirland, och av följande skäl:
(3) Enligt artikel 19.2 i stadgan skall rådet även fastställa lämpliga sanktioner vid åsidosättande av dessa skyldigheter, och i den här förordningen fastställs specifika sanktioner. I den här förordningen hänvisas det till rådets förordning (EG) nr 2532/98 av den 23 november 1998 om Europeiska centralbankens befogenhet att förelägga sanktioner (4) när det gäller principer och förfaranden samt anges ett förenklat förfarande för sanktioner avseende vissa typer av regelöverträdelser. Om bestämmelserna i rådets förordning (EG) nr 2532/98 skulle gå emot de bestämmelser i den här förordningen som ger ECB befogenhet att förelägga sanktioner skall bestämmelserna i den här förordningen gälla.
(6) I arbetet med att fastställa detaljerade regler för åläggandet av minimireserver - inbegripet fastställandet av faktiska reservkvoter, av eventuell avkastning på reserverna, av eventuella undantag från kravet på minimireserver och av eventuella ändringar av kraven på en viss grupp eller vissa grupper av institut - måste ECB sträva efter att uppnå de mål för Europeiska centralbankssystemet (nedan kallat ECBS) som anges i artikel 105.1 i fördraget och som avspeglas i artikel 2 i stadgan. Detta innebär bland annat att ECB måste sträva efter att undvika betydande, icke önskvärda effekter i fråga om undanträngning eller disintermediering. Åläggandet av sådana krav på minimireserver kan utgöra en beståndsdel i utformningen och genomförandet av gemenskapens monetära politik, något som anges som en av ECBS:s grundläggande uppgifter i första strecksatsen i artikel 105.2 i fördraget, och som avspeglas i första strecksatsen i artikel 3.1 i stadgan.
(9) Bestämmelserna i den här förordningen kan tillämpas i sin helhet på ett verkningsfullt sätt endast om de deltagande medlemsstaterna vidtar nödvändiga åtgärder så att deras myndigheter har befogenhet att fullt ut bistå och samarbeta med ECB vad gäller insamling och kontroll av uppgifter i enlighet med vad som krävs i den här förordningen och i enlighet med artikel 5 i fördraget.
3) institut: varje enhet i en deltagande medlemsstat som ECB enligt villkoren i artikel 19.1 i stadgan kan ålägga att hålla minimireserver,
Artikel 2
Artikel 3
i) institutets skyldigheter genom mottagande av medel, tillsammans med
iv) skyldigheter gentemot ECB eller gentemot nationella centralbanker.
Artikel 4
2. Med förbehåll av punkt 1 kan ECB på icke-diskriminerande grunder fastställa skilda reservkvoter för vissa kategorier av skyldigheter som ingår i basen för minimireserverna.
När det gäller artiklarna 2, 3 och 4 skall ECB, när så är lämpligt, anta förordningar eller beslut.
1. ECB skall ha rätt att från institut inhämta de uppgifter som behövs för genomförandet av kravet på minimireserver. Sådana uppgifter skall vara insynsskyddade.
a) begära att dokument överlämnas,
d) begära skriftliga eller muntliga förklaringar.
Artikel 7
a) En räntebetalning uppgående till högst fem procentenheter över ECBS:s marginallåneränta eller två gånger ECBS:s marginallåneränta; i båda fallen skall betalningen beräknas på det belopp varmed det berörda institutets reserver understiger kravet på minimireserver.
3. Om ett institut underlåter att fullgöra skyldigheter enligt den här förordningen eller enligt ECB-förordningar eller ECB-beslut som är knutna till denna förordning, utöver de skyldigheter som avses i punkt 1, skall förordning (EG) nr 2532/98 tillämpas när det gäller sanktioner för sådan underlåtenhet och vad gäller gränser och villkor för sådana sanktioner.
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
om införande av ett enhetligt formulär för inbjudan eller åtagandeförklaring
med beaktande av artikel 132 i konventionen om tillämpning av Schengenavtalet,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Dessa skillnader ökar särskilt risken för missbruk och därför skall ett dokument införas med särskilda kännetecken till skydd mot förfalskning.
- Säkerhetsdetaljerna i dessa dokument.
2. De avtalsslutande parterna i Schengenavtalet skall fylla i det enhetliga formuläret i enlighet med bestämmelserna i den nationella lagstiftningen.
5. Frankrike skall förse Schengenstaterna med de filmer som behövs för att framställa formulären. Kostnaderna skall delas mellan de avtalsslutande parterna.
8. Detta beslut träder i kraft när de avtalsslutande parterna har meddelat att åtgärderna har genomförts. Berlin den 16 december 1998. C. H. Schapper
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Enligt artikel 13.4 krävs att det förfarande som sålunda bestämts skall anges i uppdragen och i de tekniska specifikationerna. Det är därför önskvärt att definiera de produkter eller produktgrupper som används i uppdragen och i de tekniska specifikationerna.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga byggkommittén.
För de produkter och produktgrupper som anges i bilaga I skall överensstämmelsen bestyrkas genom ett förfarande där tillverkaren ensam ansvarar för ett system för tillverkningskontroll i fabriken som säkerställer att produkten överensstämmer med de tillämpliga tekniska specifikationerna.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
om ytterligare bestämmelser för de listor över sorter av prydnadsväxter som förs av leverantörer i enlighet med rådets direktiv 98/56/EG
med beaktande av rådets direktiv 98/56/EG av den 20 juli 1998 om saluföring av förökningsmaterial av prydnadsväxter(1), särskilt artikel 9.4 i detta, och av följande skäl:
3. I enlighet med artikel 9.4 i direktiv 98/56/EG får ytterligare genomförandebestämmelser antagas för de listor över sorter av prydnadsväxter som förs av leverantör och som innehåller teknisk beskrivning och benämningar.
6. Med hänsyn till utvecklingen av gemenskapens lagstiftning om växtförädlarrätt bör det garanteras att sortbeskrivning enligt direktiv 98/56/EG överensstämmer med denna lagstiftning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
ii) Uppgifter om upprätthållande av sort och om det förökningssystem som tillämpas.
2. Punkt 1 ii och iv skall inte omfatta någon leverantör vars verksamhet inskränker sig till utsläppande på marknaden av förökningsmaterial av prydnadsväxter.
Artikel 4
3. Medlemsstaterna skall underrätta kommissionen om de viktigaste bestämmelserna i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
av den 16 december 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 137 i detta,
enligt förfarandet i artikel 251 i fördraget, och mot bakgrund av det gemensamma utkast som godkändes av förlikningskommittén den 21 oktober 1999(3), och
2. Enligt den artikeln skall dessa direktiv undvika sådana administrativa, finansiella och rättsliga ålägganden som motverkar tillkomsten och utvecklingen av små och medelstora företag.
5. Detta direktiv är ett särdirektiv i den mening som avses i artikel 16.1 i rådets direktiv 89/391/EEG av den 12 juni 1989 om åtgärder för att främja förbättringar av arbetstagarnas säkerhet och hälsa i arbetet(4). Bestämmelserna i det direktivet, särskilt de som avser information till arbetstagare, samråd och samverkan med arbetstagarna samt arbetstagares utbildning, är således också fullt tillämpliga för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär, utan att det påverkar tillämpningen av strängare eller mer detaljerade bestämmelser i det här direktivet.
8. Explosionsskydd är särskilt viktigt för säkerheten. Genom explosioner äventyras arbetstagarnas liv och säkerhet till följd av okontrollerade flammor och tryckvågor, förekomsten av hälsofarliga reaktionsprodukter och förbrukningen av den omgivande luftens syre som arbetstagarna behöver för att kunna andas.
11. Förebyggande av att explosiva atmosfärer uppstår inbegriper även tillämpning av substitutionsprincipen.
14. Rådets direktiv 92/58/EEG av den 24 juni 1992 om minimikrav beträffande varselmärkning och signaler för hälsa och säkerhet i arbetet (nionde särdirektivet enligt artikel 16.1 i direktiv 89/391/EEG)(6) är fullt tillämpligt, i synnerhet beträffande områden som omedelbart gränsar till explosionsfarliga områden, där rökning, användning av vinkelslip, svetsning och andra verksamheter som medför lågor eller gnistor kan integreras med explosionsfarliga områden.
AVDELNING I
Syfte och räckvidd
a) lokaler som används direkt för och under medicinsk behandling av patienter.
d) utvinningsindustrin som omfattas av direktiv 92/91/EEG(8) eller 92/104/EEG(9).
Artikel 2
AVDELNING II
Förebyggande av och skydd mot explosioner
- undvika att explosiv atmosfär antänds, och
Artikel 4
- sannolikheten för att explosiv atmosfär uppstår, samt dess varaktighet,
- de förväntade verkningarnas omfattning.
Artikel 5
- arbetsmiljön där explosiv atmosfär kan uppstå i sådana mängder att arbetstagares eller andras säkerhet och hälsa äventyras, arbetsmiljön är sådan att arbete kan utföras på ett säkert sätt,
Samordningsskyldighet
Artikel 7
2. Arbetsgivaren skall säkerställa att de minimikrav som fastställs i bilaga II tillämpas på områden som omfattas av punkt 1 ovan.
Explosionsskyddsdokument
- att explosionsriskerna har fastställts och bedömts,
- de områden på vilka minimikraven i bilaga II tillämpas,
Explosionsskyddsdokumentet skall ha utarbetats innan arbetet påbörjas och skall ses över när väsentliga ändringar, utvidgningar eller omvandlingar av arbetsplatsen, arbetsutrustningen eller arbetsorganisationen genomförs.
Särskilda krav för arbetsutrustning och arbetsplatser
3. Arbetsplatser med områden där explosiv atmosfär kan uppstå och som tas i bruk för första gången efter den 30 juni 2003 skall uppfylla minimikraven i detta direktiv.
AVDELNING III
Ändringar i bilagorna
- den tekniska utvecklingen, ändringar i internationella regelverk eller specifikationer samt nya rön om förebyggande av och skydd mot explosioner
Handbok för god praxis
Vid tillämpningen av detta direktiv skall medlemsstaterna i möjligast mån beakta ovannämnda handbok när de utarbetar sin nationella politik för skydd av arbetstagares hälsa och säkerhet.
Medlemsstaterna skall på begäran sträva efter att göra relevant information tillgänglig för arbetsgivare i enlighet med artikel 11, med särskild hänvisning till handboken för god praxis.
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 30 juni 2003. De skall genast underrätta kommissionen om detta.
3. Medlemsstaterna skall vart femte år till kommissionen inge en rapport om den praktiska tillämpningen av bestämmelserna i detta direktiv och i denna ange synpunkter som framförts av arbetsmarknadens parter. Kommissionen skall underrätta Europaparlamentet, rådet, Ekonomiska och sociala kommittén samt Rådgivande kommittén för arbetarskyddsfrågor därom.
av den 15 december 1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets och rådets direktiv 96/79/EG av den 16 december 1996 om skydd av förare och passagerare i motorfordon vid frontalkollision och om ändring av direktiv 70/156/EEG(3), och
2. I enlighet med artikel 4.b i direktiv 96/79/EG skall kommissionen se över och vid behov ändra tillägg 7 till bilaga II så att hänsyn tas till den provning som är avsedd för bedömning av Hybrid III-provdockans fotled, inklusive provning av fordonen.
Artikel 1
1. Från och med den 1 oktober 2000 får medlemsstaterna inte, av skäl som hänför sig till den provning som är avsedd för bedömning av Hybrid III-provdockans fotled,
om den provning som är avsedd för bedömning av Hybrid III-provdockans fotled uppfyller kraven i direktiv 96/79/EG, i dess lydelse efter ändringar genom det här direktivet.
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 30 september 2000. De skall genast underrätta kommissionen om detta.
Artikel 4
EUROPAPARLAMENTET, EUROPEISKA UNIONENS RÅD OCH EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR,
med beaktande av kommissionens beslut 1999/352/EG, EKSG, Euratom av den 28 april 1999 om inrättande av en europeisk byrå för bedrägeribekämpning(2),
(3) Det är viktigt att öka bedrägeribekämpningens omfattning och effektivitet med hjälp av de experter som finns inom området för administrativa utredningar.
(6) Dessa utredningar skall utföras på samma villkor inom alla institutioner, organ och byråer inom gemenskapen utan att överlämnandet av denna uppgift till byrån skall påverka institutionernas, organens och byråernas eget ansvar eller på något sätt minska de berörda personernas rättsliga skydd.
med uppmaning till övriga institutioner, organ och byråer att ansluta sig till detta avtal,
- bekämpa bedrägerier, korruption och all annan olaglig verksamhet som riktar sig mot Europeiska gemenskapernas ekonomiska intressen,
Utredningarna skall också utföras i enlighet med de villkor och närmare bestämmelser som avses i Europeiska gemenskapens och Europeiska atomenergigemenskapens förordningar.
4. Institutionerna skall till byrån översända de bestämmelser som de har fastställt för att genomföra detta avtal.
Detta avtal träder i kraft den 1 juni 1999.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 43 i denna,
av följande skäl: Enligt artikel 1.5 i förordning (EEG) nr 2262/84 (3) skall rådet med kvalificerad majoritet, på förslag från kommissionen, före den 1 januari 1999 fastställa formen för finansieringen av organens utgifter från och med regleringsåret 1999/2000.
Artikel 1
Kommissionen skall före den 1 oktober år 2001 undersöka om det är nödvändigt att gemenskapen fortsätter att dela organens utgifter och skall vid behov presentera ett förslag för rådet. Rådet skall, enligt förfarandet i artikel 43.2 i fördraget, före den 1 januari år 2002 besluta om eventuell finansiering av de berörda utgifterna".
KOMMISSIONENS FÖRORDNING (EG) nr 568/1999 av den 16 mars 1999 om ändring av förordning (EG) nr 577/97 om vissa tillämpningsföreskrifter för rådets förordning (EG) nr 2991/94 om regler för bredbara fetter och rådets förordning (EEG) nr 1898/87 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter
med beaktande av rådets förordning (EG) nr 2991/94 av den 5 december 1994 om regler för bredbara fetter (1), särskilt artikel 8 i denna,
KOMMISSIONENS FÖRORDNING (EG) nr 676/1999 av den 26 mars 1999 om ändring för femte gången av förordning (EG) nr 785/95 om tillämpningsföreskrifter för rådets förordning (EG) nr 603/95 om den gemensamma marknaden för torkat foder
med beaktande av rådets förordning (EG) nr 603/95 av den 21 februari 1995 om den gemensamma marknaden för torkat foder (1), senast ändrad genom förordning (EG) nr 1347/95 (2), särskilt artikel 18 i denna, och
Marknadsläget för torkat foder karakteriseras av fallande försäljningspriser och ökad produktion och är sådant att det är nödvändigt att garantera tillgången på en slutprodukt av näringsmässigt hög kvalitet framställd under likartade konkurrensvillkor och att motivera det stödbelopp som beviljas till bearbetningskostnaderna. Detta kan uppnås genom att torkning av foder vid hög temperatur tillämpas allmänt.
I vissa medlemsstater används för närvarande ett litet antal bandtorkar med en temperatur på minst 110 °C vid torkningsprocessens början. Det rör sig om små installationer med låg kapacitet vars driftstemperatur inte kan höjas utan radikala tekniska justeringar. Därför bör de omfattas av undantag från minimikravet på en torkningstemperatur på 350 °C, samtidigt som det skall stå klart att ingen ny installation av denna typ får godkännas efter det att regleringsåret 1999/2000 inletts.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 2.2 a skall den första strecksatsen ersättas med följande:
2. Medlemsstaterna skall senast den 15 maj 1999 till kommissionen översända en förteckning över de bandtorkar som godkänts före inledningen av regleringsåret 1999/2000 och som därför får omfattas av undantaget i artikel 1.1.
KOMMISSIONENS FÖRORDNING (EG) nr 730/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl: I bilaga I till förordning (EG) nr 2200/96 återfinns morötter bland de produkter för vilka normer skall antas. Kommissionens förordning (EEG) nr 920/89 av den 10 april 1989 om kvalitetsnormer för morötter, citrusfrukt, äpplen och päron(3), senast ändrad genom förordning (EG) nr 2536/98(4), har genomgått ett flertal ändringar som medför att den ur juridisk synpunkt inte längre kan anses tydlig.
Normerna skall tillämpas i samtliga handelsled. Vid transport över långa sträckor, lagring under en viss tid och olika typer av hantering kan det inträffa att produkterna försämras till följd av sin biologiska utveckling eller sin benägenhet att förfaras. Hänsyn bör därför tas till sådan försämring när normerna tillämpas i de handelsled som ligger efter avsändningstillfället. Eftersom produkter i klass "Extra" skall vara mycket noggrant sorterade och förpackade bör för dem avvikelser endast medges i fråga om bristande färskhet och saftspändhet.
Artikel 1
I de handelsled som ligger efter avsändningstillfället får dock produkterna i förhållande till de föreskrivna normerna
Artikel 2
2) Bilaga I skall utgå.
KOMMISSIONENS FÖRORDNING (EG) nr 1081/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EG) nr 3066/95 av den 22 december 1995 om vissa medgivanden i form av gemenskapstullkvoter för vissa jordbruksprodukter och om autonom anpassning under en övergångsperiod av vissa jordbrukskoncessioner som föreskrivs i Europaavtalen i syfte att beakta det jordbruksavtal som ingåtts inom ramen för de multilaterala handelsförhandlingarna under Uruguayrundan(3), senast ändrad genom förordning (EG) nr 2435/98(4), särskilt artikel 8 i denna,
(2) Garantier bör särskilt ställas för att alla berörda gemenskapsaktörer skall ges lika och fortlöpande tillträde till kvoten och för att de tullar som fatställts för dessa kvoter skall tillämpas fortlöpande på all import av djuren i fråga fram till dess att kvoten är förbrukad.
(5) För kontrollen av dessa kriterier krävs att ansökningen lämnas in i den medlemsstat där importören är registrerad i ett register för mervärdesskatt.
(8) Det bör föreskrivas att systemet skall administreras med hjälp av importlicenser. I detta syfte bör närmare bestämmelser fastställas, i synnerhet om inlämnande av ansökningar och om de uppgifter som skall lämnas i ansökningarna och i licenserna, i förekommande fall som undantag från eller tillägg till vissa bestämmelser i kommissionens förordning (EEG) nr 3719/88 av den 16 november 1988 om gemensamma tillämpningsföreskrifter för systemet med import- och exportlicenser samt förutfastställelselicenser för jordbruksprodukter(6), senast ändrad genom förordning (EG) nr 168/1999(7), och i kommissionens förordning (EG) nr 1445/95 av den 26 juni 1995 om tillämpningsföreskrifter för systemet med import- och exportlicenser för nötköttssektorn och om uphävande av förordning (EEG) nr 2377/80(8), senast ändrad genom förordning (EG) nr 2648/98(9).
(11) I artikel 7.2 och 7.3 i kommissionens förordning (EG) nr 1143/98 av den 2 juni 1998 om fastställande av tillämpningsföreskrifter för en tullkvot för kor och kvigor av vissa bergraser som inte är slaktboskap med ursprung i vissa tredje länder och om ändring av förordning (EG) nr 1012/98 föreskrivs, för att garantera efterlevnaden av bestämmelsen om att slakt av de importerade djuren inte är tillåten under en viss period, identifiering av de importerade djuren i enlighet med bestämmelserna i rådets förordning (EG) nr 820/97 av den 21 april 1997 om upprättande av ett system för identifiering och registrering av nötkreatur och om märkning av nötkött och nötköttsprodukter(14) liksom vissa ytterligare relevanta uppgifter. Eftersom dessa uppgifter redan är obligatoriska bör ovan nämnda två punkter utgå.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
>Plats för tabell>
3. Tilldelning ur tullkvoten med löpnummer 09.0003 skall beviljas på villkor att följande dokument uppvisas:
Artikel 2
Medlemsstaterna får som referenskvantiteter emellertid godkänna importtillstånd som hänför sig till föregående importår men som inte har delats ut om detta beror på ett administrativt fel som begåtts av den nationella behöriga myndigheten.
2. På grundval av ansökningarna om importtillstånd skall fördelningen av den första delen mellan de olika importörerna ske i proportion till storleken på deras import av djur enligt punkt 1 a första stycket under de 36 månader som har föregått importåret i fråga.
- skall avse minst 15 djur, och
4. Import får uteslutande bevisas med hjälp av tulldokumentet om övergång till fri omsättning som vederbörligen attesterats av tullmyndigheterna.
1. De aktörer som den 1 juni före importåret i fråga inte längre utövade någon verksamhet inom nötköttssektorn skall inte beaktas vid fördelningen i enlighet med artikel 2.1 a första stycket.
1. Ansökan om importtillstånd får endast lämnas in i den medlemsstat där den sökande är registrerad i ett nationellt register för mervärdesskatt.
3. Vid tillämpningen av artikel 2.1 a och b skall importörer senast den 15 juni före importåret i fråga för varje löpnummer lämna in ansökningar om importtillstånd till de behöriga myndigheterna, tillsammans med det bevis som anges i artikel 2.4.
- När det gäller den ordning som avses i artikel 2.1 b, en förteckning över de sökande, med uppgift om deras namn och adress samt de kvantiteter som de har ansökt om.
1. Kommissionen skall besluta om i vilken utsträckning ansökningar får godkännas.
Artikel 6
3. När kommissionen har meddelat fördelningen enligt artikel 5.1, skall importlicenserna utfärdas på begäran av den importör som erhållit importtillståndet och i dennes namn.
6. Utan att det påverkar tillämpningen av bestämmelserna i den här förordningen skall bestämmelserna i förordningarna (EEG) nr 3719/88 och (EG) nr 1445/95 tillämpas.
Artikel 7
Säkerheten skall frisläppas omedelbart om bevis har lagts fram för de berörda tullmyndigheterna att djuren
Licensansökan och licensen skall innehålla följande:
c) I fält 20, en av följande uppgifter:
1. De kvantiteter som inte omfattas av en ansökan om importlicens per den 15 mars under importåret skall omfattas av en sista fördelning för samma importår som förbehålls de berörda importörer som har ansökt om importlicens för alla de kvantiteter de har rätt till, utan att hänsyn tas till bestämmelserna i artikel 2.1 a och b.
4. En ansökan om importtillstånd från en importör som avses i punkt 1 skall gälla en kvantitet på 15 djur.
Om en sökande lämnar in mer än en ansökan för en enskild kvot skall inga ansökningar från denne för den berörda kvoten godtas.
8. Vid tillämpningen av denna artikel skall bestämmelserna i artiklarna 5-8 gälla i tillämpliga delar.
Artikel 11
2) I artikel 7 skall punkterna 2 och 3 utgå.
- Bergraser (förordning (EG) nr 1143/98), importår: ..."
KOMMISSIONENS FÖRORDNING (EG) nr 1125/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
(1) I kommissionens förordning (EG) nr 111/1999(2) fastställs allmänna tillämpningsföreskrifter för genomförande av leveranser enligt den ordning som fastställs i förordning (EG) nr 2802/98.
(4) För att göra det enklare för aktörer att delta i anbudsförfarandena förefaller det lämpligt att lätta på vissa av de ursprungliga kraven i anbudsinfordran och att ange mer detaljerade bestämmelser för hur leveranserna skall genomföras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
5) I artikel 5.1 f skall punkt 4 utgå.
14) Artikel 6.5 skall utgå.
2. Vid leverans enligt artikel 2.1 a skall interventionsorganet utfärda uttagsintyget senast tre arbetsdagar efter det att samtliga varor i ett av de magasin som anges i respektive förordning om leverans tagits ut. Interventionsorganet skall stå för de omkostnader som uppstår på grund av att uttagsintyget utfärdas för sent och dessa omkostnader skall beräknas genom tillämpning av en räntesats som skall vara samma som den räntesats som anges i bilaga VII och som är tillämplig i den berörda medlemsstaten den sista dagen för inlämning av anbud, höjd med 1 1/2 punkt."
2. Begäran om betalning för leveransen skall
- övertagandeintyg i original, i enlighet med bilaga I, utfärdat av det kontrollorgan som utsetts av kommissionen och undertecknat av den företrädare för mottagarlandet som anges i bilagan till förordningen om anbudsförfarande,
b) i de fall då artikel 2.1 a tillämpas och utöver de intyg som anges ovan i a, åtföljas av det kontrolldokument som anges i artikel 14.2.
5. Vid leverans enligt artikel 2.3 skall betalningen till den anbudsgivare som tilldelats kontrakt för anskaffande av produkter ske mot uppvisande av det uttagsintyg i enlighet med bilaga V som skall utfärdas av transportören och som skall viseras av kontrollorganet enligt artikel 9.1 efter det att hela partiet lastats.
24) I artikel 13 skall följande införas som tredje stycket: "Förskottssäkerheten skall frisläppas när villkoren för betalning av leveransen i enlighet med artikel 10 har uppfyllts."
26) Bilaga II skall ersättas med bilaga A till den här förordningen.
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om godkännande av nya fodertillsatser
med beaktande av rådets direktiv 70/524/EEG av den 23 november 1970 om fodertillsatser(1), senast ändrat genom kommissionens förordning (EG) nr 866/1999(2), särskilt artiklarna 9j och 3 i detta, och av följande skäl:
(3) I vissa medlemsstater har framgångsrika försök gjorts med en annan ny fodertillsats, "Hydratiserad kalciumaluminiumsilikat av vulkaniskt ursprung" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel". Denna nya fodertillsats bör tillåtas tillfälligt.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga foderkommittén.
"Natrolit-fonolit" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel" skall tillåtas enligt direktiv 70/524/EEG som fodertillsats E 566 på de villkor som anges i bilaga I till den här förordningen.
Artikel 3
av den 17 maj 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3),
2. Med hänsyn till att den inre marknaden innebär enhetliga prissystem och en gemensam jordbrukspolitik, bör gemenskapen stå för de ekonomiska följderna. I enlighet med denna princip, som fastställs i artikel 2.2 i förordning nr 25, bör fondens garantisektion finansiera bidrag vid export till tredje land, intervention i syfte att stabilisera jordbruksmarknader, åtgärder för landsbygdsutveckling, särskilda veterinäråtgärder enligt rådets beslut 90/424/EEG av den 26 juni 1990 om utgifter inom veterinärområdet(6), åtgärder för att informera om den gemensamma jordbrukspolitiken samt vissa utvärderingar i syfte att uppnå målen i artikel 33.1 i fördraget.
5. Ansvaret för kontrollen av garantisektionens utgifter inom fonden ligger i första hand hos medlemsstaterna, som utser myndigheter och andra organ som skall verkställa utgifter. Medlemsstaterna skall fullt ut och på ett effektivt sätt ta på sig denna uppgift. Kommissionen, som är ansvarig för att verkställa gemenskapens budget, måste kontrollera de sätt på vilka dessa utbetalningar och kontroller har utförts. Kommissionen får finansiera utgifter enbart om detta sker på ett sätt som ger tillräckliga garantier för att gemenskapsbestämmelserna efterlevs. Inom ramen för ett decentraliserat system för förvaltning av gemenskapens utgifter är det av avgörande betydelse att kommissionen, som är den institution som är ansvarig för finansieringen, är berättigad till och har möjlighet att utföra alla kontroller som den anser nödvändiga, med avseende på förvaltningen av utgifterna, samt att öppenheten och det ömsesidiga biståndet mellan medlemsstaterna och kommissionen är effektiva och fullständiga.
8. Medlemsstaterna måste tillhandahålla finansiella medel i enlighet med utbetalningsställenas behov, medan kommissionen gör förskottsutbetalningar mot utbetalningsställenas verkställda utgifter. Inom ramen för åtgärder för landsbygdsutveckling bör verkliga förskottsbetalningar göras för genomförande av program. Dessa förskottsbetalningar bör behandlas enligt de finansiella mekanismer som har upprättats för förskott mot de verkställda utgifter som har betalats under en referensperiod.
11. Åtgärder måste vidtas för att förhindra och ingripa mot oegentligheter och för att återkräva belopp som förlorats till följd av sådana oegentligheter eller sådan försumlighet. Det ekonomiska ansvaret för sådana oegentligheter eller sådan försumlighet måste fastställas.
14. Med hänsyn till omfattningen av gemenskapsfinansieringen måste Europaparlamentet och rådet regelbundet informeras genom finansiella rapporter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Utvecklingssektionen.
b) intervention i syfte att stabilisera jordbruksmarknaden,
e) åtgärder avsedda att ge information om den gemensamma jordbrukspolitiken och vissa utvärderingar av åtgärder som finansieras av fondens garantisektion.
Artikel 2
3. Om det är nödvändigt skall rådet, på förslag av kommissionen, med kvalificerad majoritet fastställa föreskrifter för finansiering av de åtgärder som avses i punkterna 1 och 2.
2. Veterinära åtgärder och växtskyddsåtgärder som vidtas enligt gemenskapsbestämmelser skall finansieras enligt artikel 1.2 d.
Artikel 4
b) Om fler än ett utbetalningsställe har ackrediterats, den myndighet eller det organ, nedan kallat "samordningsorgan", som den ger i uppdrag dels att samla in och överföra de uppgifter som skall ges in till kommissionen, dels att främja en enhetlig tillämpning av gemenskapsbestämmelserna.
b) de gjorda betalningarna redovisas korrekt och fullständigt i räkenskaperna,
4. Endast utgifter som betalas av ackrediterade utbetalningsställen skall finansieras av gemenskapen.
a) Namn och stadgar.
Kommissionen skall omedelbart underrättas om dessa uppgifter ändras på något sätt.
Artikel 5
2. Till dess att förskotten på verkställda utgifter har utbetalats skall medlemsstaterna tillhandahålla de medel som är nödvändiga för att täcka nämnda utgifter, alltefter de godkända utbetalningsställenas behov.
1. Medlemsstaterna skall med jämna mellanrum tillställa kommissionen följande uppgifter om de ackrediterade utbetalningsställena och samordningsorganen och de transaktioner som finansieras av fondens garantisektion:
2. Tillämpningsföreskrifter för denna artikel, särskilt de som gäller det redovisningsintyg som avses i punkt 1 b, skall antas enligt förfarandet i artikel 13.
2. Kommissionen skall besluta om månatliga förskott på verkställda utgifter som betalas av de ackrediterade utbetalningsställena.
3. Kommissionen skall före den 30 april året efter det aktuella budgetåret på grundval av de uppgifter som avses i artikel 6.1 b granska och godkänna räkenskaperna för utbetalningsställena.
Före varje beslut om att vägra finansiering skall resultaten av kommissionens kontroller och den berörda medlemsstatens svar överlämnas skriftligen, varefter båda parter skall söka nå en överenskommelse om vilka åtgärder som skall vidtas.
En vägran att finansiera får inte omfatta följande:
Bestämmelsen i femte stycket skall emellertid inte tillämpas på de ekonomiska följderna
5. Tillämpningsföreskrifterna för denna artikel skall antas i enlighet med förfarandet i artikel 13. Dessa föreskrifter skall särskilt omfatta de förskottsbetalningar som avses i artikel 5.1 andra stycket under punkterna 2, 3 och 4 i denna artikel och förfarandena för de beslut som avses i nämnda punkterna 2, 3 och 4.
a) försäkra sig om att transaktioner som finansieras av fonden verkligen äger rum och att de genomförs korrekt,
Medlemsstaterna skall underrätta kommissionen om de åtgärder som vidtagits i dessa syften, särskilt i vilket stadium de förvaltningsmässiga och rättsliga förfarandena befinner sig.
3. Rådet skall, på förslag av kommissionen, med kvalificerad majoritet fastställa de allmänna tillämpningsföreskrifterna för denna artikel.
Medlemsstaterna skall underrätta kommissionen om alla bestämmelser i lagar och andra författningar som de har antagit för tillämpningen av gemenskapens rättsakter avseende den gemensamma jordbrukspolitiken, i den mån dessa akter har ekonomiska följder för fonden.
a) om förvaltningsrutinerna är förenliga med gemenskapsreglerna,
Kommissionen skall i god tid före kontrollen underrätta den berörda medlemsstaten eller den medlemsstat inom vars territorium kontrollen skall äga rum. Tjänstemän från den berörda medlemsstaten får delta i kontrollen.
3. Rådet skall vid behov, på förslag av kommissionen, med kvalificerad majoritet fastställa allmänna tilllämpningsföreskrifter för denna artikel:
Artikel 11
Fondkommittén skall bestå av företrädare för medlemsstaterna och för kommissionen. Varje medlemsstat skall i fondkommittén företrädas av högst fem tjänstemän. Ordförande för fondkommittén skall vara en företrädare för kommissionen.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 205.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Medlemsstaternas röster skall vägas enligt den artikeln. Ordföranden får inte rösta.
- får kommissionen uppskjuta verkställandet av de beslutade åtgärderna under den tid som inte överstiger en månad från den dag då rådet underrättats.
1. Fondkommittén skall höras
c) om utkast till rapporter om fonden som skall överlämnas till rådet.
Artikel 15
Fondkommittén skall själv fastställa sin arbetsordning.
2. Hänvisningar till den upphävda förordningen skall tolkas som hänvisningar till denna förordning och skall läsas i enlighet med jämförelsetabellen i bilagan.
Artikel 18
Kommissionen får stryka första meningen i artikel 7.2 andra stycket enligt förfarandet i artikel 13, om de budgetmedel som beviljats fondens garantisektion och som finns tillgängliga i slutet av ett visst budgetår, gör det möjligt för fonden att finansiera de tilläggsutgifter som blir följden av strykningen för samma budgetår. Om kommissionen använder sig av denna befogenhet får den i enlighet med samma förfarande senarelägga startdatum till den 1 november för de betalningsperioder för åtgärder som påbörjas för att löpa mellan den 16 till och med den 31 oktober.
KOMMISSIONENS FÖRORDNING (EG) nr 1636/1999
med beaktande av rådets direktiv 70/524/EEG av den 23 november 1970 om fodertillsatser(1), senast ändrat genom kommissionens förordning (EG) nr 1411/1999(2), särskilt artiklarna 9j och 3 i detta, och av följande skäl:
3. Nya fodertillsatser eller nya användningsområden för fodertillsatser får ges ett provisoriskt godkännande om de vid den halt som tillåts i foder inte negativt påverkar människors eller djurs hälsa eller miljön, och inte heller skadar konsumenten genom att de förändrar animalieproduktens egenskaper, om deras förekomst i fodret kan kontrolleras, och om det är rimligt att anta - med hänsyn till tillgängliga resultat - att de har en positiv effekt på fodrets eller aminalieproduktionens egenskaper om de används i sådant foder.
6. Vetenskapliga foderkommittén har i ett yttrande fastställt att dessa preparat är ofarliga.
Artikel 1
Det preparat av typen enzymer som förtecknas i bilaga II till denna förordning får godkännas som fodertillsats i enlighet med direktiv 70/524/EEG på de villkor som anges i nämnda bilaga.
KOMMISSIONENS FÖRORDNING (EG) nr 2376/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
3. Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
3. Före den 1 april 1998 skall, särskilt enligt artikel 9i i direktiv 70/524/EEG, de preliminära godkännandena för tillsatser som avses i bilaga II och som hör till grupperna antibiotika och som förts över till bilaga B, kapitel III ersättas med godkännanden som knyts till den som är ansvarig för avyttringen.
6. De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga foderkommittén.
De preliminära godkännandena av de tillsatser som förtecknas i bilaga I till denna förordning skall ersättas med ett godkännande som knyts till den som är ansvarig för avyttringen av tillsatserna och som anges i andra kolumnen i bilaga I.
Artikel 3
av den 16 december 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
1. Förordning (EG) nr 1255/1999 ersätter, från och med den 1 januari 2000, rådets förordning (EEG) nr 804/68(2), senast ändrad genom förordning (EG) nr 1587/96(3) och, bland andra, rådets förordning (EEG) nr 987/68 av den 15 juli 1968 om fastställande av allmänna bestämmelser om beviljande av stöd för skummjölk som förädlas till kasein eller kaseinater(4), senast ändrad genom förordning (EEG) nr 1435/90(5). För att ta hänsyn till denna nya ordning bör ändringar göras av bestämmelserna i kommissionens förordning (EEG) nr 2921/90 av den 10 oktober 1990 om beviljande av stöd för framställningen av kasein och kaseinater av skummjölk(6), senast ändrad genom förordning (EG) nr 2501/1999(7). Den förordningen bör kompletteras med definitioner av de produkter som berörs av denna stödordning och det bör preciseras till vilket organ ansökan om stöd skall lämnas. Dessa bestämmelser bör gälla från och med den 1 januari 2000.
Artikel 1
b) råkasein: den produkt, olöslig i vatten, som erhålls från skummjölk genom utfällning medelst syrning med bakteriekultur eller tillsats av syra, löpe eller andra mjölkkoagulerande enzymer, utan hänsyn till eventuell föregående jonbytes- eller koncentreringsbehandling,
Artikel 2
av den 22 mars 1999
Infiltratörerna och uppgiftslämnarna bidrar med viktig hjälp i kampen mot den allvarliga brottsligheten över gränserna, i synnerhet narkotikabrottsligheten, eftersom dessa personer i allmänhet åtnjuter brottslingarnas förtroende och det med hjälp av dessa personer är möjligt att skaffa sig en allmän bild av verksamheten i de i små, enskilda enheter uppdelade brottsorganisationerna och kriminella strukturerna.
av den 21 december 1999
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
3. Hänvisningarna till lagstiftning i förlagan till sundhetsintyg i bilaga A till beslut 93/436/EEG innehåller vissa misstag och bör ändras.
Artikel 1
Detta beslut riktar sig till medlemsstaterna.
om att inte uppta monolinuron som ett verksamt ämne i bilaga I till rådets direktiv 91/414/EEG och om upphävande av tillstånd för växtskyddsmedel som innehåller detta verksamma ämne
(2000/234/EG)
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(1), senast ändrat genom kommissionens direktiv 97/73/EG(2),
(1) I kommissionens förordning (EG) nr 933/94(5), senast ändrad genom förordning (EG) nr 2230/95(6) anges verksamma ämnen i växtskyddsmedel, utses de rapporterande medlemsstaterna för genomförandet av kommissionens förordning (EEG) nr 3600/92 och fastställs anmälare för varje verksamt ämne.
(4) Kommissionen och medlemsstaterna har granskat den ingivna rapporten inom Ständiga kommittén för växtskydd. I enlighet med bestämmelserna i artikel 7.6 i förordning (EEG) nr 3600/92 slutfördes denna granskning den 20 juli 1999 genom kommissionens granskningsrapport för monolinuron.
(7) Det är därför inte möjligt att uppta detta verksamma ämne i bilaga I till direktiv 91/414/EEG.
(10) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för växtskydd.
Monolinuron skall inte tas upp som ett verksamt ämne i bilaga I till direktiv 91/414/EEG.
1. tillstånden för växtskyddsmedel som innehåller monolinuron upphävs inom en period på sex månader efter den dagen för anmälan av detta beslut,
Medlemsstaterna skall bevilja ett tidsbegränsat anstånd, under vilken tid kvarvarande lager får omhändertas, lagras, släppas ut på marknaden och användas i enlighet med artikel 4.6 i direktiv 91/414/EEG, som är så kort som möjligt och upphör inom 18 månader efter dagen för anmälan av detta beslut.
Kommissionens beslut
[delgivet med nr K(2000) 2261]
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(3) Det är därför nödvändigt att ändra den förlaga till intyg som anges i bilaga IV till direktiv 90/539/EEG samt att ändra beslut 96/482/EG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Detta beslut gäller för sändningar av dagsgamla kycklingar för vilka det utfärdas intyg från och med den 1 oktober 2000.
Kommissionens beslut
(2000/520/EG)
med beaktande av Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter(1), särskilt artikel 25.6 i detta, och
(2) Kommissionen kan konstatera att ett tredje land har en adekvat skyddsnivå. I sådana fall får personuppgifter överföras från medlemsstaterna utan att det behövs några ytterligare garantier.
(5) Den adekvata skyddsnivån för överföring av uppgifter från gemenskapen till Förenta staterna i enlighet med detta beslut bör anses ha uppnåtts om organisationer följer Safe Harbor Privacy-principerna för skydd av personuppgifter som överförs från en medlemsstat till Förenta staterna (nedan kallade principerna) och de vägledande frågorna och svaren (nedan kallade FoS) som utfärdats av Förenta staternas regering den 21 juli 2000. Organisationerna bör dessutom offentliggöra sin politik för skydd av personuppgifter och vara underställda antingen Federal Trade Commission (FTC) enligt avsnitt 5 i Federal Trade Commission Act, som förbjuder illojala eller bedrägliga handlingar eller metoder i handeln och i verksamhet som påverkar handeln, eller någon annan tillsynsmyndighet som på ett effektivt sätt ser till att principerna, tillämpade i överensstämmelse med FoS, efterlevs.
(8) För att värna om öppenhet och för att bevara förmågan hos de behöriga myndigheterna i medlemsstaterna att garantera skydd av enskilda med avseende på behandlingen av deras personuppgifter är det nödvändigt att i detta beslut specificera vilka omständigheter som i undantagsfall bör medföra att vissa dataflöden avbryts, trots att skyddsnivån befunnits vara adekvat.
(11) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som inrättats genom artikel 31 i direktiv 95/46/EG.
1. Med avseende på artikel 25.2 i direktiv 95/46/EG skall i fråga om all verksamhet som omfattas av det direktivet, safe harbor-principerna om integritetsskydd (nedan kallade principerna), se bilaga I till detta beslut, tillämpade i enlighet med den vägledning som ges i de frågor och svar (nedan kallade FoS) som utfärdats av Förenta staternas handelsministerium den 21 juli 2000, se bilaga II till detta beslut, anses utgöra en adekvat skyddsnivå för personuppgifter som överförs från gemenskapen till organisationer som är etablerade i Förenta staterna med beaktande av följande dokument som utfärdats av Förenta staternas handelsministerium:
c) En skrivelse från Federal Trade Commission, bilaga V.
a) Den organisation som tar emot uppgifterna har otvetydigt och offentligt förpliktat sig att följa principerna såsom de tillämpas i enlighet med FoS, och
Artikel 2
1. Utan att det påverkar de befogenheter behöriga myndigheter i medlemsstaterna har att vidta åtgärder för att säkra efterlevnaden av nationella bestämmelser som antagits enligt andra bestämmelser i direktiv 95/46/EG än artikel 25, får dessa myndigheter utöva sin befogenhet att tillfälligt förbjuda överföringen av uppgifter till en organisation som genom självcertifiering förbundit sig att följa principerna i överensstämmelse med FoS, i syfte att skydda enskilda med avseende på behandling av deras personuppgifter i de fall då
Förbudet skall hävas så snart det säkerställts att organisationen följer principerna i överensstämmelse med FoS och de behöriga myndigheterna i Europeiska unionen har underrättats härom.
4. Om den information som inhämtats i enlighet med punkterna 1, 2 och 3 visar att någon av de myndigheter som har ansvar för att principerna tillämpade i överensstämmelse med FoS följs i Förenta staterna inte fullgör denna uppgift på ett effektivt sätt, skall kommissionen underrätta Förenta staternas handelsministerium om detta och vid behov lägga fram förslag till bestämmelser i enlighet med det förfarande som föreskrivs i artikel 31 i direktivet i syfte att helt eller tills vidare upphäva detta beslut eller begränsa dess tillämpningsområde.
Artikel 5
Detta beslut riktar sig till medlemsstaterna.
om ett principiellt erkännande av fullständigheten hos den dokumentation som inlämnats för detaljerad granskning inför ett eventuellt införande av RH-7281 (zoxamid) och B-41; E-187 (milbemectin), BAS500F (pyraclostrobin) och AEF130360 (foramsulfuron) i bilaga I till rådets direktiv 91/414/EEG om utsläppande av växtskyddsmedel på marknaden
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) Företaget Sankyo Company Limited lämnade den 6 mars 2000 in en akt med dokumentation för det verksamma ämnet B-41; E-187 (milbemectin) till de nederländska myndigheterna.
(6) Myndigheterna i fråga underrättade kommissionen om resultaten av en första undersökning av huruvida dokumentationen var fullständig vad gäller kraven på uppgifter och upplysningar enligt bilaga II och, vad beträffar åtminstone ett växtskyddsmedel som innehåller det verksamma ämnet i fråga, enligt bilaga III till direktivet. I enlighet med artikel 6.2 överlämnade de ansökande företagen därefter akterna till kommissionen och övriga medlemsstater.
(9) En sådan bekräftelse är nödvändig för att en detaljerad granskning av dokumentationen skall kunna äga rum. Den skall också göra det möjligt för medlemsstaterna att tills vidare godkänna växtskyddsmedel som innehåller det verksamma ämnet i fråga, med beaktande av de villkor som anges i artikel 8.1 i direktivet, särskilt villkoret om att en detaljerad utvärdering av de verksamma ämnena och av växtskyddsmedlen skall göras i enlighet med direktivets bestämmelser.
(12) Förenade kungariket, Nederländerna och Tyskland skall rapportera resultaten av sina undersökningar till kommissionen, och samtidigt ge rekommendationer om huruvida införande bör beviljas eller inte, samt även ange eventuella villkor för införande senast inom ett år efter det att detta beslut har offentliggjorts.
Artikel 1
2. Den dokumentation som lämnats in av Sankyo Company Limited till kommissionen och medlemsstaterna beträffande införandet av B-41; E-187 (milbemectin) som ett verksamt ämne i bilaga I till direktiv 91/414/EEG, och som överlämnades till Ständiga kommittén för växtskydd den 31 maj 2000.
Europaparlamentets och rådets direktiv 2000/13/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(1),
(1) Rådet direktiv 79/112/EEG av den 18 december 1978 om tillnärmning av medlemsstaternas lagstiftning om märkning och presentation av livsmedel samt om reklam för livsmedel(3) har undergått flera och omfattande ändringar(4). För att skapa klarhet och av rationella skäl bör därför en kodificering företas av nämnda direktiv.
(4) Syftet med detta direktiv bör vara att anta allmänna gemenskapsregler som skall gälla horisontellt för alla livsmedel som släpps ut på marknaden.
(7) Detta behov innebär att medlemsstaterna, med hänsyn tagen till bestämmelserna i fördraget, skall kunna ställa språkliga krav.
(10) Med hänsyn till att detta direktiv är horisontellt var det från början inte möjligt att bland de obligatoriska märkningsanvisningarna ta med samtliga uppgifter som gäller för varje livsmedel och som måste framgå av den förteckning som i princip gäller för samtliga livsmedel; i ett senare steg bör gemenskapsbestämmelser antas som kompletterar de bestämmelser som redan finns.
(13) Bestämmelser måste också skapas för att ge gemenskapens lagstiftare möjlighet att, i undantagsfall, avvika från vissa förpliktelser som har fastställts generellt.
(16) Medlemsstaterna bör behålla rätten att, beroende på lokala förhållanden och praktiska omständigheter, fastställa regler för märkning av livsmedel som säljs i lös vikt; informationen bör i sådana fall likväl göras tillgänglig för konsumenten.
(19) Detta direktiv får inte påverka medlemsstaternas förpliktelser vad gäller de tidsgränser för genomförande av direktiven som anges i bilaga IV del B.
3. I detta direktiv avses med
Artikel 2
i) om vad som är utmärkande för livsmedlet, särskilt dess slag, identitet, egenskaper, sammansättning, kvantitet, hållbarhet, ursprung eller härkomst, framställnings- eller produktionsmetod,
b) såvida något annat inte följer av gemenskapsbestämmelser för naturliga mineralvatten och specialdestinerade livsmedel, tillskriva livsmedel egenskaper som förebygger, behandlar eller botar någon sjukdom hos människor eller antyda sådana egenskaper.
a) presentationen av livsmedel, särskilt med avseende på deras form, utseende eller förpackning, de förpackningsmaterial som används och det sätt på vilket livsmedlen arrangeras samt den miljö i vilken de exponeras,
1. Om något annat inte följer av artiklarna 4-17, är endast följande uppgifter obligatoriska vid märkning av livsmedel:
3. Mängden av särskilda ingredienser eller kategorier av ingredienser i enlighet med bestämmelserna i artikel 7.
6. Speciella förvarings- eller användningsanvisningar.
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt andra stycket.
10. För drycker som innehåller mer än 1,2 volymprocent alkohol, den verkliga alkoholhalten uttryckt i volym.
Artikel 4
Artikel 5
Om försäljningsnamn saknas skall det namn under vilket varan säljs vara det namn som är vedertaget i den medlemsstat i vilken den säljs till konsumenter eller institutioner och storkök, eller en beskrivning av livsmedlet och om det behövs av dess användning, vilket skall vara tillräckligt klargörande för att informera köparen om livsmedlets verkliga art och göra det möjligt för köparen att särskilja det från andra varor som det skulle kunna förväxlas med.
c) I undantagsfall får försäljningsnamnet i den medlemstat där tillverkningen sker inte användas i den medlemsstat där saluföringen sker, när den produkt som betecknas i fråga om sammansättning eller framställning skiljer sig så mycket från den produkt som är känd under det namnet att bestämmelserna i punkt b inte är tillräckliga för att säkerställa att konsumenterna i den medlemsstat där varan saluförs ges korrekt information.
Alla livsmedel som har behandlats med joniserande strålning skall förses med någon av följande uppgifter:
- på danska:
"bestrahlt" eller "mit ionisierenden Strahlen behandelt".
- på franska:
"irradiato" eller "trattato con radiazioni ionizzanti"
- på portugisiska:
"säteilytetty" eller "käsitelty ionisoivalla säteilyllä"
Artikel 6
a) - färsk frukt och färska grönsaker, inklusive potatis, som inte skalats, delats i bitar elelr behandlats på liknande sätt,
b) - ost,
förutsatt att ingen ingrediens har tillsatts utom mjölkprodukter, enzymer och kulturer av mikroorganismer som är nödvändiga för framställningen, eller det salt som behövs för framställning av annan ost än färskost och smältost,
- om ingrediensen klart framgår av försäljningsnamnet utan risk för förväxling.
b) Om en ingrediens i ett livsmedel består av flera ingredienser, skall dessa anses som ingredienser i det aktuella livsmedlet.
ii) tillsatser
iii) ämnen som används i de mängder som är absolut nödvändiga som lösningsmedel för tillsatser eller aromämnen.
Undantag:
- Ingredienserna i koncentrerade eller torkade livsmedel som är avsedda att rekonstitueras genom tillsats av vatten får anges efter proportion i den rekonstituerade varan, förutsatt att ingrediensförteckningen åtföljs av uttrycket "ingredienser i den rekonstituerade varan" eller "ingredienser i den konsumtionsfärdiga varan" eller liknande uttryck.
6. Ingredienser skall vid behov anges med sina särskilda beteckningar i enlighet med de regler som fastställts i artikel 5.
Förteckningen över kategorier i bilaga I kan ändras i enlighet med förfarandet i artikel 20.2.
Ändringar av nämnda bilaga som grundas på framsteg när det gäller vetenskapligt eller tekniskt kunnande skall antas i enlighet med förfarandet i artikel 20.2.
- De särskilda gemenskapsbestämmelserna om angivelse av behandling av en ingrediens med joniserande strålning skall antas senare i enlighet med artikel 95 i fördraget.
De gemenskapsbestämmelser som avses i denna punkt skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
a) Om den sammansatta ingrediensen utgör mindre än 25 % av den färdiga varan. Detta undantag skall dock inte gälla i fråga om tillsatser som faller under bestämmelserna i punkt 4 c.
a) om vattnet används under framställningsprocessen enbart för att rekonstituera en ingrediens som använts i koncentrerad eller torkad form,
1. Mängden av en ingrediens eller av en kategori av ingredienser som används vid tillverkningen eller beredningen av ett livsmedel skall anges i enlighet med denna artikel.
b) om den berörda ingrediensen eller kategorin av ingredienser skriftligen, genom en illustration eller grafiskt, framhävs i märkningen, eller
3. Punkt 2 skall inte tillämpas
- vars mängd, på grund av gemenskapsbestämmelser, redan måste anges i märknignen,
b) om särskilda gemenskapsbestämmelser exakt föreskriver mängden av en ingrediens eller kategori av ingredienser utan att föreskriva att detta skall anges i märkningen,
4. Den angivna mängden, uttryckt i procent, skall motsvara mängden av ingrediensen eller ingredienserna vid den tidpunkt då de användes. Gemenskapsbestämmelser får emellertid tillåta avvikelser från denna princip för vissa livsmedel. Sådanna bestämmelser skall antas i enlighet med det förfarande som anges i artikel 20.2.
Artikel 8
- i viktenheter i fråga om andra varor,
Det förfarande som fastställs i artikel 19 skall tillämpas på varje sådan nationell bestämmelse.
b) Gemenskapsbestämmelser eller, som sådana saknas, nationella bestämmelser får för vissa livsmedel, som delas in i kategorier efter mängd, innehålla föreskrifter om att mängd skall anges på annat sätt.
d) Om en fördigförpackad vara består av två eller flera separata förpackningar, som vid försäljning inte betraktas som enheter, skall nettoinnehållet anges genom uppgift om det totala nettoinnehållet och det totala antalet separata förpackningar. När det gäller vissa livsmedel behöver gemenskapsbestämmelser, eller om sådana saknas, nationella bestämmelser inte innehålla föreskrifter om att det totala antalet separata förpackningar skall anges.
Utan att det påverkar den anmälningskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt denna punkt.
Denna uppräkning kan kompletteras i enlighet med det förfarande som fastställs i artikel 20.2.
a) som minskar avsevärt i volym eller vikt och som säljs styckevis eller vägs i köparens nävraro,
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemsstaterna om varje åtgärd som vidtagits enligt denna punkt.
1. Datum för minsta hållbarhetstid för ett livsmedel skall vara den dag fram till vilken livsmedlet vid rätt förvaring har kvar sina särskilda egenskaper.
- "Bäst före..." när datumet omfattar uppgift om dagen,
- antingen själva datumet, eller
4. Datumet skall bestå av dag, månad och år i okodad kronologisk form.
- med längre hållbarhetstid än tre månader men kortare än 18 månader tillräckligt att ange månad och år,
5. Om inte annat följer av gemenskapsbestämmelser som fastställer andra typer av datummärkning, skall uppgift om hållbarhetsdatum inte krävas för:
- Drycker som innerhåller minst 10 volymprocent alkohol.
- Ättika.
- Portionsförpackningar av glass.
"sista förbrukningsdag".
- en hänvisning till var på märkningen datumet finns angivet.
4. I vissa fall kan det genom det förfarande som fastställs i artikel 20.2 avgöras huruvida villkoren i punkt 1 är uppfyllda.
2. Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser får i fråga om vissa livsmedel närmare ange hur bruksanvisningarna bör vara utformade.
Artikel 12
Artikel 13
- avsedda för konsumenter men saluförs i ett handelsled före försäljningen till konsumenten och under förutsättning att försäljning till storkök inte sker i detta handelsled,
De skall inte på något sätt döljas, skymmas eller avbrytas av annan text eller av någon illustration.
4. För regurglas som har märkning som är outplånlig och därför saknar etikett, ring eller krage samt för förpackningar eller kärl med en största yta mindre än 10 cm2, behöver endast de uppgifter anges om avss i artikel 3.1.1, 3.1.4 och 3.1.5.
De skall underrätta kommissionen om varje åtgärd som vidtagits i enlighet med punkt 5.
De får besluta att samtliga eller en del av dessa uppgifter inte behöver lämnas, förutsatt att köparen ända får tillfredsställande information.
Artikel 16
3. Bestämmelserna i punkterna 1 och 2 skall inte förhindra att uppgifterna i märkningen ges på flera språk.
Artikel 18
- skydda människors hälsa,
Artikel 19
Medlemsstaterna får vidta åtgärderna tidigast tre månader efter anmälan och under förutsättning att kommissionen inte motsatt sig det.
1. Kommissionen skall biträdas av en kommitté (nedan kallad kommittén).
3. Kommittén skall själv anta sin arbetsordning.
Artikel 22
Artikel 23
Medlemsstaterna skall se till att kommissionen får del av texten till alla väsentliga bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 26
Artikel 27
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
(1) Det är nödvändigt att fastställa renhetskriterier för alla de andra tillsatser än färgämnen och sötningsmedel som anges i Europaparlamentets och rådets direktiv 95/2/EG av den 20 februari 1995 om andra livsmedelstillsatser än färgämnen och sötningsmedel(3), senast ändrat genom direktiv 98/72/EG(4).
(4) Det är nödvändigt att beakta de specifikationer och analysmetoder för tillsatser som anges i den Codex Alimentarius som utarbetats av FAO/WHO:s gemensamma expertkommitté för livsmedelstillsatser (JECFA).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1) I bilagan skall texten avseende E 320 - butylhydroxianisol (BHA) ersättas med bilaga I till detta direktiv.
1) Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 mars 2001. De skall genast underrätta kommissionen om detta.
Artikel 3
om gränsvärden för bensen och koloxid i luften
med beaktande av kommissionens förslag(1),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) Enligt artikel 152 i fördraget skall hälsoskyddskraven ingå som ett led i gemenskapens övriga politik. I artikel 3.1 p i fördraget föreskrivs också att gemenskapens verksamhet skall bidra till att uppnå en hög hälsoskyddsnivå.
(5) Enligt direktiv 96/62/EG skall numeriska värden för gränsvärdena bygga på resultaten från det arbete som utförs av internationella forskargrupper verksamma inom området. Kommissionen bör ta hänsyn till de senaste rönen från forskning om berörda områden inom epidemiologi och miljö och de senaste framstegen inom metrologin när de faktorer som gränsvärdena bygger på tas upp till förnyad undersökning.
(8) De gränsvärden som fastställs i detta direktiv är minimikrav. I enlighet med artikel 176 i fördraget får en medlemsstat behålla eller införa strängare skyddsåtgärder. Strängare gränsvärden kan i synnerhet införas för att skydda hälsan hos särskilt sårbara kategorier av befolkningen såsom barn och patienter på sjukhus. En medlemsstat kan kräva att gränsvärdena uppnås före de datum som fastställs i detta direktiv.
(11) För att underlätta översynen av detta direktiv under år 2004 bör kommissionen och medlemsstaterna överväga att uppmuntra forskning om effekterna av bensen och koloxid. I detta sammanhang bör det förutom till utomhusluft också tas hänsyn till luftföroreningar i inomhusluft.
(14) Aktuella uppgifter om koncentrationer av bensen och koloxid i luften bör finnas lätt tillgängliga för allmänheten.
Mål
b) utvärdera koncentrationerna av bensen och koloxid i luften på grundval av gemensamma metoder och kriterier,
Artikel 2
I detta direktiv avses med
c) fasta mätningar: mätningar som utförs i enlighet med artikel 6.5 i direktiv 96/62/EG.
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att koncentrationen av bensen i luften, som utvärderats i enlighet med artikel 5, inte överskrider det gränsvärde som anges i bilaga I med hänsyn till de datum som där anges.
- fastställer de zoner och/eller den tätbebyggelse som berörs,
- anger den framtida utvecklingens huvuddrag med avseende på de åtgärder som den kommer att vidta i enlighet med artikel 8.3 i direktiv 96/62/EG.
Koloxid
Artikel 5
Minst vart femte år skall klassificeringen av varje zon eller tätbebyggelse för de syften som avses i artikel 6 i direktiv 96/62/EG ses över i enlighet med det förfarande som fastställs i avsnitt II i bilaga III till detta direktiv. Klassificeringen skall ses över tidigare om betydande ändringar ägt rum i fråga om verksamhet som påverkar koncentrationerna av bensen eller koloxid i luften.
4. För zoner och tätbebyggelser där inga mätningar krävs får modelleringsmetoder eller objektiva skattningsmetoder tillämpas.
7. De ändringar som behövs för att anpassa bestämmelserna i denna artikel samt i bilagorna III-VII till den vetenskapliga och tekniska utvecklingen skall antas i enlighet med det förfarande som avses i artikel 6.2, men de får inte leda till direkta eller indirekta ändringar av gränsvärdena.
1. Kommissionen skall biträdas av den kommitté som avses i artikel 12.2 i direktiv 96/62/EG, nedan kallad kommittén.
3. Kommittén skall själv anta sin arbetsordning.
1. Medlemsstaterna skall se till att aktuell information om koncentrationerna av bensen och koloxid i luften rutinmässigt görs tillgänglig för allmänheten, liksom för berörda organisationer, såsom miljöorganisationer, konsumentorganisationer, organisationer som företräder känsliga befolkningsgruppers intressen och andra berörda hälso- och sjukvårdsorgan, till exempel via radio och TV, tidningar, informationstavlor och datanättjänster, teletext, telefon eller fax.
2. När medlemsstaterna gör planer och program i enlighet med bestämmelserna i artikel 8.3 i direktiv 96/62/EG tillgängliga för allmänheten skall de också göra dem tillgängliga för de organisationer som avses i punkt 1 i denna artikel. Detta gäller också den dokumentation som erfordras enligt bilaga VI.II.
Rapport och översyn
a) Den nuvarande luftkvaliteten och tendenserna fram till år 2010 och därefter.
d) Nuvarande och framtida krav i fråga om information till allmänheten och utbyte av information mellan medlemsstater och kommissionen.
Artikel 9
Artikel 10
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Ikraftträdande
om fastställande av de tillämpningsföreskrifter som krävs för ett korrekt bruk av vissa bestämmelser i artikel 7 i rådets direktiv 86/362/EEG och artikel 4 i rådets direktiv 90/642/EEG om arrangemang för övervakning av gränsvärdena för bekämpningsmedelsrester i och på spannmål och produkter av vegetabiliskt ursprung inklusive frukt och grönsaker
med beaktande av rådets direktiv 86/362/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på spannmål(1), senast ändrat genom kommissionens direktiv 1999/71/EG(2), särskilt artikel 7 i detta,
(1) I artikel 7 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG fastställs grundläggande bestämmelser för kontroll av bekämpningsmedelsrester i och på spannmål respektive frukt och grönsaker.
(4) Eftersom kommissionen vid sammanställning av de uppgifter som lämnas av medlemsstaterna som underlag till de rapporter Europeiska gemenskapen skall offentliggöra måste kunna lita på uppgifternas kvalitet, noggrannhet och jämförbarhet bör kommissionen bidra ekonomiskt till åtgärder som medverkar till att kontrollprogrammen uppfyller högsta möjliga kvalitetskrav. Särskilt de regelbundna kvalifikationsprövningarna samt översynen och utformningen av riktlinjer för kvalitetskontroll i samband med regelbundna expertmöten bör stödjas.
(7) Vid de kontroller som genomfördes 1996 och 1997 påvisades överträdelser av de gränsvärden som fastställs i direktiv 90/642/EEG i dess ändrade form.
(10) De tillämpningsföreskrifter bör fastställas som krävs för ett korrekt bruk av kontrollbestämmelserna. I dessa föreskrifter bör det tydligt anges vilka åtgärder och förfaranden kommissionen får stödja ekonomiskt inom ramen för tillgängliga budgetanslag.
Artikel 1
Artikel 2
2. Inom ramen för de tillgängliga budgetanslagen i Europeiska gemenskapens budget ge ekonomiskt stöd till
c) till årlig organisation av undersökningar, samråd och andra förberedelser som krävs för att kommissionen skall kunna arbeta i riktning mot ett system som gör det möjligt att på grundval av uppgifter från kontrollprogrammen beräkna det faktiska intaget av bekämpningsmedelsrester via kosten, i enlighet med andra stycket i artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG, och
1. Kommissionen skall genom ett beslut som fattas enligt förfarandena i artikel 12 i direktiv 86/362/EEG och artikel 10 i direktiv 90/642/EEG utse den eller de mottagare av ekonomiskt stöd som avses i artikel 2.2.
- den totala kostnaden för den åtgärd som skall genomföras och åtagandena från de parter som deltar i genomförandet, inbegripet Europeiska gemenskapen,
Artikel 4
- på alla sätt har strävat efter att tillämpa de kvalitetskontroll-förfaranden för analys av bekämpningsmedelsrester som avses i artikel 2.2 b i denna förordning.
1. Kommissionen skall utse särskilda tjänstemän med lämpliga kvalifikationer för att i medlemsstaterna tillsammans med nationella myndigheter följa genomförandet av nationella respektive gemenskapens kontrollprogram för bekämpningsmedelsrester i och på livsmedel av vegetabiliskt ursprung. Detta inbegriper provtagning och kvaliteten på relevanta laboratoriers arbete.
4. Efter varje besök skall kommissionen sammanställa en skriftlig rapport. Den besökta medlemsstaten skall ges möjlighet att lämna synpunkter på rapporten.
Artikel 6
Rådets förordning (EG) nr 657/2000
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande, och
(4) För att förbättra villkoren för beslutsfattandet bör också sektorn mycket tidigt informeras om planerade initiativ, och samtliga berörda grupper bör få förklaringar till olika åtgärders syften och förutsättningar inom ramen för den gemensamma fiskeripolitiken.
Kommissionen skall, enligt de villkor som föreskrivs i bilagan, svara för utgifter avseende
Även expertmöten som kommissionen organiserar för att stödja insatser som omfattas av första stycket, andra strecksatsen, kan finansieras.
Artikel 3
av den 17 april 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 28 juli 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(3) I artikel 3 i Europaparlamentet och rådets förordning (EG) nr 1784/1999 av den 12 juli 1999 om Europeiska socialfonden(4) anges vilken typ av åtgärder som ESF kan stödja.
(6) Enligt artikel 36.1 i förordning (EG) nr 1257/1999 skall förordning (EG) nr 1260/1999 och de bestämmelser som antagits för genomförandet av den förordningen, om inte något annat följer av förordning (EG) nr 1257/1999, tillämpas på landsbygdsutvecklingsåtgärder i områden som omfattas av mål 2 som finansieras av garantisektionen inom EUGFJ. Reglerna i den här förordningen skall därför tillämpas på sådana åtgärder som omfattas av programmen för de regioner som omfattas av mål 2, såvida inte något annat följer av förordning (EG) nr 1257/1999 och kommissionens förordning (EG) nr 1750/1999(7) om tillämpningsföreskrifter till förordning (EG) nr 1257/1999.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 28 september 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175.1 i detta,
i enlighet med förfarandet i artikel 251 i fördraget(2), och
(2) Förordning (EG) nr 2037/2000 bör därför ändras.
Följande punkt skall läggas till i artikel 11.1 i förordning (EG) nr 2037/2000:
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(2) Därför bör gemensamma och harmoniserade handelsnormer fastställas för hela gemenskapsmarknaden för dessa arter genom ändring av rådets förordning (EG) nr 2406/96(3).
Förordning (EG) nr 2406/96 ändras på följande sätt:
"- Mulle (Mullus barbatus, Mullus surmuletus)
"d) Stor kammussla och andra ryggradslösa vattendjur enligt KN-nummer 0307:
2. Artikel 4.3 första stycket skall ersättas med följande text:"3. Krabba, stor kammussla och vanlig valthornssnäcka enligt artikel 3 skall inte klassificeras enligt särskilda färskhetsnormer."
4. I bilaga II skall tabellen i bilagan till den här förordningen avseende de storlekskategorier för mulle, havsruda, stor kammussla och vanlig valthornssnäcka införas efter befintlig tabell.
Europaparlamentets och rådets förordning (EG) nr 2700/2000
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
(1) I rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(4) anges det i artikel 253.4 att rådet före den 1 januari 1998 på grundval av en rapport från kommissionen, som kan åtföljas av eventuella förslag, skall se över tullkodexen för att göra nödvändiga anpassningar, med särskild hänsyn till genomförandet av den inre marknaden.
(4) De olika myndigheternas befogenheter att fastställa växelkurser efter införandet av euron har ännu inte fastställts.
(7) Det bör i enlighet med kommittéförfarandet fastställas ytterligare fall där taxeringen inom ramen för förfarandet för passiv förädling beräknas på grundval av kostnaderna för processen.
(10) I bestämmelserna om platsen för en tullskulds uppkomst bör särskilda regler införas för de fall där beloppet i fråga understiger en viss nivå.
(13) I de fall där skulden har uppkommit på grund av att en vara har undandragits från tullkontroll och där det finns fler än en gäldenär bör uppskov med betalningen av tullskulden kunna beviljas för att göra det möjligt för tullmyndigheterna att inleda ett uppbördsförfarande gentemot en bestämd gäldenär före de andra gäldenärerna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 4 skall punkt 24 ersättas med följande:
3. I artikel 77 skall den nuvarande texten betecknas punkt 1 och följande punkt skall läggas till:
"4. Åtgärder avsedda att förbjuda tillämpningen av punkt 1, att underställa tillämpningen vissa villkor eller att underlätta tillämpningen kan antas enligt kommittéförfarandet."
"Artikel 124
- importvarorna omfattas av en tullförmån inom ramen för kvotsystemet,
2. Dessutom kan ingen återbetalning av importtullar enligt restitutionssystemet ske om förädlingsprodukterna vid mottagandet av deklarationen om export omfattas av krav på uppvisande av import- eller exportintyg enligt den gemensamma jordbrukspolitiken eller om det har fastställts ett exportbidrag eller en exportavgift för dessa produkter.
"Artikel 131
9. Artikel 142 skall ersättas med följande:
2. Listan på de varor för vilka förfarandet för temporär import med partiell befrielse från importtullar inte får användas, samt de villkor under vilka förfarandet får användas, skall fastställas enligt kommittéförfarandet."
"3. Med undantag för de frizoner som utses i enlighet med artikel 168a skall frizonerna vara inhägnade. Medlemsstaterna skall fastställa infarts- och utfartsplatserna för varje frizon eller frilager."
13. Följande artikel skall införas mellan artikel 168 och punkt B (Uppläggning av varor i frizoner eller frilager):
Artiklarna 170, 176 och 180 skall inte tillämpas på de frizoner som utsetts på detta vis.
"Artikel 212a
"4. Om en tullmyndighet konstaterar att en tullskuld har uppkommit i en annan medlemsstat, i enlighet med artikel 202, skall tullskulden, om skuldbeloppet är lägre än 5000 euro, anses ha uppkommit i den medlemsstat där den konstaterades."
Om en vara erhåller förmånsbehandling på grundval av ett system för administrativt samarbete mellan tullmyndigheter som omfattar myndigheter i tredje land, skall ett ursprungsintyg som utfärdats av dessa myndigheter, om det skulle visa sig vara felaktigt, betraktas som ett misstag som inte rimligen kunde ha upptäckts på det sätt som avses i första stycket.
Gäldenären kan dock inte åberopa god tro när kommissionen i Europeiska gemenskapernas officiella tidning har offentliggjort ett yttrande om att det finns välgrundade tvivel om huruvida det land som omfattas av förmånsordningen tillämpar denna korrekt."
4. När tullskulden har uppkommit på grund av en handling som när den utfördes skulle ha kunnat ge upphov till straffrättsliga påföljder, får på de villkor som anges i de gällande bestämmelserna, underrättelsen till gäldenären lämnas efter det att treårsfristen enligt punkt 3 har löpt ut."
- när en ansökan om eftergift framställs i enlighet med artiklarna 236, 238 eller 239, eller
19. Artiklarna 247, 248 och 249 skall ersättas med följande artiklar:
Artikel 247a
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
De åtgärder som krävs för att genomföra artiklarna 11, 12 och 21 skall antas i enlighet med den förvaltningskommitté som avses i artikel 248a.2.
2. När det hänvisas till denna punkt skall artiklarna 4 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 249
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EG) nr 296/96 om de uppgifter som medlemsstaterna skall sända in för månatlig bokföring av de utgifter som finansieras genom garantisektionen vid Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) samt fastställande av vissa tillämpningsföreskrifter för rådets förordning (EG) nr 1259/1999
med beaktande av rådets förordning (EG) nr 1258/1999 av den 17 maj 1999 om finansiering av den gemensamma jordbrukspolitiken(1), särskilt artiklarna 4.8, 5.3 och 7.5 i denna, och
(2) I rådets förordning (EG) nr 974/98 av den 3 maj 1998 om införande av euron(3), ändrad genom förordning (EG) nr 2596/2000(4), föreskrivs i artikel 2 andra meningen att Greklands valuta från och med den 1 januari 2001 skall vara euron.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 3.8 b skall följande läggas till:"I Greklands fall skall regeln tillämpas fr.o.m. den 1 januari 2001."
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
om ändring av förordning (EG) nr 2125/95 om öppnande och förvaltning av tullkvoter för svampkonserver
med beaktande av rådets förordningar (EG) nr 2290/2000(1), (EG) nr 2435/2000(2) och (EG) nr 2851/2000(3) om vissa medgivanden i form av gemenskapstullkvoter för vissa jordbruksprodukter och om anpassning, som en autonom övergångsåtgärd, av vissa jordbruksmedgivanden enligt Europaavtalet med, respektive, republikerna Bulgarien, Rumänien och Polen, särskilt artikel 1.3 i dessa, och
(2) Förordning (EG) nr 3066/95 har upphävts genom förordning (EG) nr 2851/2000 och ersatts av förordningarna (EG) nr 2290/2000, (EG) nr 2435/2000 och (EG) nr 2851/2000 för respektive Bulgarien, Rumänien och Polen. Ovannämnda tullmedgivanden för svampkonserver bibehålls utan ändringar - genom förordning (EG) nr 2290/2000 och (EG) nr 2435/2000 för produkter med ursprung i Bulgarien och Rumänien, å ena sidan, och beviljas utan kvantitativa begränsningar genom förordning (EG) nr 2851/2000, för produkter med ursprung i Polen, å andra sidan. Det är därför lämpligt att ändra förordning (EG) nr 2125/95 genom att stryka alla hänvisningar till Polen, med undantag av hänvisningen till artikel 5 beträffande licensansökningar som lämnas in av traditionella importörer, för att anpassa den till dessa nya bestämmelser.
Artikel 1
Kommissionens beslut
[delgivet med nr K(2000) 3866]
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
I bilaga I till rådets direktiv 92/118/EEG skall punkt 1 a i kapitel 14 del I A ersättas med följande:
och
Detta beslut träder i kraft den 1 januari 2001.
Kommissionens beslut
[delgivet med nr K(2001) 143]
med beaktande av rådets direktiv 64/432/EEG av den 26 juni 1964 om djurhälsoproblem som påverkar handeln med nötkreatur och svin inom gemenskapen(1), senast ändrat genom direktiv 2000/20/EG(2), särskilt artikel 11.6 i detta,
med beaktande av rådets direktiv 90/426/EEG av den 26 juni 1990 om djurhälsovillkor vid förflyttning och import av hästdjur från tredje land(5), senast ändrat genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 7 i detta,
av följande skäl:
(3) Det är tillåtet att bedriva handel inom gemenskapen med embryon och ägg från arter av nötkreatur om dessa embryon och ägg har samlats in, bearbetats och lagrats av embroysamlingsgrupper som godkänts av de behöriga myndigheterna i de medlemsstater där de är verksamma.
(6) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Förteckningarna över de enheter som anges i bilaga I skall skickas till kommissionen i något av följande format: Word 97 (eller tidigare versioner), Excel 97 (eller tidigare versioner) eller pdf; filerna skall skickas till följande e-postadress: Inforvet@cec.eu.int.
Artikel 2
av den 16 januari 2001
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 2 skall ersättas med följande:
- flampunkt <= 55 °C,
- ett eller flera ämnen som klassificeras som hälsoskadliga vid en total koncentration >= 25 %,
- ett eller flera irriterande ämnen som klassificeras som R41 vid en total koncentration >= 10 %,
- ett ämne som är känt för att vara cancerframkallande (kategori 3) vid en koncentration >= 1 %,
- ett mutagent ämne (kategori 1 eller 2) som klassificeras som R46 vid en koncentration >= 0,1 %,
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
om fastställande av provtagningsplaner och diagnostiska metoder för påvisande och bekräftelse av vissa fisksjukdomar och om upphävande av beslut 92/532/EEG
(2001/183/EG)
med beaktande av rådets direktiv 91/67/EEG av den 28 januari 1991 om djurhälsovillkor för utsläppande på marknaden av djur och produkter från vattenbruk(1), senast ändrat genom direktiv 98/45/EG(2), särskilt artikel 15 i detta, och
(2) Sedan beslut 92/532/EEG fattades har både tekniska och vetenskapliga framsteg skett, och direktiv 91/67/EEG har ändrats. Detta innebär att provtagningsplaner och diagnostiska metoder måste moderniseras.
(5) De provtagningsplaner och diagnostiska metoder för påvisande och bekräftelse av vissa fisksjukdomar som infördes genom beslut 92/532/EEG måste för klarhetens skull upphävas.
Artikel 1
Detta beslut upphäver beslut 92/532/EEG.
Rådets beslut
(2001/572/EG)
med beaktande av rådets beslut 90/424/EEG av den 26 juni 1990 om utgifter inom veterinärområdet(1), särskilt artikel 24.1 och 24.2 i detta,
(1) I beslut 90/424/EEG fastställs att det är möjligt att ge finansiellt stöd från gemenskapen för bekämpning och övervakning av de sjukdomar som förtecknas i en bilaga till det beslutet.
(4) Det är viktigt att infektiös laxanemi bekämpas i syfte att förhindra dess spridning till andra områden.
(7) År 1998 kom bluetongue in på gemenskapens område från utlandet och spreds via infekterade vektorer.
(10) Med hänsyn till ovanstående bör infektiös laxanemi och bluetongue läggas till i den ovan nämnda förteckningen, så att finansiellt stöd från gemenskapen kan erhållas för genomförande av programmen för utrotning och övervakning av dessa sjukdomar. Särskilda kriterier för bluetongue bör antas för att göra det möjligt att verkställa den finansiella åtgärd som avses i artikel 24.1.
(13) Beslut 90/424/EEG bör därför ändras.
I bilagan till beslut 90/424/EEG skall följande strecksatser läggas till i Grupp 1: "- Infektiös laxanemi(5)
Detta beslut riktar sig till medlemsstaterna.
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT,
med beaktande av kommissionens förslag, och
(2) Enligt artikel 1.4 i direktiv 91/689/EEG skall medlemsstaterna till kommissionen anmäla allt avfall som inte är upptaget i förteckningen över farligt avfall, och som de anser företer någon eller några av de egenskaper som anges i bilaga 3 till direktivet. Flera medlemsstater har anmält avfall som innehåller klorsilaner, avfall som innehåller silikoner och byggmaterial som innehåller asbest och begärt att förteckning över farligt avfall skall anpassas.
(5) De åtgärder som föreskrivs i detta beslut är inte förenliga med yttrandet från den kommitté som upprättats i enlighet med artikel 18 i direktiv 75/442/EEG av den 15 juli 1975 om avfall(3). De måste därför, i enlighet med artikel 18 fjärde stycket i direktiv 75/442/EEG, antas av rådet.
Bilagan till beslut 2000/532/EG skall ändras i enlighet med bilagan till det här beslutet.
Artikel 3
av den 6 augusti 2001
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(3) Genom kommissionens beslut 93/590/EG(5), senast ändrat genom beslut 2000/112/EG(6), fastställs bestämmelser för inköp av mul- och klövsjukevirusantigen A5, A22 och O1.
(6) Genom kommissionens beslut 2000/569/EG(9), fastställs bestämmelser för inköp av ytterligare mängder av mul- och klövsjukevirusantigen A22-Iraq, O1-Manisa, ASIA 1-Shamir, A Malaysia 97, SAT 1, SAT 2 (stammar från östra respektive södra Afrika) och SAT 3.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 28 maj 2001
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA RAMBESLUT
med beaktande av Europaparlamentets yttrande(2), och
(2) Det arbete som olika internationella organisationer (t.ex. Europarådet, G8-gruppen, OECD, Interpol och FN) utför är betydelsefullt, men det behöver kompletteras med åtgärder från Europeiska unionens sida.
(5) Detta rambeslut bör bidra till kampen mot bedrägeri och förfalskning som rör andra betalningsmedel än kontanter tillsammans med andra rättsakter som rådet redan har antagit, t.ex. gemensam åtgärd 98/428/RIF(5) om inrättande av ett europeiskt rättsligt nätverk, gemensam åtgärd 98/733/RIF(6) om att göra deltagande i en kriminell organisation i Europeiska unionens medlemsstater till ett brott, gemensam åtgärd 98/699/RIF(7) om penningtvätt, identifiering, spårande, spärrande, beslag och förverkande av hjälpmedel och vinning av brott samt beslut av den 29 april 1999 om utökande av Europols mandat till att omfatta bekämpning av penningförfalskning och förfalskning av betalningsmedel(8).
(8) Det är nödvändigt att en beskrivning av de olika typer av beteenden som bör kriminaliseras i samband med bedrägeri och förfalskning som rör andra betalningsmedel än kontanter omfattar all den verksamhet som i detta avseende utgör hotet från den organiserade brottsligheten.
(11) Det är nödvändigt att medlemsstaterna ger varandra största möjliga ömsesidiga bistånd och samråder med varandra när fler än en medlemsstat är behöriga i fråga om samma brott.
Definitioner
b) juridisk person: varje enhet som har denna ställning enligt tillämplig lagstiftning, med undantag av stater eller andra offentliga organ vid utövandet av de befogenheter som de har i egenskap av statsmakter samt internationella offentliga organisationer.
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att följande handlingar är straffbara när de är uppsåtliga, åtminstone när det gäller kreditkort, eurocheckkort, andra kort utgivna av finansinstitut, resecheckar, eurocheckar, andra checkar och växlar:
c) Mottagande, förskaffande, transport, försäljning eller överlämnande till en annan person eller innehav av ett betalningsinstrument som stulits eller olovligen tillgripits eller som är helt eller delvis förfalskat med syfte att använda det för bedrägeri.
Datorrelaterade brott
- att utan rätt ingripa i ett dataprograms eller datasystems funktion.
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att följande handlingar är straffbara när de är uppsåtliga:
- datorprogram som är avsedda för att begå något av de brott som avses i artikel 3.
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att deltagande i och anstiftan till sådana handlingar som avses i artiklarna 2-4 eller försök till sådana handlingar som avses i artikel 2 a, 2 b, 2 d och artikel 3 är straffbara.
Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att de handlingar som avses i artiklarna 2-5 är belagda med straffrättsliga påföljder som är effektiva, proportionella och avskräckande och som, åtminstone i allvarliga fall, omfattar påföljder som är frihetsberövande och kan medföra utlämning.
1. Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att juridiska personer kan ställas till ansvar för sådana handlingar som avses i artikel 2 b-d och artiklarna 3-4 och som till deras förmån begås av varje person som agerar antingen enskilt eller som en del av den juridiska personens organisation och har en ledande ställning inom den juridiska personen, grundad på
- befogenhet att utöva kontroll inom den juridiska personen,
3. Den juridiska personens ansvar enligt punkterna 1 och 2 utesluter inte lagföring av fysiska personer som är gärningsmän, anstiftare eller medhjälpare till de handlingar som avses i artikel 2 b-d och artiklarna 3-4.
1. Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att en juridisk person som har ställts till ansvar i enlighet med artikel 7.1 kan bli föremål för effektiva, proportionella och avskräckande påföljder, som skall innefatta bötesstraff eller administrativa avgifter och som kan innefatta andra påföljder, t.ex.
c) rättslig övervakning,
Artikel 9
a) helt eller delvis på medlemsstatens territorium,
2. Om inte annat följer av artikel 10, kan en medlemsstat besluta att inte tillämpa behörighetsregeln eller att endast i särskilda fall eller under särskilda omständigheter tillämpa regeln i
3. Medlemsstaterna skall vederbörligen underrätta rådets generalsekretariat om de beslutar att tillämpa punkt 2, om så är lämpligt med angivande av de särskilda fall eller omständigheter då beslutet gäller.
1. a) Varje medlemsstat som enligt sin lag inte utlämnar sina egna medborgare skall vidta nödvändiga åtgärder för att fastställa sin behörighet rörande brott enligt artiklarna 2, 3, 4 och 5 när de begås av en av dess egna medborgare utanför dess territorium.
Artikel 11
2. Om flera medlemsstater är behöriga i fråga om brott som avses i detta rambeslut skall dessa stater samråda med varandra i syfte att samordna sina insatser för en effektiv lagföring.
1. Medlemsstaterna skall antingen utse operativa kontaktpunkter eller också kan de använda befintliga operativa strukturer för informationsutbyte samt för annan kontakt mellan medlemsstaterna för att tillämpa detta rambeslut.
Territoriell tillämpning
Genomförande
Artikel 15
Europaparlamentets och rådets direktiv 2001/108/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
(1) Räckvidden av rådets direktiv 85/611/EEG(4) var ursprungligen begränsad till sådana företag för kollektiva investeringar av den öppna typen som utbjuder sina andelar till allmänheten inom gemenskapen och som har som enda syfte att investera i överlåtbara värdepapper (fondföretag). I ingressen till direktiv 85/611/EEG såg man framför sig att sådana företag för kollektiva investeringar som inte omfattades av direktivet skulle kunna bli föremål för samordning i ett senare skede.
(4) Penningmarknadsinstrument omfattar de kategorier av överlåtbara instrument som normalt inte handlas på reglerade marknader utan som omsätts på penningmarknaden, till exempel statsskuldväxlar, kommunala skuldväxlar, bankcertifikat, företagscertifikat, omsättningsbara medelfristiga skuldväxlar och bankaccepter.
(7) Utvecklingen av möjligheterna för ett fondföretag att investera i fondföretag och i andra företag för kollektiva investeringar bör underlättas. Det är därför väsentligt att se till att en sådan investeringsverksamhet inte minskar skyddet för investerarna. På grund av fondföretagens ökade möjligheter att investera i andelar i andra fondföretag och/eller företag för kollektiva investeringar är det nödvändigt att fastställa vissa regler om kvantitativa begränsningar, tillhandahållande av information och förhindrande av uppkomsten av s.k. kaskadfonder.
(10) Av försiktighetsskäl är det nödvändigt att fondföretag, när det gäller investeringar som utsätter dem för en motpartsrisk, undviker orimlig koncentration till samma organ eller till organ som tillhör samma grupp.
(13) Derivattransaktioner får aldrig användas för att kringgå principerna och reglerna i detta direktiv. För OTC-derivat måste det finnas ytterligare regler för riskspridningen som bör tillämpas vid exponering i förhållande till en enda motpart eller grupp av motparter.
(16) Det finns ett behov av att säkerställa fri saluföring över gränserna av andelar i ett större urval av företag för kollektiva investeringar, samtidigt som en enhetlig miniminivå för skydd av investerare tillhandahålls. De uppsatta målen kan därför endast nås genom att de överenskomna miniminormerna fastställs i ett bindande gemenskapsdirektiv. Detta direktiv gäller endast den erforderliga minimiharmoniseringen och går i enlighet med artikel 5 tredje stycket i fördraget inte utöver vad som är nödvändigt för att uppnå dessa mål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 1.2 första strecksatsen skall ersättas med följande: "- som har till enda syfte att företa kollektiva investeringar i överlåtbara värdepapper och/eller i andra likvida finansiella tillgångar som avses i artikel 19.1 med kapital från allmänheten och som tillämpar principen om riskspridning, och"
- obligationer eller andra skuldförbindelser (nedan kallade skuldförbindelser),
9. I detta direktiv avses med 'penningmarknadsinstrument' instrument som normalt omsätts på penningmarknaden och som är likvida och har ett värde som vid varje tidpunkt exakt kan fastställas."
5. Artikel 19.1 skall ändras på följande sätt:
- dessa andra företag för kollektiva investeringar är auktoriserade enligt lagstiftning som fastställer att de är föremål för tillsyn som av de behöriga myndigheterna med ansvar för fondföretaget anses motsvara den tillsyn som fastställs i gemenskapslagstiftningen och att det anses tillräckligt säkerställt att samarbete mellan myndigheterna sker, och
- de fondföretag eller andra företag för kollektiva investeringar i vars andelar förvärv planeras, enligt dessas fondbestämmelser eller bolagsordning, får investera högst 10 % av sina tillgångar i andelar i andra fondföretag eller andra företag för kollektiva investeringar, och/eller
- de underliggande tillgångarna utgörs av sådana instrument som avses i denna punkt 1, finansiella index, räntesatser, växelkurser eller utländska valutor, i vilka fondföretaget kan investera utifrån de investeringsmål som det har angett i sina fondbestämmelser eller sin bolagsordning,
h) andra penningmarknadsinstrument än de som omsätts på en reglerad marknad och som faller under artikel 1.9, om själva emissionen eller emittenten av instrumenten reglerats i syfte att skydda investerare och sparmedel och under förutsättning att de har
- emitterats eller garanterats antingen av en inrättning som är föremål för tillsyn i enlighet med de kriterier som fastställs i gemenskapslagstiftningen eller av en inrättning som omfattas av och följer sådana tillsynsregler som av de behöriga myndigheterna anses minst lika stränga som de som fastställs i gemenskapslagstiftningen, eller
7. Artikel 19.2 b och 19.3 skall utgå.
1. Förvaltnings- eller investeringsbolaget måste använda ett förfarande för riskhantering som gör det möjligt för det att vid varje tidpunkt kontrollera och bedöma den risk som är knuten till positionerna och deras bidrag till portföljens allmänna riskprofil; bolaget måste använda ett förfarande som möjliggör en exakt och oberoende bedömning av värdet på OTC-derivat. Bolaget måste underrätta de behöriga myndigheterna regelbundet och i enlighet med de detaljerade regler de skall fastställa om de typer av derivatinstrument, underliggande risker, kvantitativa begränsningar liksom de metoder som valts för att beräkna de risker som åtföljer transaktioner med derivatinstrument för varje fondföretag som det förvaltar.
3. Ett fondföretag skall säkerställa att dess totala exponering som hänför sig till derivatinstrument inte överskrider dess portföljs totala nettovärde.
När ett överlåtbart värdepapper eller ett penningmarknadsinstrument innefattar ett derivat måste detta beaktas när kraven i denna artikel skall uppfyllas.
1. Ett fondföretag får investera högst 5 % av sina tillgångar i överlåtbara värdepapper eller penningmarknadsinstrument som emitterats av samma organ. Ett fondföretag får investera högst 20 % av sina tillgångar i inlåning i samma organ.
- 5 % av fondföretagets tillgångar i andra fall.
- investeringar i överlåtbara värdepapper eller penningmarknadsinstrument som emitterats av,
Om ett fondföretag investerar mer än 5 % av sina fondtillgångar i sådana obligationer som avses i första stycket och som har samma emittent, får det totala värdet av dessa investeringar inte överstiga 80 % av värdet av fondföretagets tillgångar.
De gränser som anges i punkterna 1, 2, 3 och 4 får inte kombineras, och investeringar i överlåtbara värdepapper och penningmarknadsinstrument emitterade av samma organ eller i inlåning eller derivatinstrument från detta organ enligt bestämmelserna i punkterna 1, 2, 3 och 4 får därför under inga förhållanden överstiga sammanlagt 35 % av ett fondföretags tillgångar.
11. Följande artikel skall läggas till: "Artikel 22a
- Indexet skall utgöra en lämplig referens för den marknad det hänför sig till.
12. I artikel 23.1 skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
2. Investeringar i andelar i företag för kollektiva investeringar som ej är fondföretag får sammanlagt inte överstiga 30 % av fondföretagets tillgångar.
Ett fondföretag som investerar en betydande del av sina tillgångar i andra fondföretag och/eller företag för kollektiva investeringar, skall i sitt prospekt uppge maximinivån för de förvaltningskostnader som kan debiteras både fondföretaget självt och de andra fondföretag och/eller företag för kollektiva investeringar i vilka fondföretaget ämnar investera. Fondföretaget skall i sin årsrapport ange en maximal procentsats för de förvaltningskostnader som debiteras både fondföretaget självt och de fondföretag och/eller företag för kollektiva investeringar i vilka det investerar."
2. När ett fondföretag huvudsakligen investerar i någon annan kategori av de tillgångar som anges i artikel 19 än överlåtbara värdepapper och penningmarknadsinstrument eller efterbildar aktieindex eller index för skuldebrev enligt artikel 22a måste dess prospekt och i förekommande fall allt övrigt reklammaterial ange investeringspolicyn på framträdande plats.
15. Artikel 25.2 skall ändras enligt följande:
16. Andra meningen i artikel 25.2 skall ersättas med följande: "De gränsvärden som anges i andra, tredje och fjärde strecksatserna behöver inte iakttas vid förvärvstillfället, om bruttomängden av skuldförbindelserna eller av penningmarknadsinstrumenten eller nettomängden av de värdepapper som är föremål för emission då inte kan beräknas."
19. Artikel 26.1 skall ersättas med följande: "1. Fondföretag behöver inte iaktta de gränsvärden som anges i detta avsnitt när de nyttjar teckningsrätter för överlåtbara värdepapper eller penningmarknadsinstrument som ingår i fondtillgångarna.
22. Efter artikel 53 skall följande artikel läggas till: "Artikel 53a
- Likriktning av definitionerna i fråga om terminologi och utformning i enlighet med senare rättsakter avseende fondföretag och närstående frågor.
3. Kommittén skall själv anta sin arbetsordning.".
a) en analys av hur man kan fördjupa och vidga den inre marknaden för fondföretag, särskilt vad gäller gränsöverskridande marknadsföring av fondföretag (även tredjemansfonder), hur passet för förvaltningsföretag fungerar, hur det förenklade prospektet fungerar som informations- och marknadsföringsverktyg, en översyn av omfattningen av tillhörande verksamhet samt möjligheterna till förbättrat samarbete mellan kontrollmyndigheter vad gäller enhetlig tolkning och tillämpning av direktivet,
d) en översyn av investeringsbestämmelserna för fondföretag, till exempel användningen av derivatinstrument och andra instrument samt tekniker för värdepapper, reglering av indexfonder, reglering av penningmarknadsinstrument, inlåning, reglering av fond-till-fond-investeringar liksom de olika investeringsgränserna,
2. Medlemsstaterna får bevilja fondföretag, som är verksamma vid tidpunkten för detta direktivs ikraftträdande, en frist om högst 60 månader från denna tidpunkt för att de skall kunna anpassa sig till den nya nationella lagstiftningen.
De skall börja tillämpa dessa åtgärder senast den 13 februari 2004.
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 70/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
efter att ha offentliggjort ett utkast till denna förordning(2),
(1) Genom förordning (EG) nr 994/98 bemyndigas kommissionen att i enlighet med artikel 87 i fördraget förklara att stöd till små och medelstora företag på vissa villkor skall vara förenliga med den gemensamma marknaden och undantagna från anmälningsskyldigheten enligt artikel 88.3 i fördraget.
(4) Denna förordning påverkar inte medlemsstaternas möjligheter att anmäla stöd till små och medelstora företag. Sådana anmälningar kommer att bedömas av kommissionen särskilt utifrån kriterierna i denna förordning. Riktlinjerna för statligt stöd till små och medelstora företag bör upphävas den dag då denna förordning träder i kraft, eftersom deras innehåll förs in i den här förordningen.
(7) Denna förordning bör inte påverka tillämpningen av särskilda regler i förordningar och direktiv om statligt stöd inom vissa sektorer, såsom de gällande reglerna för varvssektorn, och den bör inte vara tillämplig inom jordbruks- samt fiske- och vattenbrukssektorn.
(10) För att fastställa huruvida stöd som omfattas av denna förordning är förenliga med den gemensamma marknaden, är det nödvändigt att ta hänsyn till stödnivån och således stödbeloppet uttryckt i bidragsekvivalenter. Vid beräkningen av bidragsekvivalenten av stöd som kan betalas ut i flera omgångar och stöd i form av mjuka lån måste de marknadsräntor som rådde när stödet beviljades användas. För att säkerställa en enhetlig, öppen och enkel tillämpning av reglerna för statligt stöd, bör med marknadsräntor i denna förordning avses referensräntorna, under förutsättning att det ställs normala säkerheter när det gäller mjuka lån och att dessa inte innebär ett onormalt risktagande. Referensräntorna bör vara de räntor som löpande fastställs av kommissionen på grundval av objektiva kriterier och som offentliggörs i Europeiska gemenskapernas officiella tidning samt på Internet.
(13) Det är lämpligt att fastställa ytterligare villkor som bör uppfyllas av varje stödordning eller enskilt stöd som beviljas undantag med stöd av denna förordning. Med hänvisning till artikel 87.3 c i fördraget bör sådana stöd normalt inte ha som enda syfte att fortlöpande eller periodiskt minska de driftskostnader som stödmottagaren normalt skall stå för, och de bör stå i proportion till de hinder som måste övervinnas för att uppnå de sociala och ekonomiska fördelar som anses vara i gemenskapens intresse. Tillämpningsområdet för denna förordning bör därför begränsas till stöd som ges till vissa materiella och immateriella investeringar, vissa tjänster som tillhandahålls stödmottagarna och viss övrig verksamhet. Mot bakgrund av den överkapacitet inom transportsektorn som råder i gemenskapen, med undantag för rullande järnvägsmateriel, bör transportmedel och transportutrustning inte ingå i de stödberättigande investeringskostnaderna för företag som har sin huvudsakliga ekonomiska verksamhet inom transportsektorn.
(16) Mot bakgrund av Världshandelsorganisationens (WTO) avtal om subventioner och kompensatoriska åtgärder(7) bör exportstöd och stöd som gynnar inhemska produkter på bekostnad av importerade produkter inte undantas enligt denna förordning. Bidrag till kostnaderna för deltagande i handelsmässor eller för undersökningar eller konsulttjänster som behövs för att lansera en ny produkt eller en befintlig produkt på en ny marknad utgör normalt inte exportstöd.
(19) Undantag bör enligt denna förordning inte medges stöd som kumuleras med annat statligt stöd, inbegripet stöd från nationella, regionala eller lokala myndigheter, eller med gemenskapsbidrag, om, i förhållande till samma stödberättigande kostnader, ett sådant kumulerat stöd, överstiger de tröskelvärden som anges i denna förordning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Denna förordning gäller för statligt stöd som beviljas små och medelstora företag inom alla sektorer, utan att det påverkar tillämpningen av särskilda gemenskapsförordningar eller gemenskapsdirektiv enligt EG-fördraget vilka styr beviljandet av statligt stöd till särskilda sektorer, oavsett om de är mer eller mindre restriktiva än denna förordning.
b) exportrelaterade stöd, d.v.s. stöd som är direkt knutna till exporterade volymer, till upprättandet eller driften av ett distributionsnät eller till andra löpande uppgifter som har samband med exportverksamhet,
Definitioner
b) små och medelstora företag: företag som definieras i bilaga I.
e) stödnivå brutto: stödbeloppet uttryckt i procent av projektets stödberättigande kostnader. Alla siffror som används skall avse belopp före eventuella avdrag för direkt skatt. Om stöd beviljas i någon annan form än som bidrag, skall stödbeloppet vara lika med stödets bidragsekvivalent. Stöd som betalas ut i flera omgångar skall aktualiseras till sitt värde vid tidpunkten för beviljandet. Den ränta som skall användas för nuvärdesberäkningar och för att räkna ut stödbeloppet i ett mjukt lån skall vara den gällande referensräntan vid den tidpunkt då lånet beviljades.
Artikel 3
2. Stödordningar som uppfyller samtliga villkor enligt denna förordning skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget, under förutsättning att
3. Stöd som beviljas enligt en sådan stödordning som avses i punkt 2 skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget, under förutsättning att det beviljade stödet direkt uppfyller samtliga villkor i denna förordning.
1. Stöd till investeringar i materiella och immateriella tillgångar inom och utom gemenskapen skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskraven i artikel 88.3 i fördraget om det uppfyller villkoren i punkterna 2-6.
b) 7,5 % för medelstora företag.
b) 15 procentenheter brutto i de områden som omfattas av artikel 87.3 a, under förutsättning att den totala stödnivån netto inte överstiger 75 %.
5. Om stödet beräknas på grundval av investeringskostnaderna, skall de stödberättigande kostnaderna för materiella investeringar utgöra kostnader som avser investeringar i mark, byggnader, maskiner och utrustning. Inom transportsektorn får, med undantag för rullande järnvägsmateriel, transportmedel och transportutrustning inte ingå i de stödberättigande kostnaderna. Stödberättigande kostnader för immateriella investeringar skall vara kostnader för förvärv av teknologi.
b) Investeringsprojektet måste leda till en nettoökning av antalet sysselsatta i den berörda anläggningen i förhållande till det genomsnittliga antalet anställda under de senaste tolv månaderna.
Rådgivningsverksamhet och andra tjänster och verksamheter
b) För deltagande i mässor och utställningar får stödet brutto inte överstiga 50 % av merkostnaderna för hyra, uppförande och drift av utställningsmontern. Detta undantag skall endast gälla för ett företags första deltagande i en viss mässa eller utställning.
Ett enskilt stöd som uppfyller ett av följande tröskelvärden får inte beviljas undantag enligt denna förordning:
ii) stödnivån netto i områden som är berättigade till regionalstöd är minst 50 % av stödtaket netto enligt regionalstödskartan för området i fråga, eller
Villkor för stödet
- har antagit bestämmelser som fastställer en laglig rätt till stöd enligt objektiva kriterier och utan vidare diskretionär prövningsrätt för medlemsstaten
1. De stödtak som fastställs i artiklarna 4, 5 och 6 skall tillämpas oavsett om stödet helt finansieras med statliga medel eller samfinansieras av gemenskapen.
Insyn och kontroll
3. Medlemsstaterna skall sammanställa en rapport om tillämpningen av denna förordning för varje helt kalenderår eller del av kalenderår under vilket denna förordning gäller, enligt den förlaga som anges i bilaga III och även i elektronisk form. Medlemsstaterna skall överlämna en sådan rapport till kommissionen senast tre månader efter utgången av den period som rapporten avser.
1. Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EG) nr 562/2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 1254/1999 vad avser systemen för offentliga interventionsuppköp inom nötköttssektorn och förordning (EG) nr 2734/2000
med beaktande av rådets förordning (EG) nr 1254/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för nötkött(1), särskilt artikel 47.8 i denna, och
(2) Med hänsyn till den exceptionella situationen på marknaden och för att de interventionsåtgärder som föreskrivs i förordning (EG) nr 2734/2000 skall ha större effekt bör det medges undantag från artikel 4.2 g i förordning (EG) nr 562/2000 vad gäller den maximala vikten för slaktkroppar genom att inte fastställa någon viktbegränsning för de två anbudsförfarandena under februari månad och genom att öka vikten till 430 kg för de resterande anbudsförfarandena under det första kvartalet 2001 och samtidigt tillåta uppköp av tyngre djur, men då begränsa priset för dessa till det pris som betalas för den högsta tillåtna vikten.
(5) I bilaga III till förordning (EG) nr 562/2000 fastställs de bestämmelser som hela och halva slaktkroppar samt kvartsparter måste följa om de skall få köpas upp för offentlig intervention. För att anpassa bestämmelserna till gällande handelssed bör beskrivningen av halva slaktkroppar i den bilagan ändras så att den tillåter viss variation.
(8) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för nötkött.
Artikel 6.1 i förordning (EG) nr 2734/2000 skall ersättas med följande:
- får slaktkroppar med en vikt över 430 kg köpas för intervention vid de resterande anbudsförfarandena under det första kvartalet 2001, men i sådana fall skall uppköpspriset högst vara det som betalas för den maximala vikten."
1. Artikel 4.3 d skall ersättas med följande:
"b) halv slaktkropp: de produkter som erhålls genom symmetrisk delning av den slaktkropp som avses i a ovan genom mitten av hals-, rygg-, länd- och korskotorna och genom mitten av bröstbenet och bäckenbensfogen. Under uppslaktning och hantering av slaktkroppen får inte rygg- och ländkotorna tydligt förskjutas. Tillhörande muskler och senor får inte skadas allvarligt av såg eller kniv."
Kommissionens förordning (EG) nr 749/2001
(Text av betydelse för EES)
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), senast ändrad genom kommissionens förordning (EG) nr 2908/2000(2), särskilt artiklarna 7 och 8 i denna, och
(2) Gränsvärden bör fastställas först efter det att Kommittén för veterinärmedicinska läkemedel har granskat all relevant information beträffande säkerheten med restmängder av ämnet i fråga för den som konsumerar livsmedel med animaliskt ursprung samt restmängdernas påverkan på den industriella bearbetningen av livsmedel.
(5) För veterinärmedicinska läkemedel som är avsedda för äggläggande fåglar, mjölkdjur eller honungsbin, måste gränsvärden även fastställas för ägg, mjölk eller honung.
(8) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
Bilaga II till förordning (EEG) nr 2377/90 skall ändras i enlighet med bilagan till den här förordningen.
Kommissionens förordning (EG) nr 939/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) I artikel 6.1 i rådets förordning (EG) nr 2406/96 av den 26 november 1996 om fastställande av gemensamma marknadsnormer för saluföring av vissa fiskeriprodukter(7), senast ändrad genom förordning (EG) nr 2578/2000(8), föreskrivs att produkter i kategori B inte skall berättiga till ekonomiskt stöd i samband med intervention inom ramen för den gemensamma organisationen av marknaden. I den mån som endast produkter av kvalitet Extra, "E" och "A" berättigar till schablonmässigt stöd enligt artikel 24 i förordning (EG) nr 104/2000, bör beräkningen av stödberättigande kvantiteter uteslutande göras på grundval av dessa produktkategorier.
(6) För beräkningen av det schablonmässiga stödet bör medlemsstaterna tillåtas att fastställa ett schablonvärde, fördelat på de återtagna produkternas avsättning enligt kommissionens förordning (EEG) nr 1501/83 av den 9 juni 1983 om omhändertagande av vissa fiskeriprodukter som varit föremål för marknadsstabiliserande åtgärder(9), ändrad genom förordning (EEG) nr 1106/90(10).
(9) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fiskeriprodukter.
Allmänna villkor
Det schablonmässiga stödet skall betalas ut till den berörda producentorganisationen först sedan medlemsstatens behöriga myndighet har konstaterat att de kvantiteter för vilka stödet har sökts inte överstiger den högsta nivå som anges i artikel 24.5 i förordning (EG) nr 104/2000.
Artikel 3
Medlemsstaterna skall fastställa ett schablonvärde för att beräkna schablonersättning och tillhörande förskott, fördelat på de återtagna produkternas avsättning enligt artikel 1 b, c och d i förordning (EEG) nr 1501/83.
Villkor för att bevilja schablonmässigt stöd enligt artikel 24.4 i förordning (EG) nr 104/2000 (nedan kallat schablonbidrag)
2. Schablonbidraget skall beräknas på grundval av de faktiska tekniska och ekonomiska kostnader för nödvändiga åtgärder vid stabiliseringsbehandling och lagring av produkterna i fråga som noterats i gemenskapen under det föregående fiskeåret.
b) Arbetskostnader i samband med lagring och uttag från lager.
e) Transportkostnader från landningsställe till plats där beredningen sker.
Artikel 6
Schablonbidraget skall betalas ut till den berörda producentorganisationen först sedan medlemsstatens behöriga myndighet har konstaterat att de kvantiteter för vilka bidraget har sökts antingen beretts och lagrats eller konserverats och sedan återförts till marknaden i enlighet med bestämmelserna i artikel 4 i förordning (EG) nr 2814/2000.
Artikel 8
3. Förskotten skall fastställas på grundval av det under perioden rådande preliminära förhållandet mellan återtagna och saluförda kvantiteter. Beräkningen av beloppet skall justeras två månader efter den aktuella månaden på grundval av de transaktioner som faktiskt genomförts och skall redovisas enligt den förlaga som finns i bilagan.
1. Medlemsstaterna skall införa en ordning för att kontrollera att den information som lämnas i ansökningarna om utbetalning överensstämmer med de kvantiteter som producentorganisationen i fråga faktiskt har salufört och återtagit från marknaden.
Artikel 10
Förordning (EEG) nr 4176/88 skall upphöra att gälla.
av den 22 maj 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 152.4 b i detta,
efter att ha hört Regionkommittén,
(1) Flera olika typer av transmissibel spongiform encefalopati (TSE) har sedan flera år tillbaka konstaterats oberoende av varandra hos människor och djur. Bovin spongiform encefalopati (BSE) upptäcktes först hos nötkreatur 1986 och under följande år också hos andra djurarter. En ny variant av Creutzfeldt-Jakobs sjukdom (CJS) beskrevs 1996. Det samlas ständigt nya bevis för likheten mellan BSE-smittämnet och det smittämne som förorsakar den nya varianten av Creutzfeldt-Jakobs sjukdom.
(4) Kommissionen har erhållit vetenskapliga yttranden om flera aspekter av TSE, bland annat från Vetenskapliga styrkommittén och Vetenskapliga kommittén för veterinära åtgärder till skydd för människors hälsa. Vissa av dessa yttranden avser åtgärder för att minska den potentiella risken för att människor och djur skall utsättas för produkter från infekterade djur.
(7) Ett förfarande bör fastställas för att bestämma den epidemiologiska statusen för en medlemsstat, ett tredje land och en av dess regioner (nedan kallade länder eller regioner) med hänsyn till BSE på grundval av en bedömning av risken för förekomst (på engelska: incident risk), spridning och risk för att människor utsätts för smitta, utifrån tillgänglig information. Medlemsstater och tredje land som väljer att inte ansöka om att få sin status fastställd bör av kommissionen placeras i en kategori, på grundval av all information som kommissionen har tillgång till.
(10) Vissa vävnader från idisslare bör betecknas som specificerat riskmaterial på grundval av de olika TSE-typernas patogener och den epidemiologiska statusen för det land eller den region där det berörda djuret har sitt ursprung eller sin hemvist. De specificerade riskmaterialen måste avlägsnas och destrueras på ett sådant sätt att människor och djur inte utsätts för några hälsorisker. Framför allt bör de inte avyttras för att användas vid tillverkning av livsmedel, foder eller gödningsmedel. Bestämmelser bör emellertid införas om möjlighet att uppnå en likvärdig hälsoskyddsnivå, med hjälp av ett TSE-test som utförs på enskilda djur, sedan full validitet fastställts. Slakttekniker som innebär en risk för att material från hjärnan infekterar andra vävnader bör inte tillåtas i andra länder eller regioner än de där BSE-risken är lägst.
(13) Om förekomst av TSE bekräftas officiellt, bör den behöriga myndigheten vidta alla nödvändiga åtgärder, i synnerhet låta destruera slaktkroppen, och genomföra en undersökning för att identifiera alla riskdjur och fastställa restriktioner för förflyttning av djur och animaliska produkter för vilka smittorisk konstaterats. Ägarna bör utan dröjsmål ersättas för förlust av djur och animaliska produkter som destruerats enligt denna förordning.
(16) Avyttring av vissa animaliska produkter som härrör från nötkreatur i högriskregioner bör förbjudas. Detta förbud bör dock inte gälla vissa animaliska produkter som framställs under kontrollerade förhållanden och som kommer från djur för vilka det kan fastställas att de inte utgör någon hög risk för infektion med TSE.
(19) Handelsåtgärderna när det gäller TSE bör bygga på internationella standarder, riktlinjer eller rekommendationer, om sådana finns. Åtgärder som är vetenskapligt underbyggda och som säkerställer ett bättre sanitärt skydd får dock vidtas om de åtgärder som är grundade på relevanta internationella standarder, riktlinjer eller rekommendationer inte skulle säkerställa ett lämpligt hälsoskydd.
(22) De åtgärder som krävs för att genomföra denna förordning bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(4).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
2. Denna förordning skall inte tillämpas på
c) animaliska produkter som är avsedda för utställning, undervisning, forskning, specialstudier eller analyser, förutsatt att de inte slutligen kan konsumeras eller användas av människor eller andra djur än de som används för de aktuella forskningsprojekten,
Separering av levande djur och animaliska produkter
Artikel 3
a) TSE: samtliga former av transmissibel spongiform encefalopati utom de som människor kan drabbas av.
d) utgångsmaterial: råvaror eller andra animaliska produkter från vilka eller med vars hjälp de produkter som avses i artikel 1.2 a och 1.2 b framställs.
g) specificerat riskmaterial: de vävnader som specificeras i bilaga V. Om inte annat anges, skall produkter som innehåller eller härrör från dessa vävnader inte inbegripas i denna definition.
j) provtagning: provtagning, med statistiskt korrekt underlag, från djur eller deras omgivning eller från animaliska produkter för att ställa en sjukdomsdiagnos eller fastställa släktskap, övervaka hälsan samt kontrollera frånvaron av mikrobiologiska agenser eller vissa material i animaliska produkter.
m) alternativt test: de test som avses i artikel 8.2 och som används i stället för avlägsnande av specificerat riskmaterial.
Artikel 4
2. Skyddsåtgärderna skall antas i enlighet med det förfarande som avses i artikel 24.2 och Europaparlamentet skall samtidigt underrättas om dessa åtgärder och om motiveringen till dem.
Artikel 5
Medlemsstaterna och de tredje länder som vill stå kvar på förteckningarna över tredje länder som är godkända för att till gemenskapen exportera de levande djur eller de produkter som avses i denna förordning, skall till kommissionen lämna en ansökan om fastställande av deras BSE-status, tillsammans med relevanta uppgifter avseende kriterierna i kapitel A i bilaga II och de potentiella riskfaktorerna i kapitel B i bilaga II samt deras utveckling över tiden.
Efter det att Internationella byrån för epizootiska sjukdomar har fastställt ett förfarande för klassificering av länder i kategorier och om den har placerat det ansökande landet i någon av dessa kategorier, får det beslutas om en förnyad bedömning av den gemenskapskategorisering som genomförts för det berörda landet i enlighet med första stycket i denna punkt, i förekommande fall i enlighet med det förfarande som avses i artikel 24.2.
Snabbtest skall godkännas för detta ändamål enligt det förfarande som avses i artikel 24.2 och införas i en förteckning i kapitel C.4 i bilaga X.
4. De medlemsstater eller tredje länder som inte lämnat in någon ansökan enligt punkt 1 inom sex månader från och med den 1 juli 2001 skall, när det gäller export från deras territorier av levande djur eller animaliska produkter, betraktas som länder i kategori 5 enligt kapitel C i bilaga II så länge de inte har lämnat in någon ansökan.
För att tredje land skall få exportera levande djur eller animaliska produkter för vilka det finns särskilda bestämmelser i denna förordning till gemenskapen enligt de villkor som grundar sig på den kategori som kommissionen fastställt, skall de förbinda sig att utan dröjsmål till kommissionen skriftligen anmäla alla epidemiologiska eller andra bevis som skulle kunna leda till ändringar i deras BSE-status.
KAPITEL III
Övervakningssystem
2. Medlemsstaterna skall underrätta kommissionen och de övriga medlemsstaterna i Ständiga veterinärkommittén om uppkomst av annan TSE än BSE.
Artikel 7
2. Dessutom skall det förbud som avses i punkt 1 även gälla djur och animaliska produkter i enlighet med punkt 1 i bilaga IV.
Tredje land eller regioner i tredje land som har placerats i kategori 5 skall inte tillåtas att till gemenskapen exportera sådant foder för livsmedelsproducerande djur som innehåller protein som härrör från däggdjur eller foder som är avsett för däggdjur, med undantag av hundar och katter, och som innehåller bearbetat protein som härrör från däggdjur.
Specificerat riskmaterial
2. Punkt 1 skall inte tillämpas på vävnader från djur som har genomgått ett alternativt test som godkänts för detta särskilda syfte i enlighet med det förfarande som avses i artikel 24.2 och som införts i förteckningen i kapitel C.5 i bilaga X och tillämpas enligt de villkor som anges i punkt 5 i bilaga V, och där testresultaten är negativa.
4. De uppgifter om ålder som anges i bilaga V skall anpassas regelbundet. Denna anpassning skall genomföras på grundval av de senaste säkra vetenskapliga rönen om den statistiska sannolikheten för att TSE förekommer inom de berörda åldersgrupperna av gemenskapens bestånd av nötkreatur, får och getter.
6. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
1. De animaliska produkter som räknas upp i bilaga VI får inte framställas av material som härrör från idisslare från länder eller regioner som är placerade i kategori 5, såvida de inte framställs i enlighet med de produktionsprocesser som har godkänts i enlighet med det förfarande som avses i artikel 24.2.
4. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
1. Medlemsstaterna skall se till att personalen vid den behöriga myndigheten, diagnostiska laboratorier samt utbildningsanstalter för lantbruk och veterinärmedicin, officiella veterinärer, praktiserande veterinärer, slakteripersonal samt personer som föder upp, håller och hanterar djur får utbildning när det gäller kliniska tecken, epidemiologi samt, när det gäller personal som har ansvar för inspektionerna, utbildning i att tolka laboratorieresultat som rör TSE.
KONTROLL OCH UTROTNING AV TSE
Utan att det påverkar tillämpningen av direktiv 82/894/EEG(12) skall medlemsstaterna se till att alla djur som misstänks vara smittade med TSE omedelbart anmälas till de behöriga myndigheterna.
Artikel 12
Om man misstänker BSE hos ett nötkreatur på en anläggning i en medlemsstat, skall alla övriga nötkreatur på denna anläggning vara föremål för officiella restriktioner vad avser förflyttning i avvaktan på att resultaten av undersökningen blir tillgängliga.
En medlemsstat får, enligt det förfarande som avses i artikel 24.2 och med avvikelse från kraven i andra, tredje och fjärde styckena i denna punkt, undantas från tillämpning av officiella restriktioner vad avser förflyttning av djur, om medlemsstaten tillämpar åtgärder som erbjuder likvärdiga garantier.
4. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
1. Om förekomst av TSE har bekräftats officiellt, skall följande åtgärder vidtas utan dröjsmål:
c) Alla djur och animaliska produkter som avses i punkt 2 i bilaga VII och som vid den undersökning som avses i punkt b har konstaterats vara riskdjur, skall avlivas och destrueras fullständigt i enlighet med punkterna 3 och 4 i bilaga V.
Om det kan styrkas att anläggningen där det smittade djuret befann sig när TSE bekräftades förmodligen inte är den anläggning där djuret exponerats för TSE, får den behöriga myndigheten besluta att båda anläggningarna eller bara den anläggning där djuret exponerats skall placeras under officiell övervakning.
5. Utan att det påverkar tillämpningen av direktiv 82/894/EEG skall varje bekräftat fall av en annan typ av TSE än BSE anmälas till kommissionen på årlig basis.
Beredskapsplan
KAPITEL V
Levande djur, deras sperma, embryon och ägg
3. Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
1. Följande animaliska produkter från friska idisslare skall inte vara föremål för restriktioner när de avyttras eller i förekommande fall exporteras enligt denna artikel och enligt bestämmelserna i kapitlen C och D i bilaga VIII och i kapitlen A, C, F och G i bilaga IX:
ii) Mjölk avsedd för framställning av mjölkbaserade produkter enligt definitionen i direktiv 92/46/EEG.
v) Hudar och skinn i den mening som avses i direktiv 92/118/EEG(14).
2. Animaliska produkter från tredje land som har placerats i kategorierna 2, 3, 4 och 5 skall härröra från nötkreatur, får och getter som inte har utsatts för sådan laceration av vävnad från centrala nervsystemet som anges i artikel 8.3, eller avlivats med gas som har injicerats i hjärnskålen.
b) djur som är födda, har fötts upp och hållits i besättningar som bevisligen varit BSE-fria sedan minst 7 år tillbaka i tiden.
5. De animaliska produkter för vilka det anges särskilda regler i denna artikel skall åtföljas av sådana lämpliga hälsointyg eller handelsdokument som föreskrivs i gemenskapslagstiftningen i enlighet med artiklarna 17 och 18 eller, om det inte finns något sådant krav i gemenskapslagstiftningen, av ett hälsointyg eller ett handelsdokument, för vilka modeller skall fastställas i enlighet med det förfarande som avses i artikel 24.2.
Artikel 17
Artikel 18
REFERENSLABORATORIER, PROVTAGNING, UNDERSÖKNINGAR OCH KONTROLLER
1. De nationella referenslaboratorierna i varje medlemsstat samt deras behörighet och uppgifter fastställs i kapitel A i bilaga X.
Provtagning och metoder för laboratorieanalyser
Artikel 21
Tillämpningsföreskrifter för denna artikel, särskilt sådana som syftar till att reglera formerna för samarbete med de nationella myndigheterna, skall fastställas enligt det förfarande som avses i artikel 24.2.
ÖVERGÅNGSBESTÄMMELSER OCH SLUTBESTÄMMELSER
1. Bestämmelserna i del A i bilaga XI skall tillämpas under en period på minst sex månader räknat från den 1 juli 2001; denna period upphör samma dag som ett beslut har antagits i enlighet med bestämmelserna i artikel 5.2 eller 5.4; från och med den dagen skall artikel 8 tillämpas.
4. De minimikriterier som denna statistiska undersökning skall uppfylla fastställs i del B i bilaga XI.
Efter samråd med den relevanta vetenskapliga kommittén om sådana frågor som kan ha konsekvenser för folkhälsan skall bilagorna ändras eller kompletteras och lämpliga övergångsbestämmelser antas, i enlighet med det förfarande som avses i artikel 24.2.
Kommittéer
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader, och när det gäller skyddsåtgärder enligt artikel 4.2 i denna förordning skall tiden vara 15 dagar.
Samråd med vetenskapliga kommittéer
Ikraftträdande
av den 28 juni 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I artikel 18 i förordning (EG) nr 1493/1999 föreskrivs att producenter av druvor avsedda för vinframställning och producenter av druvmust och vin varje år skall deklarera vilka mängder som producerats av den senaste skörden, samt att både producenter av druvmust och vin och andra näringsidkare än detaljhandlare varje år skall deklarera sina lager av druvmust och vin.
(4) Det är inte nödvändigt att kräva två deklarationer från producenter som kan lämna alla nödvändiga uppgifter i produktionsdeklarationen. Småproducenter kan undantas från deklarationsskyldighet eftersom deras sammanlagda produktion utgör en relativt blygsam andel av produktionen inom gemenskapen.
(7) Uppgifterna om vinarealerna kan vara oriktiga på grund av att deklaranten inte har haft de kontrollmöjligheter som krävs. I sådana fall bör påföljden stå i proportion till hur grava felen är i den inlämnade deklarationen.
(10) Enligt rådets förordning (EEG) nr 2392/86(3), senast ändrad genom förordning (EG) nr 1631/98(4), skall ett gemenskapsregister över vinodlingar upprättas. De medlemsstater som förfogar över ett fullständigt register bör tillåtas att använda vissa uppgifter ur registret om de inte finns i deklarationen.
(13) För att uppnå nödvändig överensstämmelse mellan de påföljder som föreskrivs i denna förordning och påföljderna enligt kommissionens förordning (EG) nr 1623/2000(5), senast ändrad genom förordning (EG) nr 545/2001(6), är det lämpligt att ändra sistnämnda förordning och införa en lämplig formulering om påföljderna.
Artikel 1
1. Fysiska eller juridiska personer eller sammanslutningar av sådana personer som odlar druvor, nedan kallade skördare, skall varje år till de behöriga myndigheter som har utsetts av medlemsstaterna överlämna en skördedeklaration till den administrativa enhet som fastställs. Skördedeklarationen skall minst innehålla de uppgifter som framgår av tabell A och, i förekommande fall, tabell B i bilagan.
a) Skördare vars hela produktion av druvor är avsedd för konsumtion i färskt tillstånd, för torkning eller för omedelbar bearbetning till druvsaft.
i) vinodlarens förnamn, efternamn och adress,
I det sista fallet skall vinkooperativet eller sammanslutningen kontrollera att uppgifterna i deklarationen stämmer med de uppgifter som kooperativet har.
b) Skördare som är anslutna till eller tillhör ett vinkooperativ eller en sammanslutning och som levererar hela sin skörd, i form av vin eller druvmust, till detta vinkooperativ eller denna sammanslutning, inklusive sådana skördare som avses i artikel 4.4.
1. Fysiska eller juridiska personer eller sammanslutningar av sådana personer, inbegripet vinkooperativ, som av innevarande vinårs skörd har framställt vin och/eller vid de tidpunkter som anges i artikel 11.1 innehar andra produkter än vin, skall varje år till de behöriga myndigheter som har utsetts av medlemsstaterna överlämna en produktionsdeklaration som innehåller minst de uppgifter som skall anges enligt tabell C i bilagan.
4. Undantagna från skyldigheten att lämna produktionsdeklaration är även skördare som tillhör ett vinkooperativ som skall lämna produktionsdeklaration och som levererar hela sin druvskörd till kooperativet, men som förbehåller sig rätten att för sin familjs bruk framställa mindre än 10 hektoliter vin.
Oaktat bestämmelserna i artikel 4 får medlemsstater, som i enlighet med förordning (EEG) nr 2392/86 har upprättat ett fullständigt register över vinodlingar som uppdateras varje år eller ett annat liknande administrativt kontrollinstrument, undanta de fysiska eller juridiska personer, sammanslutningar av sådana personer eller skördare som avses i denna artikel från skyldigheten att deklarera areal.
1. Fysiska eller juridiska personer eller sammanslutningar av sådana personer, med undantag av privata konsumenter och detaljister, skall varje år till de behöriga myndigheter som har utsetts av medlemsstaterna deklarera de lager av druvmust, koncentrerad druvmust, rektifierad koncentrerad druvmust och vin som de innehar den 31 juli. Vinprodukter från gemenskapen skall inte tas med i denna deklaration om de framställts av druvor som skördats under innevarande kalenderår.
De mängder som avses i första stycket skall fastställas enskilt av varje medlemsstat med hänsyn till handelns och distributionens särskilda egenskaper.
1. Medlemsstaterna skall utarbeta formulär för de olika deklarationerna och säkerställa att dessa innehåller minst de uppgifter som anges i tabellerna A, B, C och D i bilagan.
Medlemsstaterna skall besluta om nödvändiga kontrollåtgärder för att säkerställa att deklarationerna överensstämmer med verkligheten.
- fått vissa av de uppgifter som skall anges i deklarationerna enligt kapitlen I och II från andra administrativa handlingar behöver inte kräva att dessa uppgifter skall finnas med i deklarationerna,
- fått vissa av de uppgifter som skall anges i deklarationerna enligt kapitel III från andra administrativa handlingar behöver inte kräva att dessa uppgifter skall finnas med i deklarationerna,
Vid utformningen av deklarationer enligt artiklarna 2 och 4 skall följande viner betraktas som "annat vin" vara vin som härrör från druvsorter som i medlemsstaternas klassificering i enlighet med artikel 19 i förordning (EG) nr 1493/1999, samtidigt för samma administrativa enhet anges som druvsorter för vinframställning och i förekommande fall som bordsdruvor, som druvsorter som är avsedda att torkas eller som sorter avsedda för framställning av vinsprit.
De produktmängder som skall tas upp i de deklarationer som avses i artiklarna 2, 4 och 6 skall uttryckas i hektoliter vin. De mängder koncentrerad druvmust och rektifierad koncentrerad druvmust som skall tas upp i de deklarationer som avses i artikel 4 skall uttryckas i hektoliter.
Den mängd vin som skall anges i de produktionsdeklarationer som föreskrivs i artikel 4 skall vara den totala mängd som erhålls efter huvudjäsningen, inklusive vindruv.
Artikel 11
Artikel 12
Artikel 13
a) När det gäller de åtgärder som avses i artiklarna 24, 34 och 35 i förordning (EG) nr 1493/1999, skall stödet minskas med
Stöd skall inte betalas ut om felet medför att den deklarerade volymen justeras med mer än 20 %, vare sig för vinåret i fråga eller för det därpå följande vinåret.
- Med samma procentsats som det konstaterade felet om felet medför att den deklarerade volymen justeras med 5 % eller mindre.
De behöriga myndigheterna skall anpassa de stöd som skall utbetalas till destillatören i förhållande till det pris som betalats till producenten.
a) En sammanställning på nationell nivå av de produktionsdeklarationer som avses i artikel 4 i denna förordning och om sådana finns, också av de koefficienter som används för att konvertera volymer av andra produkter än vin uttryckta i deciton till hektoliter vin för de olika produktionsområdena.
d) En bedömning för pågående vinår av uppgifter som gör det möjligt att uppskatta de tillgängliga mängderna vinprodukter och deras användning i medlemsstaten.
1. För prisnoteringarna skall medlemsstaterna, förutom de i vilka kapitlen I och II i avdelning II i förordning (EG) nr 1493/1999 inte tillämpas i enlighet med artikel 21 i den förordningen, definiera sammanhängande produktionsområden som omfattar flera mindre produktionsområden vars produktion är tillräckligt homogen.
4. Ovannämnda priser skall gälla en nettovara fritt producenten.
a) senast den 15 september och den 30 november under innevarande vinår, en bedömning av den volym vinprodukter som kan förväntas framställas i medlemsstaten enligt artikel 14 c,
d) den provisoriska försörjningsbalansen för senast föregående vinår senast den 15 november och den slutliga försörjningsbalansen för det näst senaste vinåret senast den 15 mars, enligt artikel 14 e; försörjningsbalanserna skall skickas till Eurostat, gemenskapens statistikkontor.
a) före den 1 augusti 2001:
- De platser som valts i varje produktionsområde för prisnotering.
Artikel 17
Utöver att de används för statistiska ändamål används uppgifterna i deklarationerna även vid tillämpningen av förordning (EG) nr 1493/1999. Särskilt uppgifter om uppdelningen av produktionen i bordsvin, kvalitetsvin fso och annat vin avgör rättigheter och skyldigheter för producenterna vid tillämpning av den förordningen.
Artikel 20
Det belopp som skall återvinnas fastställs enligt reglerna i artikel 12 i kommissionens förordning (EG) nr 1282/2001(7).
c) Producenten har inte fullgjort skyldigheterna i artikel 37 i förordning (EG) nr 1493/1999 och överträdelsen har konstaterats eller meddelats destillatören efter det att det lägsta priset har betalats på grundval av tidigare deklarationer.
Upphävanden
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av bilagorna I och III i rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I enlighet med förordning (EEG) nr 2377/90 måste gränsvärden för högsta tillåtna restmängder successivt fastställas för samtliga farmakologiskt verksamma substanser som används inom gemenskapen i veterinärmedicinska läkemedel som är avsedda att ges till livsmedelsproducerande djur.
(4) För kontroll av resthalter bör enligt tillämplig gemenskapslagstiftning gränsvärden vanligtvis fastställas för målvävnaderna lever eller njure. I den internationella handeln avlägsnas dock ofta lever och njure från slaktkroppen, och gränsvärden bör därför alltid fastställas även för muskel- eller fettvävnader.
(7) För att möjliggöra komplettering av vetenskapliga studier, bör giltighetstiden för temporär MRL, tidigare definierad i bilaga III till förordning (EEG) nr 2377/90, förlängas för cefalonium, morantel och metamizol.
Artikel 1
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av rådets förordning (EEG) nr 3880/91 om avlämnande av statistikuppgifter om nominell fångst för medlemsstater som bedriver fiske i Nordatlantens östra del
med beaktande av rådets förordning (EEG) nr 3880/91 av den 17 december 1991 om avlämnande av statistikuppgifter över nominell fångst för medlemsstater som bedriver fiske i Nordatlantens östra del(1), särskilt artikel 2.3 och artikel 4 i denna, och
(2) Vid sitt 87:e stadgeenliga sammanträde 1999 beslöt Internationella rådet för utnyttjande av havet (ICES) att uppta de artgrupper av Elasmobranchii-fiskar, som beskrivs i rapporten från arbetsgruppen om Elasmobranchii-arter, och uppmana FAO att införa dessa arter i sitt Statlant 27A-frågeformulär om fångststatistik för nordöstra Atlanten.
(5) Flera medlemsstater har begärt att få inlämna uppgifter i annan form eller med annat medium än enligt vad som som föreskrivs i bilaga IV till förordning (EG) nr 3880/91 (som motsvarar ovannämnda Statlant-frågeformulär).
Artikel 1
Medlemsstaterna får inlämna uppgifter i enlighet med det format som specificeras i bilaga II till denna förordning.
Kommissionens förordning (EG) nr 1660/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) I artiklarna 86-102 föreskrivs avsättningsregler för alkohol som innehas av interventionsorganen. Vissa sakfel bör rättas, bland annat bör priset för prover ändras. Vidare bör det för rektifieringsprodukter beviljas samma avvikelse för bioetanol som för nya industriella användningsområden.
Artikel 1
2. Artikel 63 skall ändras på följande sätt:
b) Följande punkt skall läggas till som punkt 10: "10. Det vin som levereras till destilleri skall destilleras senast den 30 september påföljande vinår."
a) under alla förhållanden till 15 %,
Interventionsorgan som innehar alkohol kan, i synnerhet av logistikskäl, ersätta alkohol i de behållare som anges i medlemsstaternas meddelande enligt punkt 1 i den här artikeln med en annan alkohol, som är av samma typ eller som blandats med annan alkohol som levererats till interventionsorganet fram till dess att en uttagsorder utfärdas. Medlemsstaternas interventionsorgan skall meddela kommissionen om att alkoholen ersatts."
b) Punkt 2 skall ersättas med följande: "2. Efter tidsfristen för inlämnande av anbud eller efter trettio dagar efter meddelandet om offentlig auktion
Dessa prover kan fås från interventionsorganet mot betalning av 10 euro per liter, varvid kvantiteten skall begränsas till 5 liter per behållare."
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EG) nr 174/1999 om fastställande av särskilda tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 i fråga om exportlicenser och exportbidrag inom sektorn för mjölk och mjölkprodukter och av förordning (EG) nr 1498/1999 om tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 beträffande meddelanden mellan medlemsstaterna och kommissionen med avseende på mjölk och mjölkprodukter
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), senast ändrad genom förordning (EG) nr 1670/2000(2), särskilt artikel 26.3, artikel 30, artikel 31.14 och artikel 40 i denna, och
(2) En rättelse bör göras av ett fel som insmugit sig i artikel 9 i förordning (EG) nr 174/1999.
(5) För att förenkla säkerheterna för de tillfälliga licenser som avses i artikel 20 är det lämpligt att justera säkerheterna för sådana licenser och att precisera hur säkerheterna för slutliga licenser skall fungera.
Artikel 1
2. I artikel 9 skall led a ersättas med följande: "a) 5 % för produkter med KN-nummer 0405."
5. Artikel 20.10 skall ersättas med följande: "10. Före utgången av det år för vilket de tillfälliga licenserna utfärdats skall den berörda parten, även om det rör sig om delkvantiteter, ansöka om en slutlig exportlicens som skall utfärdas omedelbart, varvid den säkerhet som avses i punkt 2 skall höjas till det totalbelopp som föreskrivs i artikel 9 för de kvantiteter för vilka licenser tilldelas. I ansökan om slutlig licens och i licensen skall följande anges i fält 20: 'För export till Amerikas förenta stater: artikel 20 i förordning (EG) nr 174/1999.'
Artikel 2
i) som avses i artikel 1 i förordning (EG) nr 174/1999, med undantag för sådana produkter som avses i artikel 17 i den förordningen (kod för IDES-meddelanden: 1),
d) I förekommande fall den justerade kvantiteten i en anbudsinfordran enligt b ovan."
Rådets förordning (EG) nr 2136/2001
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(2), och
(2) Kommissionen har lämnat en rapport till rådet om tilllämpningen av förordning (EG) nr 723/97 under perioden 1997-2000. Av de utvärderingsrapporter som sammanställts av medlemsstaterna och de genomförda programmens effektivitet drar kommissionen slutsatsen att medlemsstaterna bör få fortsatt finansiellt bidrag för att genomföra programmen enligt artikel 1 i förordning (EG) nr 723/97.
(5) Förordning (EG) nr 723/97 bör därför ändras.
Förordning (EG) nr 723/97 ändras på följande sätt:
av den 28 december 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen
(1) Spanien har i enlighet med artikel 5 i förordning (EEG) nr 2081/92 till kommissionen översänt en ansökan om registrering av "Manzana Reineta del Bierzo" som ursprungsbeteckning och en ansökan om registrering av "Salchichón de Vic" "Llonganissa de Vic" som geografisk beteckning.
(4) Dessa produktnamn kan därför tas upp i Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar och därmed vara skyddade inom gemenskapen såsom skyddad ursprungsbeteckning eller skyddad geografisk beteckning.
Artikel 1
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Jordnötter som har sitt ursprung i eller försänds från Kina har vid ett flertal tillfällen visat sig innehålla alltför höga halter av aflatoxin B1 eller alltför hög total aflatoxinhalt.
(4) Detta utgör en allvarlig fara för folkhälsan inom gemenskapen. Det är därför nödvändigt att anta skyddsåtgärder på gemenskapsnivå.
(7) De kinesiska myndigheterna bör se till att alla sändningar av jordnötter som har sitt ursprung i eller försänds från Kina åtföljs av skriftlig dokumentation som anger under vilka förhållanden varorna producerats, sorterats, hanterats, bearbetats, förpackats och transporterats samt resultaten från en laboratorieanalys av halterna av aflatoxin B1 och den totala aflatoxinhalten i sändningen.
(10) Ständiga livsmedelskommittén rådfrågades den 2 april 2001 och den 19 juli 2001.
1. Medlemsstaterna får inte importera produkter som tillhör nedanstående kategorier och som har sitt ursprung i eller försänds från Kina och är avsedda som livsmedel eller att användas som ingrediens i livsmedel, om inte sändningen åtföljs av resultaten av en officiell provtagning och analys samt av ett sådant hälsointyg som återges i bilaga I, ifyllt och undertecknat av en företrädare för den kinesiska myndigheten State Administration for Entry/Exit Inspection and Quarantine:
- Rostade jordnötter som omfattas av KN-nummer 2008 11 92 (i förpackningar med en nettovikt på mer än 1 kg) och KN-nummer 2008 11 96 (i förpackningar med en nettovikt på mindre än 1 kg).
4. De behöriga myndigheterna i varje medlemsstat skall se till att handlingarna för importerade jordnötter som har sitt ursprung i eller försänds från Kina kontrolleras, för att garantera att de krav på hälsointyg och provresultat som avses i punkt 1 är uppfyllda.
Europaparlamentets beslut
(2002/262/EG, EKSG, Euratom)
med beaktande av Fördraget om upprättandet av Europeiska kol- och stålgemenskapen, särskilt artikel 20 d.4,
med beaktande av kommissionens yttrande,
(1) Enligt artikel 22.5 i budgetförordningen av den 21 december 1977 för Europeiska gemenskapernas allmänna budget(2) skall ombudsmannen vid tillämpningen av denna förordning behandlas som en institution.
(4) Följaktligen bör artiklarna 12 och 16 i detta beslut utgå.
Artiklarna 12 och 16 i beslut 94/262/EKSG, EG och Euratom skall utgå.
av den 29 juli 2002
(2002/627/EG)
av följande skäl:
(3) De sätt på vilka de nationella regleringsmyndigheternas ansvar och uppgifter är fastlagda i detalj skiljer sig åt mellan medlemsstaterna, men gemensamt är att alla har minst en nationell regleringsmyndighet som har som uppdrag att tillämpa bestämmelserna - särskilt dem som rör den löpande tillsynen över marknaden - när de väl har omsatts i nationell lagstiftning.
(6) Gruppen bör fungera som en förmedlande länk mellan nationella regleringsmyndigheter och kommissionen på sådant sätt att den bidrar till den inre marknadens utveckling. I gruppen bör medlemsstaterna också kunna bedriva öppet redovisat samarbete med nationella regleringsmyndigheter och kommissionen för att på så sätt sörja för att regelverket för nät och tjänster inom området elektronisk kommunikation tillämpas på ett enhetligt sätt i alla medlemsstater.
(9) Verksamheten bör samordnas med arbetet i den radiospektrumkommitté som inrättats i enlighet med Europaparlamentets och rådets beslut nr 676/2002/EG av den 7 mars 2002 om ett regelverk för radiospektrumpolitiken i Europeiska gemenskapen (det s.k. radiospektrumbeslutet)(5), i den grupp för radiospektrumpolitik som inrättats i enlighet med kommissionens beslut 2002/622/EG av den 26 juli 2002 om inrättande av en grupp för radiospektrumpolitik(6) samt i den kontaktkommitté för television utan gränser som inrättats i enlighet med Europaparlamentets och rådets direktiv 97/36/EG av den 30 juni 1997 om samordning av vissa bestämmelser som fastställts i medlemsstaternas lagar och andra författningar om utförandet av sändningsverksamhet för television(7).
Innehåll
Definition
Arbetsuppgifter
Artikel 4
Kommissionen skall vara företrädd på en nivå som är avpassad till gruppens uppgifter, och kommissionen skall även tillhandahålla ett sekretariat för gruppens behov.
Gruppen skall - på eget initiativ eller på kommissionens begäran - ge råd till och bistå kommissionen i alla frågor som rör nät och tjänster inom området elektronisk kommunikation.
Gruppen skall enhälligt anta sin arbetsordning eller, om enhällighet inte kan uppnås, genom omröstning med två tredjedels majoritet, varvid varje medlemsstat har en röst, och arbetsordningen skall godkännas av kommissionen.
Artikel 6
Artikel 7
Artikel 8
Artikel 9
Kommissionens beslut
(2002/916/EG)
med beaktande av rådets direktiv 93/5/EEG av den 25 februari 1993 om hjälp till kommissionen och samarbete från medlemsstaternas sida vid den vetenskapliga granskningen av livsmedelsfrågor(1), särskilt artikel 3.2 fjärde strecksatsen i detta, och
(2) I kommissionens beslut 94/652/EG(3), senast ändrat genom beslut 2001/773/EG(4), fastställs inventeringen och fördelningen av uppgifterna inom ramen för medlemsstaternas samarbete vid den vetenskapliga granskningen av livsmedelsfrågor.
(5) Beslut 94/652/EG bör ändras i enlighet med detta.
Artikel 1
Detta beslut riktar sig till medlemsstaterna.
om inrättande av en allmän ram för information till och samråd med arbetstagare i Europeiska gemenskapen
med beaktande av kommissionens förslag(1),
i enlighet med förfarandet i artikel 251(4), på grundval av det gemensamma utkast som förlikningskommittén godkände den 23 januari 2002 och
(2) I punkt 17 i gemenskapsstadgan om arbetstagares grundläggande sociala rättigheter föreskrivs bland annat att "information till, samråd med och deltagande av arbetstagare måste utvecklas på ett lämpligt sätt med hänsyn till gällande förfaranden i de olika medlemsstaterna".
(5) Efter denna andra samrådsetapp har arbetsmarknadens parter inte underrättat kommissionen om att de önskar inleda det förfarande som kan leda till att ett avtal ingås.
(8) Det finns i synnerhet ett behov av att främja och stärka informationen och samrådet om den rådande situationen och den förväntade utvecklingen av sysselsättningen inom företaget och, när arbetsgivaren bedömer att sysselsättningen i företaget kan komma att hotas, om vilka eventuella föregripande åtgärder som planeras, i synnerhet i form av utbildning och kompetensutveckling för arbetstagarna, för att motverka den negativa utvecklingen eller mildra dess följder samt för att öka anställbarheten och anpassningsförmågan hos de arbetstagare som kan komma att påverkas.
(11) Den inre marknaden måste utvecklas på ett balanserat sätt med bibehållande av de viktiga värderingar som ligger till grund för våra samhällen, och genom att alla medborgare får del av den ekonomiska utvecklingen.
(14) Hela denna politiska, ekonomiska, sociala och rättsliga utveckling gör det nödvändigt att anpassa den befintliga rättsliga ramen inom vilken de rättsliga och praktiska instrument som gör det möjligt att utöva rätten till information och samråd föreskrivs.
(17) Eftersom målen för den planerade åtgärden, såsom den beskrivs ovan, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna, eftersom syftet är att inrätta en ram för information till och samråd med arbetstagare, vilken är anpassad till de nya europeiska förutsättningar som beskrivs ovan, och därför på grund av den planerade åtgärdens omfattning och verkningar bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
(20) Detta tar hänsyn till och påverkar inte andra nationella åtgärder och förfaranden som syftar till att främja en social dialog inom företag som inte omfattas av detta direktiv, och inom den offentliga förvaltningen
(23) Målet i detta direktiv uppnås genom inrättandet av en allmän ram med principer, definitioner och villkor för informationen och samrådet, som medlemsstaterna skall respektera och anpassa i förhållande till sina nationella förutsättningar, där det vid behov säkerställs att arbetsmarknadens parter får en ledande roll genom att de får rätt att genom avtal fritt fastställa de arrangemang för information och samråd som bäst överensstämmer med deras behov och önskemål.
(26) Arbetsgivaren bör ges möjlighet att underlåta att informera och samråda, när detta skulle innebära allvarlig skada för företaget eller driftstället eller när han omedelbart måste hörsamma en anvisning som en övervaknings- eller tillsynsmyndighet givit honom.
(29) Detta direktiv bör inte påverka andra mer specifika bestämmelser i rådets direktiv 98/59/EG av den 20 juli 1998 om tillnärmning av medlemsstaternas lagstiftning om kollektiva uppsägningar(5) och i rådets direktiv 2001/23/EG av den 12 mars 2001 om tillnärmning av medlemsstaternas lagstiftning om skydd för arbetstagares rättigheter vid överlåtelse av företag, verksamheter eller delar av företag eller verksamheter(6).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Detta direktiv syftar till att inrätta en allmän ram med minimikrav avseende arbetstagarnas rätt till information och samråd i företag eller driftställen inom gemenskapen.
Artikel 2
a) företag: offentligt eller privat företag som bedriver ekonomisk verksamhet med eller utan vinstsyfte och som är beläget inom medlemsstaternas territorium,
d) arbetstagare: varje person som i den berörda medlemsstaten åtnjuter skydd som arbetstagare inom ramen för den nationella arbetslagstiftningen och enligt nationell praxis,
g) samråd: diskussion och upprättande av en dialog mellan arbetstagarrepresentanterna och arbetsgivaren.
1. I enlighet med medlemsstaternas val skall detta direktiv tillämpas på
Medlemsstaterna skall själva besluta om hur tröskelvärdena för anställda arbetstagare skall beräknas.
Artikel 4
2. Information och samråd skall omfatta följande:
c) Information och samråd om beslut som kan medföra väsentliga förändringar i arbetsorganisationen eller anställningsavtalen, inklusive de beslut som avses i de gemenskapsbestämmelser som anges i artikel 9.1.
a) med säkerställande av att tillfället, sättet och innehållet är lämpligt,
d) på ett sådant sätt som gör det möjligt för arbetstagarrepresentanterna att sammanträda med arbetsgivaren och få motiverade svar på eventuella yttranden,
Avtalsreglerad information och avtalsreglerat samråd
Konfidentiell information
3. Utan att det påverkar befintliga nationella förfaranden skall medlemsstaterna säkerställa att det finns tillgång till rättsligt eller administrativt överklagandeförfarande i de fall arbetsgivaren hävdar att informationen är konfidentiell eller inte lämnar ut information i enlighet med punkt 1 och 2. De får dessutom införa förfaranden som säkerställer att den berörda informationen förblir konfidentiell.
Medlemsstaterna skall se till att arbetstagarrepresentanterna, när de utför sina uppdrag, får tillräckligt skydd och tillräckliga garantier, så att de på ett adekvat sätt kan utföra sina uppgifter.
1. Medlemsstaterna skall föreskriva lämpliga åtgärder för de fall då arbetsgivaren eller arbetstagarrepresentanterna inte följer detta direktiv. De skall särskilt se till att det finns administrativa eller rättsliga förfaranden för att säkerställa att de skyldigheter som följer av detta direktiv iakttas.
Förhållandet mellan detta direktiv och andra bestämmelser på gemenskapsnivå och nationell nivå
3. Detta direktiv skall inte påverka övriga gällande rättigheter till information, samråd och medverkan enligt nationell lagstiftning.
Övergångsbestämmelser
b) företag med minst 100 anställda eller driftställen med minst 50 anställda under det år som följer efter den tidpunkt som anges i a).
1. Medlemsstaterna skall anta de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 23 mars 2005 eller se till att arbetsmarknadens parter inför de nödvändiga bestämmelserna genom avtal, varvid medlemsstaterna skall var skyldiga att vidta alla nödvändiga åtgärder för att alltid kunna garantera de resultat som införs genom detta direktiv. De skall genast underrätta kommissionen om detta.
Översyn av kommissionen
Ikraftträdande
Adressater
av den 19 juli 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 95 i detta,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) Textilier och läderartiklar som innehåller vissa azofärgämnen kan avge arylaminer som kan innebära risk för cancer.
(5) För att skydda människors hälsa bör användning av farliga azofärgämnen och utsläppande på marknaden av vissa artiklar som färgats med sådana färgämnen förbjudas.
(8) Mot bakgrund av nya vetenskapliga rön bör analysmetoderna ses över, inbegripet metoder för att analysera 4-aminoazobensen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 5
av den 5 november 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 71 i detta,
efter att ha hört Regionkommittén,
(1) Säkerheten vid transporter samt miljöfrågor i samband med transporter är mycket viktiga för en hållbar rörlighet.
(4) Utvidgningen av tillämpningsområdet för direktiv 92/6/EEG till att omfatta fordon på över 3,5 ton avsedda för godstransport eller personbefordran var en av de åtgärder som rådet förordade i sin resolution av den 26 juni 2000 om ökad vägtrafiksäkerhet(5), i enlighet med kommissionens meddelande av den 20 mars 2000 om prioriteringar när det gäller vägtrafiksäkerheten inom Europeiska unionen.
(7) Direktiv 92/6/EEG bör ändras i enlighet härmed.
Direktiv 92/6/EEG ändras på följande sätt:
I detta direktiv avses med motorfordon sådana motordrivna fordon som tillhör någon av kategorierna M2, M3, N2 eller N3, är avsedda att användas på väg, har minst fyra hjul och är konstruerade för en högsta hastighet som överstiger 25 km/h.
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att de motorfordon i kategorierna M2 och M3 som avses i artikel 1 används på väg endast om de är utrustade med en hastighetsbegränsande anordning som ställts in så att fordonens hastighet inte kan överskrida 100 km/h.
1. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att motorfordon i kategorierna N2 och N3 används på väg endast om de är utrustade med en hastighetsbegränsande anordning som ställts in så att fordonens hastighet inte kan överskrida 90 km/h.
1. När det gäller motorfordon i kategori M3 med en totalvikt på över 10 ton och motorfordon i kategori N3, skall artiklarna 2 och 3 tillämpas på
i) från och med den 1 januari 1995 om det rör sig om fordon som används för såväl nationella som internationella transporter,
a) fordon som registrerats den 1 januari 2005 eller senare, från och med den 1 januari 2005,
ii) från och med den 1 januari 2007, om det rör sig om fordon som endast används för nationella transporter.
1. De hastighetsbegränsande anordningar som avses i artiklarna 2 och 3 skall uppfylla de tekniska krav som fastställs i bilagan till direktiv 92/24/EEG(8). Alla fordon som omfattas av det här direktivet och registrerats före den 1 januari 2005 får dock även i fortsättningen vara utrustade med sådana hastighetsbegränsande anordningar som uppfyller de tekniska krav som fastställts av de behöriga nationella myndigheterna.
"Artikel 6a
Artikel 2
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat och om ändring av rådets direktiv 73/239/EEG, 79/267/EEG, 92/49/EEG, 92/96/EEG, 93/6/EEG och 93/22/EEG samt Europaparlamentets och rådets direktiv 98/78/EG och 2000/12/EG
med beaktande av kommissionens förslag(1),
med beaktande av Europeiska centralbankens yttrande(3),
(1) Den nuvarande gemenskapslagstiftningen innehåller ett omfattande regelverk om tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag på enskild nivå samt över kreditinstitut, försäkringsföretag och värdepappersföretag som utgör en del av en bank- eller investeringsgrupp respektive en försäkringsgrupp, det vill säga grupper med en homogen finansiell verksamhet.
(4) Även inom andra internationella forum har behovet av att utveckla lämpliga tillsynsformer för finansiella konglomerat slagits fast.
(7) De behöriga myndigheterna bör kunna bedöma den finansiella ställningen på gruppnivå för kreditinstitut, försäkringsföretag och värdepappersföretag som ingår i ett finansiellt konglomerat, särskilt vad gäller solvens (inbegripet att eliminera dubbelt utnyttjande av poster i kapitalbasen), riskkoncentration och transaktioner inom det finansiella konglomeratet.
(10) Samordnarens uppgifter bör inte påverka de behöriga myndigheternas uppgifter och ansvar enligt särreglerna.
(13) Kreditinstitut, försäkringsföretag och värdepappersföretag som har sitt huvudkontor i gemenskapen kan ingå i ett finansiellt konglomerat vars ledande enhet ligger utanför gemenskapen. Dessa reglerade enheter bör också vara föremål för sådana likvärdiga och lämpliga ordningar för extra tillsyn som medför att liknande mål och resultat som de som anges i bestämmelserna i detta direktiv uppnås. Insyn i bestämmelserna och informationsutbyte med myndigheter i tredje land om alla viktiga omständigheter är här av stor vikt.
(16) Eftersom målet för den föreslagna åtgärden, nämligen att fastställa regler för extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och därför, på grund av den planerade åtgärdens omfattning eller verkningar, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå detta mål. Eftersom det i direktivet anges minimistandarder, kan medlemsstaterna införa strängare regler.
(19) Teknisk vägledning och genomförandeåtgärder för de bestämmelser som fastställs i detta direktiv kan ibland vara nödvändiga med hänsyn till ny utveckling på finansmarknaderna. Kommissionen bör följaktligen bemyndigas att anta genomförandeåtgärder, förutsatt att dessa inte ändrar det väsentliga innehållet i detta direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 2
1. kreditinstitut: ett kreditinstitut i den mening som avses i artikel 1.1 andra stycket i direktiv 2000/12/EG.
4. reglerad enhet: ett kreditinstitut, ett försäkringsföretag eller ett värdepappersföretag.
7. särregler: gemenskapslagstiftning som rör tillsynen över reglerade enheter, särskilt den som fastställs i direktiv 73/239/EEG, 79/267/EEG, 98/78/EG, 93/6/EEG, 93/22/EEG och 2000/12/EG.
b) Ett försäkringsföretag, ett återförsäkringsföretag eller ett försäkringsholdingbolag enligt artikel 1 led i i direktiv 98/78/EG (försäkringssektorn).
9. moderföretag:ett moderföretag i den mening som avses i artikel 1 i rådets sjunde direktiv 83/349/EEG av den 13 juni 1983 om sammanställd redovisning(15) och varje företag som enligt de behöriga myndigheterna i praktiken utövar ett bestämmande inflytande över ett annat företag.
12. grupp: en grupp av företag som består av ett moderföretag, dess dotterföretag och enheter i vilka moderföretaget och dess dotterföretag har ägarintressen samt företag som är knutna till varandra genom ett sådant förhållande som avses i artikel 12.1 i direktiv 83/349/EEG.
b) kontroll, innebärande förbindelse mellan ett moderföretag och ett dotterföretag i alla de fall som omfattas av artikel 1.1 och 1.2 i direktiv 83/349/EEG, eller en likartad förbindelse mellan någon fysisk eller juridisk person och ett företag. Varje dotterföretag till ett dotterföretag skall också anses som dotterföretag till moderföretaget vilket står över dessa företag.
a) En reglerad enhet i den mening som avses i artikel 1 finns i toppen av gruppen eller minst ett av dotterföretagen i gruppen är en reglerad enhet i den mening som avses i artikel 1.
d) Minst en av gruppens enheter ingår i försäkringssektorn och minst en i bank- eller värdepapperssektorn.
15. blandat finansiellt holdingföretag: ett moderföretag som inte utgör en reglerad enhet men som tillsammans med sina dotterföretag, varav minst ett är en reglerad enhet med huvudkontor inom gemenskapen, och andra enheter utgör ett finansiellt konglomerat.
a) de behöriga myndigheter i medlemsstaterna som har ansvar för den sektoriella tillsynen på gruppnivå över de reglerade enheterna i ett finansiellt konglomerat,
18. transaktioner inom det finansiella konglomeratet: alla transaktioner genom vilka reglerade enheter inom ett finansiellt konglomerat direkt eller indirekt anlitar andra företag inom samma grupp eller en fysisk eller juridisk person som har "nära förbindelser" med företagen i den gruppen, för att uppfylla en skyldighet, oavsett om den är avtalsenlig eller ej och om den sker mot betalning eller ej.
Tröskelvärden för identifiering av ett finansiellt konglomerat
I detta direktiv är den minsta finansiella sektorn i ett finansiellt konglomerat den sektor som har det lägsta genomsnittet och den mest betydande finansiella sektorn i ett finansiellt konglomerat den sektor som har det högsta genomsnittet. Vid beräkningen av genomsnittet för den minsta finansiella sektorn och den mest betydande finansiella sektorn skall banksektorn och värdepapperssektorn beaktas tillsammans.
b) Marknadsandelen överstiger inte 5 % i någon medlemsstat, mätt i termer av balansomslutningen för bank- och värdepapperssektorerna och i termer av tecknade bruttopremier inom försäkringssektorn.
a) undanta en enhet från beräkningen av procentsatserna i de fall som avses i artikel 6.5,
5. Vid tillämpningen av punkterna 1 och 2 får de relevanta behöriga myndigheterna, i exceptionella fall och i samförstånd, ersätta balansomslutningen som kriterium med en av följande parametrar eller båda eller lägga till en eller båda av dessa parametrar, om de anser att de är av särskild relevans för den extra tillsynen enligt detta direktiv: intäktsstruktur, poster utanför balansräkningen.
Under den period som avses i denna punkt får samordnaren, med medgivande från de övriga relevanta behöriga myndigheterna, besluta att de lägre procentsatser eller det lägre belopp som anges i denna punkt inte längre skall tillämpas.
Artikel 4
För detta ändamål
2. Den samordnare som utsetts enligt artikel 10 skall informera det moderföretag som finns i toppen av en grupp eller, i avsaknad av moderföretag, den reglerade enhet som har den största balansomslutningen inom den största finansiella sektorn i en grupp, om att gruppen har identifierats som ett finansiellt konglomerat och om utnämningen av samordnare. Samordnaren skall också informera de behöriga myndigheter som har auktoriserat reglerade enheter i gruppen och de behöriga myndigheterna i den medlemsstat i vilken det blandade finansiella holdingföretaget har sitt huvudkontor samt kommissionen.
AVSNITT I
Räckvidd för den extra tillsynen över de reglerade enheter som avses i artikel 1
a) Varje reglerad enhet i toppen av ett finansiellt konglomerat.
Om ett finansiellt konglomerat är en undergrupp till ett annat finansiellt konglomerat som uppfyller kraven i första stycket, får medlemsstaterna tillämpa artiklarna 6-17 enbart på reglerade enheter i den senare gruppen, och alla hänvisningar i direktivet till begreppen grupp och finansiellt konglomerat skall då anses syfta på denna.
För att sådan extra tillsyn skall kunna utövas, skall minst en av enheterna vara en reglerad enhet enligt artikel 1 och de villkor som anges i artikel 2.14 d och e skall vara uppfyllda. De relevanta behöriga myndigheterna skall fatta sitt beslut med beaktande av de mål för extra tillsyn som anges i detta direktiv.
AVSNITT 2
Kapitaltäckning
Medlemsstaterna skall också kräva att reglerade enheter följer en adekvat kapitaltäckningsstrategi på nivån finansiellt konglomerat.
Resultatet av beräkningen och relevanta uppgifter för beräkningen skall överlämnas till samordnaren av den reglerade enhet i den mening som avses i artikel 1 som finns i toppen av det finansiella konglomeratet eller, när det finansiella konglomeratet inte har en reglerad enhet i den mening som avses i artikel 1 i toppen, av det blandade finansiella holdingföretaget eller av den reglerade enhet i det finansiella konglomeratet som identifierats av samordnaren efter samråd med de övriga relevanta behöriga myndigheterna och med det finansiella konglomeratet.
b) Försäkringsföretag, återförsäkringsföretag eller försäkringsholdingbolag i den mening som avses i artikel 1 i i direktiv 98/78/EG.
4. Vid beräkning av de extra kapitaltäckningskraven avseende ett finansiellt konglomerat genom tillämpning av metod 1 (metod baserad på sammanställd redovisning) som avses i bilaga I skall kapitalbas och solvenskrav för enheterna i gruppen beräknas genom tillämpning av de motsvarande särregler för sammanställningens form och omfattning som fastställs framför allt i artikel 54 i direktiv 2000/12/EG och i punkt 1 B i bilaga I till direktiv 98/78/EG.
a) Om enheten finns i ett tredje land där det finns rättsliga hinder för att överföra erforderliga upplysningar, utan att detta påverkar tillämpningen av särreglernas bestämmelser om de behöriga myndigheternas skyldighet att vägra auktorisation när de är förhindrade att effektivt utöva sin tillsyn.
Om flera enheter utesluts till följd av b i första stycket, måste de dock inkluderas om de tillsammans inte är av försumbar betydelse.
Artikel 7
2. Medlemsstaterna skall kräva att reglerade enheter eller blandade finansiella holdingföretag regelbundet och minst en gång per år till samordnaren rapporterar varje betydande riskkoncentration på nivån finansiellt konglomerat enligt reglerna i denna artikel och i bilaga II. Den nödvändiga informationen skall överlämnas till samordnaren av den reglerade enhet i den mening som avses i artikel 1 som finns i toppen av det finansiella konglomeratet eller, när det finansiella konglomeratet inte leds av en reglerad enhet i den mening som avses i artikel 1, av det blandade finansiella holdingföretaget eller av den reglerade enhet i det finansiella konglomeratet som identifierats av samordnaren efter samråd med de övriga relevanta behöriga myndigheterna och med det finansiella konglomeratet.
4. När ett finansiellt konglomerat leds av ett blandat finansiellt holdingföretag, skall eventuella särregler om riskkoncentration i den största finansiella sektorn i det finansiella konglomeratet gälla för hela den sektorn, inklusive det blandade finansiella holdingföretaget.
1. Utan att särreglerna åsidosätts skall extra tillsyn över reglerade enheters transaktioner inom det finansiella konglomeratet, utövas enligt reglerna i artikel 9.2-9.4 i avsnitt 3 i detta kapitel och bilaga II.
Samordnaren skall övervaka dessa transaktioner inom det finansiella konglomeratet.
Artikel 9
2. Metoderna för riskhantering skall inbegripa följande:
c) Lämpliga förfaranden för att säkerställa att systemen för övervakning av risker är väl integrerade i organisationen och att alla åtgärder har vidtagits för att se till att de system som genomförts i alla de företag som omfattas av extra tillsyn är samstämmiga, så att riskerna kan mätas, övervakas och kontrolleras på nivån finansiellt konglomerat.
b) Sunda rapporterings- och redovisningsförfaranden, för att identifiera, mäta, övervaka och kontrollera transaktionerna inom det finansiella konglomeratet och riskkoncentrationen.
AVSNITT 3
Behörig myndighet ansvarig för utövandet av extra tillsyn (samordnaren)
a) Om ett finansiellt konglomerat leds av en reglerad enhet, skall samordningen utövas av den behöriga myndighet som har auktoriserat denna reglerade enhet enligt gällande särregler.
ii) Om två eller flera reglerade enheter med huvudkontor inom gemenskapen har samma blandade finansiella holdingföretag som moderföretag och en av dessa enheter har auktoriserats i den medlemsstat där det blandade finansiella holdingföretaget har sitt huvudkontor, skall samordningen utövas av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som auktoriserats i denna medlemsstat.
iii) Om två eller flera reglerade enheter med huvudkontor inom gemenskapen har samma blandade finansiella holdingföretag som moderföretag och ingen av dessa enheter har auktoriserats i den medlemsstat där det blandade finansiella holdingföretaget har sitt huvudkontor, skall samordningen utövas av den behöriga myndighet som har auktoriserat den reglerade enhet som har den största balansomslutningen inom den största finansiella sektorn.
Artikel 11
a) Samordning av insamling och spridning av relevanta eller väsentliga uppgifter, såväl löpande som i krissituationer, inbegripet spridning av uppgifter som är av betydelse för en behörig myndighets tillsynsuppgifter enligt särreglerna.
d) Bedömning av det finansiella konglomeratets struktur, organisation och system för intern kontroll enligt artikel 9.
För att den extra tillsynen skall kunna underlättas och få en bred rättslig grund, skall samordnaren, de andra relevanta behöriga myndigheterna och vid behov andra berörda behöriga myndigheter införa samordningsåtgärder. Genom dessa kan samordnaren anförtros ytterligare uppgifter och förfaranden specificeras för de relevanta behöriga myndigheternas beslutsprocesser enligt artiklarna 3 och 4, artikel 5.4, artikel 6, artikel 12.2 samt artiklarna 16 och 18, samt för samarbetet med andra behöriga myndigheter.
Artikel 12
Detta samarbete skall åtminstone omfatta insamling och utbyte av uppgifter avseende följande punkter:
c) Det finansiella konglomeratets finansiella ställning, särskilt när det gäller kapitaltäckning, transaktioner inom det finansiella konglomeratet, riskkoncentration och lönsamhet.
f) Förfaranden för insamling av uppgifter från enheterna i ett finansiellt konglomerat samt kontroll av de uppgifterna.
När det är nödvändigt för utförandet av deras respektive uppgifter, kan de behöriga myndigheterna också utbyta uppgifter om reglerade enheter i ett finansiellt konglomerat med följande myndigheter i enlighet med bestämmelserna i särreglerna: centralbanker, Europeiska centralbankssystemet och Europeiska centralbanken.
b) Större sanktioner eller exceptionella åtgärder som de behöriga myndigheterna vidtar.
Om de uppgifter som avses i artikel 14.2 redan har lämnats till en behörig myndighet enligt särreglerna, kan de behöriga myndigheter som ansvarar för att utöva extra tillsyn vända sig till den förstnämnda myndigheten för att erhålla dessa uppgifter.
Artikel 13
Artikel 14
2. Medlemsstaterna skall föreskriva att deras behöriga myndigheter med ansvar för att utöva extra tillsyn skall få tillgång till alla uppgifter som kan vara relevanta för den extra tillsynen, genom att direkt eller indirekt vända sig till enheterna i ett finansiellt konglomerat, vare sig dessa är reglerade enheter eller ej.
Om de behöriga myndigheterna vid tillämpningen av detta direktiv i specifika fall önskar kontrollera uppgifter om en reglerad eller icke reglerad enhet i en annan medlemsstat vilken ingår i ett finansiellt konglomerat, skall de begära att de behöriga myndigheterna i denna medlemsstat låter utföra kontrollen.
Artikel 16
- av samordnaren när det gäller det blandade finansiella holdingföretaget,
Då så krävs skall de berörda behöriga myndigheterna, inklusive samordnaren, samordna sina tillsynsåtgärder.
1. I avvaktan på ytterligare harmonisering av särreglerna skall medlemsstaterna se till att de behöriga myndigheterna har befogenhet att vidta alla tillsynsåtgärder som anses nödvändiga för att undvika eller bemöta att reglerade enheter i ett finansiellt konglomerat kringgår särreglerna.
TREDJE LÄNDER
1. Utan att detta påverkar särreglerna skall de behöriga myndigheterna i det fall som avses i artikel 5.3 kontrollera huruvida reglerade enheter, vilkas moderföretag har huvudkontor utanför gemenskapen, är föremål för sådan tillsyn som utövas av en behörig myndighet i tredje land som är likvärdig med den extra tillsyn som föreskrivs i detta direktiv beträffande sådana reglerade enheter som avses i artikel 5.2. Kontrollen skall utföras av den behöriga myndighet som skulle vara samordnare om kriterierna i artikel 10.2 hade varit tillämpliga, på begäran av moderföretaget eller av någon av de reglerade enheter som auktoriserats i gemenskapen eller på egen begäran. Den behöriga myndigheten skall samråda med de andra relevanta behöriga myndigheterna och beakta varje tillämplig vägledning som Kommittén för finansiella konglomerat har utarbetat enligt artikel 21.5. Den behöriga myndigheten skall med anledning därav rådfråga kommittén innan beslut fattas.
Artikel 19
2. Kommissionen, Rådgivande bankrörelsekommittén, Försäkringskommittén och Kommittén för finansiella konglomerat skall granska resultatet av de förhandlingar som avses i punkt 1 och den därigenom uppkomna situationen.
Artikel 20
a) En mer precis formulering av definitionerna i artikel 2 i syfte att beakta utvecklingen på finansmarknaderna vid tillämpningen av detta direktiv.
d) En mer precis definition av beräkningsmetoderna i bilaga I för att beakta utvecklingen på finansmarknaderna och av tillsynsmetoderna.
Artikel 21
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av artikel 8 i det beslutet.
4. Utan att det påverkar redan antagna genomförandeåtgärder, skall tillämpningen av de bestämmelser i detta direktiv i vilka föreskrivs att tekniska regler och beslut skall antas i enlighet med förfarandet i punkt 2 upphöra fyra år efter det att detta direktiv har trätt i kraft. Europaparlamentet och rådet kan på förslag av kommissionen förnya bestämmelserna i fråga i enlighet med förfarandet i artikel 251 i fördraget och skall därvid granska dem före utgången av ovannämnda period.
KAPITEL IV
Ändringar av direktiv 73/239/EEG
"Artikel 12a
b) är dotterföretag till moderföretaget till ett försäkringsföretag som är auktoriserat i en annan medlemsstat, eller
a) är dotterföretag till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen,
3. De relevanta behöriga myndigheter som avses i punkterna 1 och 2 skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla de uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet som är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
a) Ägarintressen som försäkringsföretaget har i
- försäkringsholdingbolag i den mening som avses i artikel 1 led i i direktiv 98/78/EG,
b) Var och en av följande poster som ett försäkringsföretag innehar i de enheter som definierats i a i vilka det har ägarintresse:
- Fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 i direktiv 2000/12/EG.
För beräkningen av solvensmarginalen enligt detta direktiv får medlemsstaterna föreskriva att försäkringsföretag som är föremål för extra tillsyn enligt direktiv 98/78/EG eller direktiv 2002/87/EG inte behöver dra ifrån poster enligt a och b i fjärde stycket i de kreditinstitut, värdepappersföretag, finansiella institut, försäkrings- eller återförsäkringsföretag eller försäkringsholdingbolag som ingår i den extra tillsynen.
Ändringar av direktiv 79/267/EEG
"Artikel 12a
b) är dotterföretag till moderföretaget till ett försäkringsföretag som är auktoriserat i en annan medlemsstat, eller
a) är dotterföretag till ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen,
3. De relevanta behöriga myndigheter som avses i punkterna 1 och 2 skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla de uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet som är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
a) Ägarintressen som försäkringsföretaget har i
- försäkringsholdingbolag i den mening som avses i artikel 1 led i i direktiv 98/78/EG,
b) Var och en av följande poster som ett försäkringsföretag innehar i de enheter som definierats under a i vilka det har ägarintresse:
- Fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 i direktiv 2000/12/EG.
Artikel 24
1. I artikel 15 skall följande punkt införas:
"5c. Denna artikel skall inte hindra en behörig myndighet från att
överföra uppgifter för att dessa skall kunna utföra sina uppgifter, och den skall inte heller hindra sådana myndigheter eller organ från att vidarebefordra sådana uppgifter som de kan behöva enligt punkt 4. Uppgifter som erhålls i detta sammanhang skall omfattas av de bestämmelser om tystnadsplikt som fastställs i denna artikel.".
Direktiv 92/96/EEG skall ändras på följande sätt:
2. Artikel 15.5c skall ersättas med följande:
- i förekommande fall till andra myndigheter med ansvar för övervakning av betalningssystem,
Ändring av direktiv 93/6/EEG
- holdingföretag med blandad verksamhet: ett moderföretag som inte utgör ett finansiellt holdingföretag, ett värdepappersföretag eller ett blandat finansiellt holdingföretag i den mening som avses i direktiv 2002/87/EG, bland vars dotterföretag det finns minst ett värdepappersföretag.".
Direktiv 93/22/EEG ändras på följande sätt:
a) är dotterföretag till ett kreditinstitut eller försäkringsföretag som är auktoriserat i gemenskapen,
De relevanta behöriga myndigheter som avses i första och andra stycket skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla de uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet som är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
Artikel 28
1. I artikel 1 skall g, h, i och j ersättas med följande:
i) försäkringsholdingbolag: ett moderföretag vars huvudsakliga verksamhet består i att förvärva och ha ägarintresse i dotterföretag, vilka enbart eller huvudsakligen är försäkringsföretag, återförsäkringsföretag eller försäkringsföretag i tredje land, där minst ett av dotterföretagen är ett försäkringsföretag, och vilket inte är ett blandat finansiellt holdingföretag i den mening som avses i Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(30).
"Den behöriga myndighet som har framställt begäran får om den så önskar delta i kontrollen, om den inte själv utför den.".
4. Följande artiklar skall läggas till:
1. Kommissionen kan antingen på begäran av en medlemsstat eller på eget initiativ ställa förslag till rådet i fråga om förhandlingar om avtal med ett eller flera tredje länder om metoderna för att utöva extra tillsyn över
2. Av de avtal som avses i punkt 1 skall särskilt framgå både
3. Kommissionen och Försäkringskommittén skall granska resultaten av de förhandlingar som avses i punkt 1 och den därigenom uppkomna situationen.
Medlemsstaterna skall kräva att de personer som faktiskt leder affärsverksamheten i ett holdingföretag med blandad verksamhet har ett tillräckligt gott anseende och tillräcklig erfarenhet för att kunna fullgöra dessa åligganden.".
6. I punkt 2 i bilaga I skall följande punkt läggas till:
Artikel 29
1. Artikel 1 skall ändras på följande sätt:
b) Punkterna 21 och 22 skall ersättas med följande:
2. I artikel 12 skall följande stycken läggas till:
b) är dotterföretag till moderföretaget till ett försäkringsföretag som är auktoriserat i gemenskapen, eller
3. Artikel 16.2 skall ersättas med följande:
a) I det första stycket skall punkterna 12 och 13 ersättas med följande:
14. Ägarposter i andra kreditinstitut och finansiella institut, motsvarande högst 10 % av deras kapital, fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 som ett kreditinstitut innehar hos andra kreditinstitut och finansiella institut än de som anges i punkterna 12 och 13 i detta stycke, i den mån dessa ägarposter, fordringar och instrument tillsammans överstiger 10 % av kreditinstitutets kapitalbas beräknad före avdrag för posterna enligt punkterna 12-16 i detta stycke.
- återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG,
- de instrument som avses i artikel 16.3 i direktiv 73/239/EEG,
"Om aktier i ett annat kreditinstitut, finansiellt institut, försäkringsföretag, återförsäkringsföretag eller försäkringsholdingföretag innehas tillfälligt i syfte att ge finansiellt bistånd för att rekonstruera och rädda denna enhet, får den behöriga myndigheten bevilja undantag från bestämmelserna om avdrag i punkterna 12-16.
Denna bestämmelse skall tillämpas på alla försiktighetsregler som är harmoniserade genom gemenskapsakten.".
6. Artikel 52.2 sista meningen skall ersättas med följande:
a) I punkt 1 skall följande stycke läggas till:
8. Följande artikel skall införas:
Medlemsstaterna skall kräva att de personer som faktiskt leder affärsverksamheten i ett finansiellt holdingföretag har ett tillräckligt gott anseende och tillräcklig erfarenhet för att kunna fullgöra dessa åligganden.".
Transaktioner inom det finansiella konglomeratet med holdingföretag med blandad verksamhet
Om ovannämnda transaktioner inom det finansiella konglomeratet utgör ett hot mot kreditinstitutets finansiella ställning, skall den behöriga myndighet som ansvarar för tillsynen över institutet vidta lämpliga åtgärder.".
11. Följande artikel skall läggas till:
Om ett kreditinstitut, vars moderföretag är ett kreditinstitut eller ett finansiellt holdingföretag med huvudkontor utanför gemenskapen, inte är föremål för gruppbaserad tillsyn enligt artikel 52, skall de behöriga myndigheterna kontrollera huruvida kreditinstitutet är föremål för gruppbaserad tillsyn av en behörig myndighet i tredje land, vilken är likvärdig med den som styrs av de principer som anges i artikel 52. Kontrollen skall utföras av den behöriga myndighet som skulle vara ansvarig för den extra tillsynen om fjärde stycket hade varit tillämpligt, på begäran av moderföretaget eller av någon av de reglerade enheter som auktoriserats i gemenskapen eller på eget initiativ. Denna behöriga myndighet skall samråda med de andra berörda behöriga myndigheterna.
KAPITEL V
Kapitalförvaltningsbolag
b) tillämpningsområdet för extra tillsyn i den mening som avses i detta direktiv, om gruppen är ett finansiellt konglomerat.
KAPITEL VI
Rapport från kommissionen
- vilka kapitaltäckningsmetoder i bilaga I som bör väljas och hur de bör tillämpas,
Kommissionen skall samråda med kommittén innan den lägger fram sina förslag.
Införlivande
Ikraftträdande
Adressater
av den 16 december 2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av rådets direktiv 86/363/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på livsmedel av animaliskt ursprung(3), senast ändrat genom direktiv 2002/79/EG, särskilt artikel 10 i detta,
av följande skäl:
(3) Om det inte finns något permanent eller provisoriskt gränsvärde för bekämpningsmedelsrester på gemenskapsnivå måste medlemsstaterna fastställa ett provisoriskt nationellt gränsvärde i enlighet med artikel 4.1 f i direktiv 91/414/EEG innan växtskyddsmedel som innehåller detta verksamma ämne kan godkännas.
(6) Även om gemenskapen fastställer sådana provisoriska gränsvärden hindrar detta inte att medlemsstaterna själva fastställer provisoriska gränsvärden enligt artikel 4.1 f i direktiv 91/414/EEG och bilaga VI till det direktivet. Fyra år anses vara en tillräckligt lång period för att utveckla ytterligare användningsområden för de berörda verksamma ämnena. De provisoriska gränsvärdena bör därefter bli permanenta.
(9) Detta direktiv är förenligt med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
Följande gränsvärde för bekämpningsmedelsrester skall läggas till i del A i bilaga II till direktiv 86/362/EEG:
Följande gränsvärden för bekämpningsmedelsrester skall läggas till i del B i bilaga II till direktiv 86/363/EEG:
Gränsvärdena för bekämpningsmedelsrester av de berörda verksamma ämnena i bilagan till detta direktiv skall läggas till i bilaga II till direktiv 90/642/EEG.
De skall tillämpa dessa bestämmelser från och med den 1 juli 2003.
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Kommissionens förordning (EG) nr 204/2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Med anledning av revideringen av Harmoniserade systemet och Kombinerade nomenklaturen (HS/KN) enligt kommissionens förordning (EG) nr 2031/2001 av den 6 augusti 2001 om ändring av bilaga I till rådets förordning (EEG) nr 2658/87 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(3) är det nödvändigt att göra ändringar i CPA samt att anpassa och förtydliga texterna.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för det statistiska programmet.
Bilagan till förordning (EEG) nr 3696/93 skall ersättas med bilagan till den här förordningen.
Kommissionens förordning (EG) nr 315/2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Priset skall vara det som noteras på den eller de representativa marknaderna i varje medlemsstat för de olika kategorierna av färska eller kylda slaktkroppar av får. I de medlemsstater som har mer än en representativ marknad bör det aritmetiska eller, om nödvändigt, det viktade genomsnittet av de priser som har noterats på dessa marknader användas.
(6) För att förklara de grunder på vilka medlemsstaterna genererar priserna skall de lämna uppgifter till kommissionen om den valda representativa marknaden och kategorierna av slaktkroppar samt vikten eller den relativa betydelsen av de uppgifter som används för att beräkna priserna.
Artikel 1
Artikel 2
2. Priserna på slaktkroppar av lamm som väger mellan 9 och 16 kg kan dock noteras före borttagande av slaktbiprodukter och huvud i överensstämmelse med normal handelspraxis.
Artikel 3
3. Om det inte finns någon tillgänglig information skall dock priserna på medlemsstatens representativa marknader fastställas med hjälp särskilt av de senast noterade priserna.
a) Varje prisnoteringsområdes representativa marknader.
Medlemsstaterna skall underrätta kommissionen om eventuella ändringar i förfarandena senast en månad efter det att ändringarna gjorts.
Artikel 6
av den 25 mars 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Grekland har i enlighet med artikel 5 i förordning (EEG) nr 2081/92 till kommissionen översänt en ansökan om registrering av "Πατατα Κατω Νευροκοπιου" (Patata Kato Nevrokopiou) som geografisk beteckning.
(4) Detta produktnamn kan därför tas upp i "Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar" och därmed vara skyddat inom gemenskapen såsom skyddad geografisk beteckning.
Artikel 1
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EG) nr 3063/93 om tillämpningsföreskrifter för rådets förordning (EEG) nr 2019/93 angående stödordningen för produktion av kvalitetshonung
med beaktande av rådets förordning (EEG) nr 2019/93 av den 19 juli 1993 om införandet av särskilda bestämmelser för de mindre Egeiska öarna rörande vissa jordbruksprodukter(1), senast ändrad genom förordning (EG) nr 442/2002(2), särskilt artikel 12.3 i denna, och
(2) I syfte att aktualisera förordning (EG) nr 3063/93 bör de undantag för år 1993 strykas som berör sista ansökningsdag, sista utbetalningsdag för stöd och sista datum för inlämnande av uppgifter till kommissionen om utbetalade stöd och andelen stödansökningar som omfattas av kontroll på plats. Dessutom bör hänvisningen till jordbruksomräkningskursen strykas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) I punkt 1 skall andra stycket utgå.
5. Artikel 5 skall ändras på följande sätt:
b) Det andra stycket utgå.
Artikel 2
av den 27 juni 2002
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) Byrån bör allmänt sett fungera som ett tekniskt organ, som gör det möjligt för gemenskapen att agera effektivt för att förbättra bestämmelserna om den övergripande sjösäkerheten och förhindrandet av förorening från fartyg. Byrån bör bistå kommissionen i det fortgående arbetet med att uppdatera och utveckla gemenskapens lagstiftning när det gäller området för sjösäkerhet och förhindrande av förorening från fartyg och tillhandahålla det stöd som behövs för att se till att lagstiftningen tillämpas enhetligt och effektivt i hela gemenskapen genom att bistå kommissionen i utförandet av de uppgifter som den tilldelats genom nuvarande och framtida gemenskapslagstiftning om sjösäkerhet och förhindrande av förorening från fartyg.
(6) För att byrån skall kunna utföra sina arbetsuppgifter på vederbörligt sätt, bör dess tjänstemän besöka medlemsstaterna för att kontrollera att gemenskapens system för sjösäkerhet och förhindrande av förorening från fartyg fungerar. Besöken bör genomföras i enlighet med en praxis som byråns styrelse fastställer, och de bör underlättas av medlemsstaternas myndigheter.
(9) För att effektivt kunna se till att byrån fullgör sina uppgifter bör medlemsstaterna och kommissionen vara företrädda i en styrelse som har de befogenheter som är nödvändiga för att fastställa budgeten och kontrollera att den genomförs, anta lämpliga finansiella bestämmelser, utarbeta tydliga förfaranden för byråns beslutsfattande, godkänna dess arbetsprogram, behandla ansökningar från medlemsstater om tekniskt bistånd, fastställa riktlinjer för besök i medlemsstaterna samt utnämna den verkställande direktören. Med tanke på denna särskilda byrås synnerligen tekniska och vetenskapliga uppdrag och uppgifter bör styrelsen bestå av en företrädare för varje medlemsstat och fyra företrädare för kommissionen som är ledamöter med en hög nivå av sakkunskap. För att ytterligare säkerställa högsta möjliga nivå när det gäller sakkunskap och erfarenhet i styrelsen och för att de mest berörda branschsektorerna skall kunna delta aktivt i byråns verksamhet, bör kommissionen utnämna oberoende yrkesverksamma personer inom dessa sektorer som ledamöter i styrelsen, utan rösträtt, på grundval av personliga meriter och personlig erfarenhet inom området för sjösäkerhet och förhindrande av förorening från fartyg och inte som företrädare för särskilda branschorganisationer.
(12) I takt med att allt fler decentraliserade organ har inrättats på senare år har budgetmyndigheten de gångna åren försökt förbättra insynen i och kontrollen av förvaltningen av gemenskapsanslagen till organen, särskilt när det gäller budgetering av avgifter, finansiell kontroll, befogenheter att bevilja ansvarsfrihet, avsättning till pensionssystemet samt det interna budgetförfarandet (uppförandekodex). På liknande sätt bör Europaparlamentets och rådets förordning (EG) nr 1073/1999 av den 25 maj 1999 om utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF)(6) oinskränkt tillämpas när det gäller byrån, som bör ansluta sig till det interinstitutionella avtalet av den 25 maj 1999 mellan Europaparlamentet, Europeiska unionens råd och Europeiska gemenskapernas kommission om interna utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF)(7).
KAPITEL I
Mål
Artikel 2
a) Den skall vid behov bistå kommissionen i det förberedande arbetet med att uppdatera och utveckla gemenskapslagstiftningen när det gäller sjösäkerhet och förhindrande av förorening från fartyg, särskilt med beaktande av den internationella lagstiftningens utveckling på området. I denna uppgift ingår att analysera forskningsprojekt som utförs inom området för sjösäkerhet och förhindrande av förorening från fartyg.
ii) ge kommissionen det tekniska stöd den behöver för att delta i arbetet i de tekniska arbetsgrupper som inrättats inom ramen för det i Paris ingångna samförståndsavtalet om hamnstatskontroll (the Paris Memorandum of Understanding on Port State Control),
i) vid behov anordna relevant utbildningsverksamhet på områden som står under hamnstatens och flaggstatens ansvar,
i) främja samarbete mellan kuststater i de sjöfartsområden som omfattas av det direktivet,
f) Byrån skall förse kommissionen och medlemsstaterna med objektiva, tillförlitliga och jämförbara uppgifter och data om sjösäkerhet och förorening från fartyg, så att dessa kan vidta nödvändiga åtgärder för att förbättra sjösäkerheten [och förhindrandet av förorening från fartyg] och utvärdera befintliga åtgärders effektivitet. I dessa uppgifter ingår att samla in, registrera och utvärdera tekniska data om sjösäkerhet, sjöfart och marina föroreningar, oavsiktliga eller avsiktliga, att systematiskt utnyttja och samköra befintliga databaser och att vid behov skapa nya databaser. Byrån skall, på grundval av insamlade data, bistå kommissionen när den var sjätte månad offentliggör uppgifter om fartyg som vägrats tillträde till hamnar i gemenskapen med tillämpning av rådets direktiv 95/21/EG av den 19 juni 1995 om tillämpning av internationella normer för säkerhet på fartyg, förhindrande av förorening samt boende- och arbetsförhållanden ombord på fartyg som anlöper gemenskapens hamnar och framförs i medlemsstaternas territorialvatten (hamnstatskontroll)(8). Byrån skall också bistå kommissionen och medlemsstaterna i deras verksamhet för att förbättra identifiering och lagföring av fartyg som gjort sig skyldiga till olagliga utsläpp.
Besök i medlemsstaterna
3. Efter varje besök skall byrån upprätta en rapport och skicka den till kommissionen och den berörda medlemsstaten.
1. Byrån skall tillämpa principerna i Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar(9), när den behandlar ansökningar om tillgång till de handlingar som den innehar.
4. Den information som kommissionen och byrån samlar in i enlighet med denna förordning skall omfattas av Europaparlamentets och rådets förordning (EG) nr 45/2001 av den 18 december 2000 om skydd för enskilda då gemenskapsinstitutionerna och gemenskapsorganen behandlar personuppgifter och om den fria rörligheten för sådana uppgifter(10).
Artikel 5
2. Byrån skall i varje medlemsstat ha den mest vittgående rättskapacitet som tillerkänns juridiska personer enligt den nationella lagstiftningen. Den skall särskilt kunna förvärva och avyttra lös och fast egendom samt föra talan inför domstolar och andra myndigheter.
Artikel 6
2. Om inte annat föreskrivs i artikel 16, skall byrån, när det gäller dess egen personal, utöva de befogenheter som enligt tjänsteföreskrifterna och anställningsvillkoren för övriga anställda tillkommer tillsättningsmyndigheten.
Privilegier och immunitet
Ansvar
3. Vad beträffar utomobligatoriskt ansvar skall byrån, i enlighet med de allmänna principer som är gemensamma för medlemsstaternas rättsordningar, ersätta skada som orsakats av dess enheter eller av dess anställda under tjänsteutövning.
Artikel 9
2. De översättningar som krävs för byråns arbete skall utföras av Översättningscentrum för Europeiska unionens organ.
1. En styrelse inrättas härmed för byrån.
b) senast den 30 april varje år anta byråns allmänna rapport för föregående år och skicka den till medlemsstaterna, Europaparlamentet, rådet och kommissionen,
Detta arbetsprogram skall antas utan att det påverkar gemenskapens årliga budgetförfarande. Om kommissionen inom 15 dagar från den tidpunkt då arbetsprogrammet antagits meddelar att den inte samtycker till det antagna arbetsprogrammet, skall styrelsen behandla det igen och inom två månader, vid den andra behandlingen, anta det eventuellt ändrade arbetsprogrammet, antingen med två tredjedels majoritet, inbegripet kommissionens företrädare, eller med enhällighet bland medlemsstaternas företrädare,
g) fastställa riktlinjer för de besök som skall genomföras enligt artikel 3,
j) fastställa sin arbetsordning.
1. Styrelsen skall bestå av en företrädare för varje medlemsstat och fyra företrädare för kommissionen samt av fyra yrkesverksamma personer som kommissionen utsett inom de mest berörda sektorerna, vilka personer inte skall ha rösträtt.
3. Mandatperioden skall vara fem år. Mandatet kan förnyas en gång.
Styrelsens ordförande
Artikel 13
2. Byråns verkställande direktör skall delta i överläggningarna.
5. Styrelsen får bjuda in alla personer vars åsikter kan vara av intresse att delta som observatörer vid sammanträdena.
Artikel 14
2. Varje ledamot skall ha en röst. Den verkställande direktören får inte rösta.
Artikel 15
2. Den verkställande direktören skall ha följande arbetsuppgifter och befogenheter:
c) Han/hon skall vidta nödvändiga åtgärder för att se till att byrån fungerar i enlighet med bestämmelserna i denna förordning, bl.a. genom att anta anvisningar för den interna administrationen och offentliggöra meddelanden.
f) Han/hon skall göra beräkningar av byråns intäkter och utgifter i enlighet med artikel 18 och genomföra budgeten i enlighet med artikel 19.
Utnämning av verkställande direktör
2. Den verkställande direktörens mandatperiod skall vara fem år. Mandatet får förnyas en gång.
1. Tredjeländer får delta i byråns arbete, om de genom avtal med Europeiska gemenskapen har antagit och tillämpar gemenskapslagstiftningen inom området för sjösäkerhet och förhindrande av förorening från fartyg.
FINANSIELLA KRAV
1. Byråns intäkter skall bestå av
c) avgifter för publikationer, utbildning och/eller andra tjänster som byrån tillhandahåller.
4. Intäkter och utgifter skall balansera varandra.
6. När budgetmyndigheten har antagit Europeiska unionens allmänna budget, skall styrelsen anta byråns budget och slutliga arbetsprogram och vid behov anpassa dem till gemenskapens bidrag. Den skall utan dröjsmål överlämna dem till kommissionen, budgetmyndigheten och de tredjeländer som deltar i byråns arbete.
1. Den verkställande direktören skall genomföra byråns budget.
Revisionsrätten skall granska räkenskaperna i enlighet med artikel 248 i fördraget. Den skall årligen offentliggöra en rapport om byråns verksamhet.
Bekämpning av bedrägeri
3. I beslut om finansiering samt i de avtal om och instrument för genomförande som ingåtts till följd av dessa beslut skall det uttryckligen föreskrivas att revisionsrätten och OLAF vid behov skall få utföra kontroller på plats hos dem som mottagit anslag från byrån och hos de ombud som fördelat dessa anslag.
Styrelsen skall, efter att ha mottagit kommissionens godkännande och revisionsrättens yttrande, anta byråns budgetförordning. I denna budgetförordning skall det särskilt anges vilket förfarande som skall användas vid utarbetandet och genomförandet av byråns budget i enlighet med artikel 142 i budgetförordningen av den 21 december 1977 för Europeiska gemenskapernas allmänna budget(12).
Artikel 22
2. I utvärderingen skall det bedömas i vilken utsträckning förordningen, byrån och dess arbetsmetoder bidragit till att etablera en hög sjösäkerhetsnivå och en hög nivå på förhindrandet av förorening från fartyg. Styrelsen skall utarbeta särskilda riktlinjer i samförstånd med kommissionen och efter samråd med de berörda parterna.
Inledande av byråns verksamhet
Ikraftträdande
Europaparlamentets och rådets förordning (EG) nr 1774/2002
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) Mot bakgrund av dessa vetenskapliga yttranden bör det göras skillnad mellan de åtgärder som skall vidtas beroende på vilken typ av animaliska biprodukter som används. De möjliga användningsområdena för vissa animalieprodukter bör begränsas. Regler bör fastställas för annan användning av animaliska biprodukter än i foder och för bortskaffandet av dessa.
(6) I Europaparlamentets resolution om BSE och säkert djurfoder av den 16 november 2000(5) krävde Europaparlamentet ett förbud mot användning av animaliskt protein i foder fram till dess att denna förordning träder i kraft.
(9) Sedan oktober 1996 har kontoret för livsmedels- och vetrinärfrågor (FVO) genomfört ett antal inspektioner i medlemsstaterna för att ta reda på vilka de viktigaste riskfaktorerna är och hur dessa hanteras samt hur övervakningen av BSE sker. Bedömningen gällde bland annat systemen för kommersiell konvertering och andra metoder för att hantera animaliskt avfall. Dessa inspektioner har utmynnat i allmänna slutsatser och ett antal rekommendationer, särskilt beträffande möjligheten att spåra animaliska biprodukter.
(12) Särskilda bestämmelser bör fastställas om kontroll av bearbetningsanläggningar, särskilt när det gäller detaljförfaranden för validering av bearbetningsmetoder och för egentillsyn av produktionen.
(15) För att säkerställa att hälsobestämmelserna genomförs på ett enhetligt sätt bör gemenskapsinspektioner utföras i medlemsstaterna. Sådana inspektioner bör också omfatta kontrollförfaranden.
(18) Mot bakgrund av vad som angetts ovan verkar det vara nödvändigt att göra en genomgripande revidering av de av gemenskapens bestämmelser som gäller animaliska biprodukter.
(21) Animaliska biprodukter som passerar gemenskapen i transit, eller som har sitt ursprung i gemenskapen och är avsedda för export, kan medföra risk för djurs och människors hälsa inom gemenskapen. Vissa krav som fastställs i denna förordning bör därför tillämpas på sådan befordran.
(24) Rådet och kommissionen har antagit flera beslut om genomförande av direktiven 90/667/EEG och 92/118/EEG. Direktiv 92/118/EEG har dessutom ändrats på ett genomgripande sätt, och ytterligare ändringar skall göras. Följaktligen finns det för närvarande ett stort antal gemenskapsrättsakter som reglerar sektorn för animaliska biprodukter och det finns behov av förenkling.
(27) Produkter som importeras till gemenskapen bör genomgå noggranna kontroller. Detta kan uppnås genom tillämpning av de kontroller som fastställs i rådets direktiv 97/78/EG av den 18 december 1997 om principerna för organisering av veterinärkontroller av produkter från tredje land som förs in i gemenskapen(12).
(30) De åtgärder som krävs för att genomföra denna förordning bör antas enligt rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(16).
b) utsläppande på marknaden samt, i vissa särskilda fall, export och transitering av animaliska biprodukter och därav framställda produkter enligt bilagorna VII och VIII.
b) Flytande mjölk och råmjölk som bortskaffats eller använts på det ursprungliga jordbruksföretaget.
e) Matavfall såvida inte detta
iii) är avsett att användas i en biogasanläggning eller för kompostering.
3. Denna förordning skall inte påverka tillämpningen av sådan veterinärlagstiftning som syftar till att utrota och bekämpa vissa sjukdomar.
1. I denna förordning avses med
c) kategori 2-material: animaliska biprodukter som avses i artikel 5.
f) produktionsdjur: alla djur som hålls, göds eller föds upp av människor och används för framställning av livsmedel (bland annat kött, mjölk och ägg), ull, päls, fjädrar, skinn eller andra produkter av animaliskt ursprung.
i) behörig myndighet: den centrala myndighet i en medlemsstat som har till uppgift att se till att kraven i denna förordning följs, eller någon annan myndighet till vilken denna centrala myndighet har delegerat denna befogenhet, särskilt när det gäller kontroll av djurfoder. Den skall även i tillämpliga fall inbegripa motsvarande myndighet i tredje land.
l) transitering: en befordran genom gemenskapen från ett tredje land till ett annat.
o) specificerat riskmaterial: det material som avses i bilaga V till Europaparlamentets och rådets förordning (EG) nr 999/2001 av den 22 maj 2001 om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati(17).
Allmänna skyldigheter
3. Medlemsstaterna skall, antingen var för sig eller i samarbete, se till att det finns ändamålsenliga arrangemang och tillräcklig infrastruktur för att säkerställa att kravet i punkt 1 uppfylls.
i) Djur som misstänks vara infekterade med TSE enligt förordning (EG) nr 999/2001 eller som officiellt bekräftats vara infekterade med TSE.
iv) Försöksdjur enligt definitionen i artikel 2 i rådets direktiv 86/609/EEG av den 24 november 1986 om tillnärmning av medlemsstaternas lagar och andra författningar om skydd av djur som används för försök och andra vetenskapliga ändamål(18).
ii) Hela kroppar från döda djur som innehåller specificerat riskmaterial om det specificerade riskmaterialet inte har avlägsnats vid tidpunkten för bortskaffandet.
e) Matavfall som härrör från transportmedel i internationell trafik.
a) direkt bortskaffas som avfall genom förbränning i en förbränningsanläggning som godkänts i enlighet med artikel 12,
d) när det gäller matavfall enligt punkt 1 e bortskaffas som avfall genom nedgrävning på en deponi som godkänts i enlighet med direktiv 1999/31/EG, eller
4. Kategori 1-material får endast importeras eller exporteras i enlighet med denna förordning eller regler som fastställts i enlighet med förfarandet i artikel 33.2. Import eller export av specificerat riskmaterial får emellertid endast ske i enlighet med artikel 8.1 i förordning (EG) nr 999/2001.
1. Kategori 2-material skall omfatta animaliska biprodukter som motsvarar följande beskrivning och allt material som innehåller sådana biprodukter:
c) Produkter av animaliskt ursprung som innehåller restsubstanser av veterinärmedicinska läkemedel och föroreningar som förtecknas i grupperna B.1 och B.2 i bilaga I till direktiv 96/23/EG, om restsubstanserna av dessa ämnen överskrider gällande gränsvärden enligt gemenskapslagstiftningen.
f) Blandningar av kategori 2- och kategori 3-material, inbegripet allt material som är avsett för bearbetning i en bearbetningsanläggning för kategori 2-material.
a) direkt bortskaffas som avfall genom förbränning i en förbränningsanläggning som godkänts i enlighet med artikel 12,
ii) när det gäller utsmält fett, bearbetas vidare till fettderivat för användning i organiska gödningsmedel eller jordförbättringsmedel eller för annan teknisk användning, förutom i kosmetika, läkemedel och medicintekniska produkter, i en kategori 2-oleokemisk anläggning som godkänts i enlighet med artikel 14,
ii) omvandlas i en biogas- eller komposteringsanläggning som godkänts i enlighet med artikel 15, eller
e) när det gäller naturgödsel, från mag- och tarmsystemet avskilt mag- och tarminnehåll, mjölk och råmjölk om den behöriga myndigheten inte anser att det medför risk för spridning av allvarliga överförbara sjukdomar,
iii) omvandlas i en biogasanläggning eller komposteras i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2,
3. Mellanhantering eller mellanlagring av kategori 2-material med undantag av naturgödsel får bara genomföras på hanteringsställen för kategori 2 som godkänts i enlighet med artikel 10.
Kategori 3-material
b) Delar från slaktade djur som förklaras otjänliga som livsmedel trots att de inte visar några tecken på sjukdomar som kan överföras till människor eller djur, och som kommer från slaktkroppar som är tjänliga som livsmedel i enlighet med gemenskapslagstiftningen.
e) Animaliska biprodukter som erhållits vid framställning av produkter som är avsedda som livsmedel, exempelvis avfettade ben och fettgrevar.
h) Fisk och andra havslevande djur, utom havslevande däggdjur, som fångats på öppet hav för tillverkning av fiskmjöl.
k) Blod, hudar, skinn, hovar, fjädrar, ull, horn, hår och päls från djur som inte visat några kliniska tecken på sådana sjukdomar som kan överföras till människor eller djur via produkten i fråga.
a) direkt bortskaffas som avfall genom förbränning i en förbränningsanläggning som godkänts i enlighet med artikel 12,
d) omvandlas i en teknisk anläggning som godkänts i enlighet med artikel 18,
g) när det gäller matavfall enligt punkt 1 l, omvandlas i en biogasanläggning eller komposteras i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2, eller i väntan på att sådana bestämmelser skall antas, i enlighet med nationell lagstiftning,
3. Mellanhantering eller mellanlagring av kategori 3-material får bara genomföras på hanteringsställen för kategori 3 som godkänts i enlighet med artikel 10.
1. Animaliska biprodukter och bearbetade produkter, med undantag för matavfall av kategori 3, skall samlas in, transporteras och identifieras i enlighet med bilaga II.
4. I enlighet med artikel 4 i rådets direktiv 75/442/EEG av den 15 juli 1975 om avfall(21) skall medlemsstaterna vidta nödvändiga åtgärder för att se till att matavfall av kategori 3 insamlas, transporteras och bortskaffas utan att människors hälsa äventyras eller miljön skadas.
Artikel 8
2. Mottagande medlemsstat skall ha godkänt att ta emot kategori 1-material, kategori 2-material, bearbetade produkter som härrör från kategori 1- eller kategori 2-material och bearbetat animaliskt protein. Medlemsstaten får ställa som krav för mottagandet att bearbetningsmetod 1 skall tillämpas före avsändandet.
b) transporteras direkt till den mottagande anläggningen, som skall ha godkänts i enlighet med denna förordning.
6. Den mottagande medlemsstaten skall genom regelbundna kontroller se till att de berörda anläggningarna i det egna landet endast använder sändningarna för godkända ändamål och att de för ett fullständigt register som visar att denna förordning har följts.
1. Den som avsänder, transporterar eller tar emot animaliska biprodukter skall föra register över sändningarna. Registren skall innehålla de upplysningar och bevaras under den tid som anges i bilaga II.
1. Hanteringsställen för material i kategori 1, 2 och 3 skall godkännas av den behöriga myndigheten.
b) hantera och lagra kategori 1- eller kategori 2-material i enlighet med kapitel II del B i bilaga III,
3. För att kunna godkännas skall ett hanteringsställe för kategori 3-material
c) genomgå hanteringsställets egenkontroll på det sätt som föreskrivs i artikel 25,
Godkännande av lagringsanläggningar
a) uppfylla kraven i kapitel III i bilaga III,
Godkännande av förbrännings- och samförbränningsanläggningar
a) de allmänna kraven i kapitel I i bilaga IV,
d) kraven i kapitel IV i bilaga IV beträffande restsubstanser,
3. För att godkännas av den behöriga myndigheten för bortskaffande av animaliska biprodukter, skall en förbränningsanläggning eller samförbränningsanläggning med låg kapacitet som inte omfattas av direktiv 2000/76/EG
c) uppfylla de allmänna villkoren i kapitel I i bilaga IV,
f) uppfylla de tillämpliga temperaturmätningskraven i kapitel V i bilaga IV, och
5. Kraven i punkterna 2 och 3 får ändras med beaktande av nya vetenskapliga rön i enlighet med förfarandet i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén.
1. Bearbetningsanläggningar för kategori 1- och kategori 2-material skall godkännas av den behöriga myndigheten.
b) hantera, bearbeta och lagra kategori 1- eller kategori 2-material i enlighet med kapitel II i bilaga V samt kapitel I i bilaga VI,
e) kontrolleras av den behöriga myndigheten i enlighet med artikel 26,
Artikel 14
a) bearbeta utsmält fett som härrör från kategori 2-material i enlighet med kraven i kapitel III i bilaga VI,
d) kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
Artikel 15
2. För att kunna godkännas skall biogas- och komposteringsanläggningar
c) kontrolleras av den behöriga myndigheten i enlighet med artikel 26,
3. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
1. Medlemsstaterna skall vidta alla åtgärder som behövs för att säkerställa att de animaliska biprodukter, och därav framställda produkter som avses i bilagorna VII och VIII, inte avsänds från något jordbruksföretag som ligger i en zon som är föremål för restriktioner som införts sedan zonen drabbats av en sjukdom för vilken den djurart som produkterna härrör från är mottaglig, eller från någon anläggning eller zon från vilka förflyttning eller handel skulle medföra risker för den djurhälsostatus som berör medlemsstaterna eller vissa områden i medlemsstaterna, utom då produkterna hanteras i enlighet med denna förordning.
b) inte har slaktats i en anläggning där det vid tidpunkten för slakt fanns djur som var infekterade eller som misstänktes vara infekterade med någon av de sjukdomar som omfattas av de bestämmelser som avses i punkt a.
b) har genomgått en behandling som är tillräcklig för att eliminera de aktuella djurhälsoriskerna i enlighet med denna förordning vid en anläggning som har godkänts för detta ändamål av den medlemsstat där djurhälsoproblemet förekom,
Andra villkor än de som anges i första stycket får fastställas i särskilda situationer genom beslut som antas i enlighet med det förfarande som avses i artikel 33.2. I sådana beslut skall de åtgärder som rör djuren eller de prov som djuren skall bli föremål för beaktas, liksom de egenskaper hos sjukdomen som är kännetecknande för arten i fråga, och alla åtgärder som krävs för att säkerställa skyddet av djurhälsan i gemenskapen skall specificeras.
1. Bearbetningsanläggningar för kategori 3-material skall godkännas av den behöriga myndigheten.
b) hantera, bearbeta och lagra endast kategori 3-material i enlighet med kapitel II i bilaga V och bilaga VII,
e) kontrolleras av den behöriga myndigheten i enlighet med artikel 26,
Artikel 18
2. För att en anläggning för tillverkning av sällskapsdjursfoder eller en teknisk anläggning skall kunna godkännas, skall följande krav vara uppfyllda:
ii) införa och genomföra rutiner för övervakning och kontroll av kritiska kontrollpunkter i de processer som används,
v) underrätta den behöriga myndigheten om resultatet av den laboratorieanalys som avses i iii eller annan information som de ansvariga för anläggningen har tillgång till, visar att det föreligger allvarlig fara för djurs eller människors hälsa.
Artikel 19
a) har framställts i en bearbetningsanläggning för kategori 3-material som har godkänts och står under tillsyn i enlighet med artikel 17,
d) uppfyller de särskilda kraven i bilaga VII.
1. Medlemsstaterna skall se till att sällskapsdjursfoder, tuggben, tekniska produkter, med undantag av dem som avses i punkterna 2 och 3, samt de animaliska biprodukter som avses i bilaga VIII släpps ut på marknaden eller exporteras endast om de
ii) om en produkt kan användas både som en teknisk produkt och som foderråvara och bilaga VIII inte innehåller några särskilda krav, uppfyller de särskilda kraven i det relevanta kapitlet i bilaga VII,
3. Medlemsstaterna skall se till att fettderivat som är framställda av kategori 2-material släpps ut på marknaden eller exporteras endast om de
c) uppfyller eventuella särskilda krav i bilaga VIII.
Artikel 10 i direktiv 90/425/EEG skall tillämpas på de produkter som omfattas av bilagorna VII och VIII till denna förordning.
1. Följande användningar av animaliska biprodukter och bearbetade produkter skall vara förbjudna:
c) Användning av andra typer av organiska gödningsmedel eller jordförbättringsmedel än naturgödsel på betesmark.
Undantag när det gäller användning av animaliska biprodukter
b) Användning av animaliska biprodukter för taxidermiska ändamål i tekniska anläggningar som godkänts för detta syfte i enlighet med artikel 18.
i) Kategori 2-material under förutsättning att det kommer från djur som inte avlivats eller dött till följd av bekräftad eller förmodad förekomst av en sjukdom som kan överföras till människor eller djur.
i) djurparksdjur,
iv) pälsdjur,
vii) fluglarver som skall användas som fiskagn.
a) användningen av de undantag som avses i punkt 2,
Den behöriga myndigheten skall utöva tillsyn över de i föregående stycke omnämnda användarnas och uppsamlingscentralernas anläggningar och skall när som helst kunna få tillträde till alla delar av anläggningarna, för att kunna kontrollera att de krav som avses i punkt 2 har uppfyllts.
Artikel 24
a) döda sällskapsdjur omedelbart får bortskaffas som avfall genom nedgrävning,
ii) kategori 2-material,
2. Inget undantag får beviljas för kategori 1-material som avses i artikel 4.1 a i.
a) huruvida de använder möjligheterna enligt punkt 1 b när det gäller kategori 1- och kategori 2-material,
a) säkerställa att förbränningen eller nedgrävningen av animaliska biprodukter inte hotar djurs eller människors hälsa,
Artikel 25
a) identifiera och kontrollera de kritiska kontrollpunkterna i anläggningarna,
i) varje bearbetad sats uppfyller produktkraven enligt denna förordning, och
e) införa ett system som säkerställer att varje avsänt parti kan spåras.
b) fastställa orsakerna till att bestämmelserna inte uppfyllts,
e) göra fler provtagningar och kontroller av produktionen,
3. Närmare bestämmelser för genomförandet av denna artikel, inbegripet regler om hur ofta kontroller skall ske och om referensmetoder för mikrobiologiska analyser, får fastställas i enlighet med förfarandet i artikel 33.2.
1. Den behöriga myndigheten skall genomföra regelbundna inspektioner och utöva regelbunden tillsyn vid anläggningar som godkänts i enlighet med denna förordning. Inspektioner och tillsyn vid bearbetningsanläggningar skall utföras i enlighet med kapitel IV i bilaga V.
4. Varje medlemsstat skall upprätta en förteckning över de anläggningar på dess territorium som godkänts i enlighet med denna förordning. Varje anläggning skall av medlemsstaten tilldelas ett officiellt nummer som identifierar anläggningen med hänsyn till den typ av verksamhet som bedrivs. Medlemsstaten skall sända kopior av förteckningen samt uppdaterade versioner till kommissionen och övriga medlemsstater.
Gemenskapens kontroller i medlemsstaterna
Allmänna bestämmelser
Artikel 29
2. De produkter som avses i bilagorna VII och VIII får importeras till eller transiteras genom gemenskapen endast om de uppfyller kraven i punkterna 3-6.
När förteckningen upprättas skall särskilt följande beaktas:
c) De faktiska hälsovillkor som tillämpas på produktion, framställning, hantering, lagring och avsändande av produkter av animaliskt ursprung som är avsedda för gemenskapen.
f) Resultatet från eventuella gemenskapsinspektioner i det tredje landet.
i) De bestämmelser om förebyggande och bekämpning av infektiösa eller smittsamma djursjukdomar som gäller i det tredje landet samt tillämpningen av dessa, inklusive bestämmelser om import från andra länder.
a) Kommissionen skall underrätta medlemsstaterna om det tredje landets förslag till ändringar av förteckningen över anläggningar inom fem arbetsdagar från det att förslaget till ändringar från det tredje landet tagits emot.
d) Om kommissionen inte har erhållit några synpunkter från medlemsstaterna inom den tidsfrist som anges i punkt b, skall medlemsstaterna anses ha godtagit ändringarna i förteckningen. Kommissionen skall underrätta medlemsstaterna om dessa ändringar inom fem arbetsdagar, och import från de berörda anläggningarna skall vara tillåten fem arbetsdagar efter det att medlemsstaterna tagit emot denna underrättelse.
7. I väntan på att förteckningen enligt punkt 4 skall upprättas och att de förlagor till intyg som avses i punkt 6 skall antas, får medlemsstaterna behålla de kontroller som föreskrivs i direktiv 97/78/EG och de intyg som föreskrivs enligt gällande nationella bestämmelser.
1. I enlighet med förfarandet i artikel 33.2 får det fattas ett beslut genom vilket det erkänns att de hälsobestämmelser som tillämpas av ett tredje land, en grupp av tredje länder eller en region i ett tredje land vid produktion, framställning, hantering, lagring och transport av en eller flera av de produktkategorier som avses i bilagorna VII och VIII, innebär garantier som är likvärdiga med dem som tillämpas i gemenskapen förutsatt att det tredje landet kan visa detta på ett objektivt sätt.
a) vilken typ av hälsointyg som skall åtfölja produkten samt intygets innehåll,
3. Närmare bestämmelser för tillämpningen av denna artikel skall fastställas i enlighet med förfarandet i artikel 33.2.
1. Experter från kommissionen får, när så är lämpligt, tillsammans med experter från medlemsstaterna genomföra kontroller på plats för att
i) villkoren för införande i en gemenskapsförteckning över tredje länder,
iv) alla slags nödåtgärder som tillämpas med stöd av gemenskapslagstiftningen.
3. Hur ofta samt på vilket sätt kontrollerna i punkt 1 skall utföras får fastställas i enlighet med förfarandet i artikel 33.2.
Ändring av bilagor samt övergångsbestämmelser
Artikel 33
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i beslutet.
Artikel 34
Artikel 35
2. I synnerhet skall medlemsstaterna informera kommissionen om de åtgärder som vidtas för att se till att bestämmelserna i denna förordning iakttas senast ett år efter dess ikraftträdande. På grundval av den information som den erhåller skall kommissionen lägga fram en rapport för Europaparlamentet och rådet, i förekommande fall åtföljd av lagförslag.
Finansiella arrangemang
Upphävande
Artikel 38
Kommissionens förordning (EG) nr 1802/2002
(Text av betydelse för EES)
med beaktande av rådets direktiv 92/65/EEG av den 13 juli 1992 om fastställande av djurhälsokrav i handeln inom och importen till gemenskapen av djur, sperma, ägg (ova) och embryon som inte faller under de krav som fastställs i de specifika gemenskapsregler som avses i bilaga A.I till direktiv 90/425/EEG(1), senast ändrat genom kommissionens förordning (EG) nr 1282/2002(2), särskilt artikel 22 i detta, och
(2) För att ge tillräckligt med tid för att de nya bestämmelserna skulle kunna införas i samtliga medlemsstater borde det ha fastställts ett datum då förordning (EG) nr 1282/2002 skulle börja att tillämpas.
(5) Det är nödvändigt att rättelsen gäller från och med det datum då förordning (EG) nr 1282/2002 träder i kraft.
Artikel 1
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
om rättelse av förordning (EG) nr 2200/96 när det gäller startdatum för övergångsperioden för erkännande av producentorganisationer
med beaktande av kommissionens förslag(1),
av följande skäl:
(3) Således bör nämnda misstag i artikel 13.1 i förordning (EG) nr 2200/96 rättas. Eftersom effekterna av misstaget kan ha haft negativa effekter för producentorganisationer som har utnyttjat övergångsperioderna bör motsvarande bestämmelser tillämpas från och med tillämpningsdatumet för förordning (EG) nr 2200/96.
Artikel 13.1 i förordning (EG) nr 2200/96 skall ersättas med följande: "1. De producentorganisationer som före den här förordningens ikraftträdande har erkänts med stöd av förordning (EEG) nr 1035/72, och som inte utan en övergångsperiod kan erkännas med stöd av artikel 11 i den här förordningen, får fortsätta att verka inom ramen för avdelning IV under två år från och med den 1 januari 1997, om dessa organisationer uppfyller kraven i berörda artiklar i förordning (EEG) nr 1035/72."
Kommissionens förordning (EG) nr 1921/2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Artikel 8 i förordning (EEG) nr 3149/92, som inte längre tillämpas eftersom ersättning för transportkostnaderna betalas ut på basis av faktiska utgifter, bör utgå.
Artikel 1
2. Artikel 5 skall ersättas med följande:
För nötkött skall bokföringsvärdet vara detsamma som gällande interventionspris den 30 juni 2002. Detta pris skall multipliceras med den koefficient som anges i bilagan.
3. Artikel 8 skall utgå.
Kommissionens förordning (EG) nr 1947/2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"- Italien: Milano".
Europaparlamentets och rådets förordning (EG) nr 2099/2002
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) COSS roll består av att centralisera uppgifterna för de kommittéer som inrättats enligt gemenskapslagstiftningen om sjösäkerhet, förhindrande av förorening från fartyg och skydd av boende- och arbetsförhållanden ombord på fartyg samt att bistå och ge kommissionen råd i alla frågor som rör sjösäkerhet och förebyggande eller minskning av miljöföroreningar från sjöfartsverksamhet.
(6) De åtgärder som behövs för att genomföra nämnda lagstiftning bör antas i enlighet med beslut 1999/468/EG.
(9) Skillnad måste emellertid göras mellan sådana bestämmelser i en gemenskapsrättsakt för vilkas tillämpning det hänvisas till ett internationellt instrument och sådana gemenskapsbestämmelser som ordagrant återger ett internationellt instrument helt eller delvis. I det sistnämnda fallet kan de senaste ändringarna av internationella instrument ändå inte tillämpas på gemenskapsnivå förrän de berörda gemenskapsbestämmelserna har ändrats.
(12) Ett särskilt förfarande för kontroll av överensstämmelse bör dock införas, så att kommissionen, efter samråd med COSS, kan vidta nödvändiga åtgärder för att undvika att ändringar av internationella instrument blir oförenliga med nämnda gällande lagstiftning eller gemenskapspolitik på områdena sjösäkerhet, förhindrande av förorening från fartyg samt skydd av boende- och arbetsförhållanden ombord på fartyg, eller med de mål som eftersträvas i denna lagstiftning. Ett sådant förfarande bör även göra det möjligt att förhindra att internationella ändringar försämrar den sjösäkerhet som uppnåtts inom gemenskapen.
Artikel 1
a) centralisera uppgifterna för de kommittéer som inrättats enligt gemenskapens sjöfartslagstiftning och som upphävs genom denna förordning, genom inrättande av en enda kommitté för sjösäkerhet och förhindrande av förorening från fartyg, kallad COSS,
Definitioner
b) Rådets direktiv 93/75/EEG.
e) Rådets direktiv 95/21/EG av den 19 juni 1995 om hamnstatskontroll.(14)
h) Rådets direktiv 97/70/EG av den 11 december 1997 om att införa harmoniserade säkerhetsregler för fiskefartyg som har en längd av 24 meter och däröver.(16)
k) Rådets direktiv 1999/35/EG av den 29 april 1999 om ett system med obligatoriska besiktningar för en säker drift av ro-ro-passagerarfartyg och höghastighetspassagerarfartyg i reguljär trafik.(19)
n) Europaparlamentets och rådets direktiv 2001/96/EG av den 4 december 2001 om fastställande av harmoniserade krav och förfaranden för säker lastning och lossning av bulkfartyg.(22)
Inrättande av en kommitté
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara en månad.
Genomförande i gemenskapens lagstiftning av ändringar av internationella instrument
Förfarande för kontroll av överensstämmelse
Förfarandet för kontroll av överensstämmelse får användas enbart för att ändra gemenskapens sjöfartslagstiftning på de områden som uttryckligen omfattas av det föreskrivande förfarandet och strikt inom ramen för kommissionens genomförandebefogenheter.
Förfarandet för kontroll av överensstämmelse, i förekommande fall inbegripet förfarandena enligt artikel 5.6 i beslut 1999/468/EG, skall slutföras senast en månad innan den period löper ut som fastställts internationellt för underförstått godkännande av ändringen i fråga eller senast en månad före den planerade tidpunkten för ändringens ikraftträdande.
Information
COSS befogenheter
Ändring av förordning (EEG) nr 613/91
"a) Konventioner: 1974 års internationella konvention om säkerheten för människoliv till sjöss (Solas 1974), 1996 års internationella lastlinjekonvention (LL 66) och den internationella konventionen om förhindrande av förorening från fartyg (Marpol 73/78), i gällande version, och tillhörande bindande resolutioner, som har antagits av Internationella sjöfartsorganisationen (IMO)."
1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i Europaparlamentets och rådets förordning (EG) nr 2099/2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(23).
3. Kommittén skall själv anta sin arbetsordning.
Artikel 9
1. Artikel 3 g skall ersättas med följande:
3. Artikel 7 skall ersättas med följande:
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(26) tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 10
1. Följande stycke skall läggas till i artikel 9:"Ändringarna av de internationella instrument som avses i artikel 2 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i Europaparlamentets och rådets förordning (EG) nr.../2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(27)."
1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i förordning (EG) nr 2099/2002.
3. Kommittén skall själv anta sin arbetsordning."
Förordning (EG) nr 417/2002 ändras på följande sätt:
3. Följande stycke läggas till i artikel 11:"Ändringarna av de internationella instrument som avses i artikel 3.1 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i förordning (EG) nr 2099/2002."
Kommissionens förordning (EG) nr 2104/2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från kommittén för det statistiska programmet, inrättad genom rådets beslut 89/382/EEG, Euratom(5).
Artikel 4.1 h i rådets förordning (EG) nr 577/98 skall ersättas med följande:
- nivå
- total längd
- om den senaste undervisningsaktiviteten skett på arbetstid
- inriktning för denna högsta nivå av utbildning
Koderna för de variabler för utbildning som skall användas för överföring av data under 2003 och framgent som anges i bilagan till denna förordning, ersätter motsvarande variabler i bilagan till kommissionens förordning (EG) nr 1575/2000.
Kommissionens beslut
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Många framsteg har gjorts sedan nätverket för europeiska arbetsförmedlingar (EURES-nätverket) inrättades genom kommissionens beslut 93/569/EEG(3) om genomförandet av rådets förordning (EEG) nr 1612/68.
(4) De möjligheter som ny informations- och kommunikationsteknik ger att ytterligare förbättra och rationalisera de tjänster som erbjuds bör också beaktas.
(7) För tydlighetens skull är det lämpligt att återupprätta EURES-nätverket och samtidigt tydligare fastställa dess sammansättning, uppbyggnad och funktioner. Detta innebär att beslut 93/569/EEG bör ersättas.
Artikel 1
Artikel 2
EURES-nätverket skall särskilt till förmån för arbetssökande, arbetstagare och arbetsgivare sträva efter att främja
c) öppenhet och utbyte av information om europeiska arbetsmarknader, inklusive om levnadsvillkor och utbildningsmöjligheter,
Sammansättning
b) EURES samarbetspartner, enligt artikel 17.1 i förordning (EEG) nr 1612/68, dvs.
iii) särskilda arbetsförmedlingar som anmälts till kommissionen enligt artikel 17.2 i förordning (EEG) nr 1612/68.
Europeiska samordningsbyråns roll
EURES samordningsbyrå skall särskilt
c) ansvara för den övergripande övervakningen och utvärderingen av EURES-verksamheten och vidta åtgärder för att kontrollera att den genomförs enligt bestämmelserna i förordning (EEG) nr 1612/68 och i det här beslutet.
Akronymen EURES får användas endast för verksamhet inom EURES-nätverket. Den skall illustreras med en logotyp som är definierad i ett grafiskt dokument.
Högnivågrupp för strategiska frågor
a) EURES-stadgan, enligt artikel 8.2,
d) den rapport som kommissionen vartannat år skall lämna till Europaparlamentet, rådet och Europeiska ekonomiska och sociala kommittén enligt artikel 19.3 i förordning (EEG) nr 1612/68.
EURES samordningsbyrå skall ställa sekreterartjänster till förfogande.
För att bistå högnivågruppen med utvecklingen, genomförandet och övervakningen av EURES-verksamheten skall EURES samordningsbyrå inrätta en arbetsgrupp som består av EURES-ansvariga ("EURES-managers"), som var och en företräder en EURES-medlem. EURES samordningsbyrå skall bjuda in företrädare för arbetsmarknadens parter på EU-nivå och, i lämpliga fall, företrädare för andra samarbetspartner och experter inom EURES att delta i arbetsgruppens möten.
1. EURES samordningsbyrå skall anta EURES-stadgan enligt de förfaranden som anges i artiklarna 14.2 och 15.2, artikel 22.1 a, b och c samt artikel 23 i förordning (EEG) nr 1612/68, efter samråd med den högnivågrupp för strategiska frågor som inrättas genom artikel 6 i det här beslutet.
i) arbetsförmedling, inklusive personlig vägledning och rådgivning till kunder, antingen de är arbetssökande, arbetstagare eller arbetsgivare,
b) Verksamhetsmål för EURES-systemet, de kvalitetskrav som skall gälla samt EURES medlemmars och samarbetspartners skyldigheter, vilket inbegriper
iii) utbildning och kvalifikationer som krävs av EURES-personal samt villkor och förfaringssätt för att organisera besök och uppdrag för tjänstemän,
vi) principer för övervakning och utvärdering av EURES-verksamheten.
Riktlinjer och verksamhetsplaner
2. Utifrån dessa riktlinjer skall EURES-medlemmarna lämna sina verksamhetsplaner för den period som riktlinjerna omfattar till EURES samordningsbyrå. Verksamhetsplanerna skall innehålla uppgifter om
c) formerna för övervakning och utvärdering av den planerade verksamheten, inklusive den information som skall lämnas till kommissionen varje år.
4. Kommissionen får bevilja ekonomiskt stöd för genomförandet av verksamhetsplanerna i enlighet med bestämmelserna om de relevanta budgetmedlen.
Beslut 93/569/EEG upphävs härmed. Det skall dock fortsätta att tillämpas på verksamhet för vilken en ansökan hade lämnats in innan det här beslutet trädde i kraft.
Detta beslut skall tillämpas från och med den 1 mars 2003.
Detta beslut riktar sig till medlemsstaterna.
om ändring av rådets direktiv 98/18/EG om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg
med beaktande av kommissionens förslag(1),
i enlighet med förfarandet i artikel 251 i fördraget(3), och
(2) Definitionen av fartområden är avgörande för hur direktiv 98/18/EG skall tillämpas på olika passagerarfartygsklasser. Direktivet innehåller ett förfarande för offentliggörandet av förteckningar av fartområden som visat sig vara svårt att genomföra. Det är därför nödvändigt att skapa ett praktiskt genomförbart och öppet förfarande som möjliggör en effektiv övervakning av direktivets genomförande.
(5) Med tanke på de ombyggnader av existerande ro-ro-passagerarfartyg som kan vara nödvändiga för att de skall uppfylla de särskilda stabilitetskraven, bör dessa krav införas successivt under ett antal år, så att den del av branschen som berörs får tillräcklig tid att uppfylla kraven. En tidtabell för infasning av existerande fartyg bör därför fastställas. Denna tidtabell för infasning bör inte påverka tillämpningen av de särskilda stabilitetskraven i de fartområden som omfattas av bilagorna till Stockholmsöverenskommelsen av den 28 februari 1996.
(8) Det är viktigt att vidta lämpliga åtgärder för att garantera att personer med nedsatt rörlighet under säkra former kan ta sig ombord på passagerarfartyg och höghastighetspassagerarfartyg i inrikes trafik i medlemsstaterna.
Artikel 1
"ea) ro-ro-passagerarfartyg: ett fartyg som medför fler än tolv passagerare och som har ro-ro-lastutrymmen eller lastutrymmen av särskild kategori enligt definitionen i regel II-2/A/2 i bilaga I."
2. I artikel 4 skall punkt 2 ersättas med följande:
b) offentliggöra förteckningen i en offentlig databas som är tillgänglig på den behöriga sjöfartsmyndighetens webbplats på Internet, och
"Artikel 6a
2. Ro-ro-passagerarfartyg i klasserna A och B som kölsträcks eller är på motsvarande byggnadsstadium före den 1 oktober 2004 skall uppfylla artiklarna 6, 8 och 9 i direktiv 2003/25/EG före den 1 oktober 2010 såvida de inte har tagits ur trafik den dagen eller vid en senare tidpunkt vid vilken de har uppnått en ålder av 30 år, dock senast den 1 oktober 2015.
1. Medlemsstaterna skall se till att lämpliga åtgärder vidtas, när så är praktiskt möjligt på grundval av riktlinjerna i bilaga III, för att passagerare med nedsatt rörlighet skall kunna ta sig ombord under säkra former på alla passagerarfartyg i klasserna A-D och alla höghastighetspassagerarfartyg som används för allmänna transporter och som kölsträcks eller befinner sig på motsvarande byggnadsstadium den 1 oktober 2004 eller senare.
Medlemsstaterna skall utarbeta nationella handlingsplaner för hur riktlinjerna skall tillämpas på sådana fartyg. Medlemsstaterna skall till kommissionen översända dessa handlingsplaner senast den 17 maj 2005.
Artikel 2
Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 17 november 2004. De skall genast underrätta kommissionen om detta.
Kommissionens direktiv 2003/26/EG
(Text av betydelse för EES)
med beaktande av Europaparlamentets och rådets direktiv 2000/30/EG av den 6 juni 2000 om vägkontroller av trafiksäkerheten hos nyttofordon i trafik i gemenskapen(1), särskilt artikel 8 i detta, och
(2) Området trafiksäkerhet omfattas av rådets direktiv 96/96/EG av den 20 december 1996 om tillnärmning av medlemsstaternas lagstiftning om provning av motorfordons och tillhörande släpfordons trafiksäkerhet(2), senast ändrat genom kommissionens direktiv 2001/11/EG(3), som omfattar reguljära trafiksäkerhetsprovningar, samt av direktiv 2000/30/EG, som gäller vägkontroller av trafiksäkerheten hos tunga nyttofordon. I bägge direktiven förekommer samma kommitté och förfarande för tekniska anpassningar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
2. Medlemsstaterna skall till kommissionen överlämna texterna till bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
av den 8 maj 2003
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175.1 i detta,
med beaktande av Regionkommitténs yttrande(3),
(1) Europeiska rådet enades vid mötet i Göteborg den 15 och 16 juni 2001 om en gemenskapsstrategi för hållbar utveckling som omfattar ett antal åtgärder, däribland utvecklingen av biodrivmedel.
(4) Transportsektorn, som svarar för mer än 30 % av den slutliga energiförbrukningen i gemenskapen, expanderar och trenden kommer med all säkerhet att förstärkas och koldioxidutsläppen öka; denna expansion kommer att bli procentuellt högre i kandidatländerna efter deras anslutning till Europeiska unionen.
(7) En ökad användning av biodrivmedel - utan att för den skulle utesluta användning av andra möjliga alternativa drivmedel, inbegripet motorgas (LPG) och komprimerad naturgas (CNG) för motorfordon - är ett av flera sätt för gemenskapen att minska sitt beroende av importerad energi och påverka drivmedelsmarknaden och således energiförsörjningstryggheten på medellång och lång sikt. Detta bör dock inte på något sätt minska vikten av att gemenskapslagstiftningen om bränslekvalitet, fordonsutsläpp och luftkvalitet efterlevs.
(10) Att främja användningen av biodrivmedel utgör ett steg mot en utökad användning av biomassa, vilket gör det möjligt att utveckla biodrivmedlen ytterligare i framtiden samtidigt som andra alternativ inte utesluts, särskilt inte vätgasalternativet.
(13) Nya typer av drivmedel bör uppfylla erkända tekniska standarder för att accepteras i större omfattning av konsumenter och fordonstillverkare, och därmed få spridning på marknaden. Tekniska standarder utgör också utgångspunkten för krav när det gäller utsläpp och övervakning av utsläpp. Nya drivmedelstyper kan ha svårt att uppfylla dagens tekniska standarder, som i stor utsträckning har utvecklats för konventionella fossila drivmedel. Kommissionen och standardiseringsorganen bör övervaka utvecklingen och aktivt anpassa och utveckla standarder, i synnerhet flyktighetsparametrar, så att nya typer av drivmedel kan införas med bibehållna krav på miljöprestanda.
(16) I sin resolution av den 8 juni 1998(5) godkände rådet kommissionens strategi och handlingsplan för förnybara energikällor och efterlyste särskilda åtgärder när det gäller biodrivmedel.
(19) I sin resolution av den 18 juni 1998(6) krävde Europaparlamentet att marknadsandelen för biodrivmedel skulle öka till 2 % under de kommande fem åren genom ett åtgärdspaket som bland annat omfattar skattebefrielse, finansiellt stöd till förädlingsindustrin och fastställande av en obligatorisk andel biodrivmedel för oljeföretag.
(22) Främjande av produktion och användning av biodrivmedel kan bidra till att beroendet av importerad energi och utsläppen av växthusgaser minskar. Dessutom kan biodrivmedel, i ren form eller i blandad form, i princip användas i befintliga motorfordon och användas i nuvarande bränslesystem för fordon. Blandning av biodrivmedel och fossila drivmedel kan underlätta en potentiell minskning av kostnaderna för distributionssystemet i gemenskapen.
(25) Ökad användning av biodrivmedel bör åtföljas av en noggrann analys av de miljömässiga, ekonomiska och sociala konsekvenserna för att man skall kunna avgöra huruvida det är lämpligt att öka andelen biodrivmedel i förhållande till konventionella drivmedel.
(28) Stödet för att främja användningen av biodrivmedel bör ske i överensstämmelse med försörjningstrygghet och miljömål, liksom de politiska målen och åtgärderna på området i varje medlemsstat. När så är fallet kan medlemsstaterna överväga vilka kostnadseffektiva sätt som finns för att informera om möjligheterna att använda biodrivmedel.
Artikel 1
1. I detta direktiv avses med
c) andra förnybara drivmedel: andra förnybara bränslen än biodrivmedel, som framställs från förnybara energikällor enligt definitionen i direktiv 2001/77/EG(8) och som används för transportändamål,
a) bioetanol: etanol som framställs av biomassa och/eller den biologiskt nedbrytbara delen av avfall och som skall användas som biodrivmedel.
d) biometanol: metanol som framställs av biomassa och skall användas som biodrivmedel.
g) bio-MTBE (metyltertiärbutyleter): bränsle som framställs av biometanol. Volymandelen biodrivmedel i bio-MTBE beräknas till 36 %.
j) ren vegetabilisk olja: olja framställd från oljeväxter genom pressning, extraktion eller jämförbara metoder, rå eller raffinerad men kemiskt oförändrad, då den är förenlig med motortyperna och motsvarande utsläppskrav.
b) i) Ett referensvärde för dessa mål skall vara 2 %, beräknat på energiinnehållet, av all bensin och diesel för transportändamål som släpps ut på deras marknader, senast den 31 december 2005.
a) Rena biodrivmedel eller mineraloljederivat med hög halt av biodrivmedel i enlighet med särskilda kvalitetsnormer för transporttillämpningar.
3. Medlemsstaterna skall övervaka effekterna av en användning i icke-anpassade fordon av dieselblandningar som består av mer än 5 % biodrivmedel och skall, om så krävs, vidta åtgärder för att se till att den tillämpliga gemenskapslagstiftningen om utsläppsnormer följs.
Artikel 4
- de nationella resurser som anslagits för produktion av biomassa för annan energianvändning än transport, och
I rapporterna skall avvikelser från de nationella målen i förhållande till referensvärdena i artikel 3.1 b motiveras och kan grundas på följande faktorer:
c) Nationella strategier för att anslå jämförbara resurser till produktionen av andra drivmedel som baseras på förnybara energikällor och är förenliga med målen för detta direktiv.
a) Kostnadseffektiviteten för de åtgärder som medlemsstaterna har vidtagit för att främja användningen av biodrivmedel och andra förnybara drivmedel.
d) Hållbarheten vid odling av grödor som används för att framställa biodrivmedel, särskilt markanvändning, grad av odlingsintensitet, växelbruk och användning av bekämpningsmedel.
Utifrån denna rapport skall kommissionen när det är lämpligt för Europaparlamentet och rådet lägga fram förslag om en anpassning av de mål som anges i artikel 3.1. Om rapportens slutsats blir att de vägledande målen sannolikt inte kommer att uppnås av skäl som är oberättigade och/eller inte hänför sig till nya vetenskapliga rön, skall dessa förslag ta upp nationella mål, inklusive eventuella bindande mål, i en lämplig form.
Artikel 6
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 december 2004. De skall genast underrätta kommissionen om detta.
Artikel 8
Detta direktiv riktar sig till medlemsstaterna.
om ändring av bilagorna till rådets direktiv 76/895/EEG, 86/362/EEG, 86/363/EEG och 90/642/EEG beträffande fastställande av gränsvärden för vissa bekämpningsmedelsrester i och på spannmål, livsmedel av animaliskt ursprung och vissa produkter av vegetabiliskt ursprung, inklusive frukt och grönsaker
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 86/363/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på livsmedel av animaliskt ursprung(4), senast ändrat genom direktiv 2002/79/EG(5), särskilt artikel 10 i detta,
av följande skäl:
(3) Införandet av de berörda verksamma ämnena i bilaga I till direktiv 91/414/EEG grundades på en utvärdering av de uppgifter som lämnats in om det föreslagna användningsområdet. Uppgifterna om användningen har lämnats in av vissa medlemsstater i enlighet med artikel 4.1 f i direktiv 91/414/EEG. Tillgängliga uppgifter har nu gåtts igenom, och de har befunnits vara tillräckliga för att vissa gränsvärden för bekämpningsmedelsrester skall kunna fastställas.
(6) För att berättigade förväntningar beträffande användning av befintliga lager av bekämpningsmedel skall kunna uppfyllas ges i kommissionens beslut om att inte godkänna de verksamma ämnena möjlighet till en utfasningsperiod, och därför bör beslut om gränsvärden för bekämpningsmedelsrester där ingen användning av det berörda ämnet är tillåten inom gemenskapen inte börja gälla förrän efter utgången av utfasningsperioden för det ämnet.
(9) För att konsumenterna skall få tillräckligt skydd mot exponering för bekämpningsmedelsrester till följd av otillåten användning av växtskyddsprodukter, bör de provisoriska gränsvärden som fastställs för de berörda kombinationerna av produkter/bekämpningsmedel motsvara den lägsta analytiska bestämningsgränsen.
(12) För att möjliggöra att det fastställs gränsvärden för resthalter av dikvat måste bestämmelserna i direktiv 76/895/EEG överföras till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG, och dessa bestämmelser måste strykas i direktiv 76/895/EEG. En del av dessa bestämmelser bör ändras som ett resultat av vetenskapliga och tekniska framsteg och på grund av förändrad användning och ändrade godkännanden på nationell nivå och gemenskapsnivå.
Artikel 1
De gränsvärden för bekämpningsmedelsrester som anges i bilaga I till detta direktiv skall läggas till i del A i bilaga II till direktiv 86/362/EEG.
Artikel 4
Medlemsstaterna skall senast den 30 juni 2003 sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv, med undantag för bestämmelserna för fentinhydroxid, fentinacetat och klorfenapyr, som skall sättas i kraft senast den 30 juni 2004. De skall genast underrätta kommissionen om detta.
Artikel 6
Detta direktiv riktar sig till medlemsstaterna.
om rättelse av de engelska och nederländska versionerna av förordning (EG) nr 2603/1999 om regler för övergången till den ordning för stöd till landsbygdens utveckling som föreskrivs i rådets förordning (EG) nr 1257/1999
med beaktande av rådets förordning (EG) nr 1257/1999 av den 17 maj 1999 om stöd från Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ) till utveckling av landsbygden och om ändring och upphävande av vissa förordningar(1), särskilt artikel 53.1 i denna, och
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för jordbrukets struktur och landsbygdens utveckling.
Artikel 2
av den 19 juni 2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Det företag som marknadsför ett av de snabbtest som har godkänts för TSE-övervakning har meddelat kommissionen att det har för avsikt att marknadsföra testet under ett nytt handelsnamn.
(6) Förordning (EG) nr 999/2001 bör därför ändras.
Artikel 1
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
om ändring av Europaparlamentets och rådets förordning (EG) nr 999/2001 när det gäller övervakningsprogram och specificerat riskmaterial
med beaktande av Europaparlamentets och rådets förordning (EG) nr 999/2001 av den 22 maj 2001 om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati(1), senast ändrad genom kommissionens förordning (EG) nr 1053/2003(2), särskilt artikel 23 i denna, och
(2) I förordning (EG) nr 999/2001 föreskrivs utrotningsåtgärder efter det att TSE har bekräftats hos får och getter. För att samla in epidemiologisk information bör riktade prov tas av djur som destruerats genom åtgärderna.
(5) Vetenskapliga styrkommittén har fastställt att kontaminering med vävnader från det centrala nervsystemet och tonsiller måste undvikas när tunga och kött från huvud tas ut från nötkreatur för att användas som livsmedel, för att undvika alla BSE-risker.
(8) Europaparlamentets og rådets förordning (EG) nr 1774/2002(3), ändrad genom kommissionens förordning (EG) nr 808/2003(4), innehåller bestämmelser om djur- och folkhälsa vid insamling, transport, lagring, hantering, bearbetning och användning eller bortskaffande av alla animala biprodukter som inte skall användas som livsmedel, inklusive deras avyttring och, i vissa undantagsfall, export och transitering. Särskilda bestämmelser om avlägsnande och bortskaffande av sådana produkter i bilaga XI till förordning (EG) nr 999/2001 bör därför utgå.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 16 juni 2003
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europeiska centralbankens yttrande(2),
(1) Rådets förordning (EG) nr 2223/96 av den 25 juni 1996 om det europeiska national- och regionalräkenskapssystemet(4), innehåller en referensram bestående av gemensamma standarder, definitioner, klassifikationer och bokföringsregler för sammanställande av medlemsstaternas räkenskaper för gemenskapens statistikbehov, för att sinsemellan jämförbara resultat skall erhållas från medlemsstaterna.
(4) För att den kvartalsvisa statistiken skall kunna sammanställas för euroområdet, bör den beviljade tidsfristen för sändningen av huvudaggregaten i nationalräkenskaperna minskas till 70 dagar.
(7) Kommittén för det statistiska programmet och kommittén för valuta-, finans- och betalningsbalansstatistik har rådfrågats i enlighet med artikel 3 i rådets beslut 89/382/EEG, Euratom(5) och rådets beslut 91/115/EEG(6).
Bilaga B till förordning (EG) nr 2223/96 ändras enligt följande:
b) Texten till tabell 1, "Huvudaggregat - kvartalsvis och årlig redovisning" skall ersättas med texten i bilaga II.
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
om ändring av förordning (EG) nr 1488/2001 om tillämpningsföreskrifter för rådets förordning (EG) nr 3448/93 när det gäller att hänföra vissa kvantiteter av vissa basprodukter enligt bilaga I till Fördraget om upprättandet av Europeiska gemenskapen till förfarandet för aktiv förädling utan förhandskontroll av de ekonomiska kraven
av följande skäl:
(3) De åtgärder som föreskrivs i denna förordning står i överensstämmelse med yttrandet från Kommittén för övergripande frågor rörande handel med bearbetade jordbruksprodukter som inte omfattas av bilaga I till fördraget.
Förordning (EG) nr 1488/2001 ändras enligt följande:
2. I artikel 22 skall det andra stycket ersättas med följande:"Om de bidrag som skall betalas ut beräknas bli större än de tillgängliga ekonomiska medlen, skall den återstående kvantiteten för varje basprodukt fastställas i enlighet med artikel 11.1 i förordning (EG) nr 3448/93 med beaktande av redan licensierade kvantiteter och av de icke-utnyttjade kvantiteter som kommissionen informerats om i enlighet med artikel 25 i denna förordning. Denna kvantitet skall offentliggöras i Europeiska unionens officiella tidning en andra gång senast den 31 januari varje år och en tredje gång senast den 31 maj varje år."
Utfärdande av AF-licenser i nödfall
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Uppbyggnaden av och koderna i CPV bör uppdateras för att ta hänsyn till de särskilda behov som medlemsstaterna och användarna av CPV gett uttryck för samt för att rätta sakfel i de olika språkversionerna.
(6) Berörda parter och CPV-användare har bidragit med förslag till förbättring av CPV.
(9) I och med att kommissionens förordning (EG) nr 204/2002 av den 19 december 2001 om ändring av rådets förordning (EEG) nr 3696/93 om den statistiska indelningen av produkter efter näringsgren (CPA) inom Europeiska ekonomiska gemenskapen(3) trädde i kraft, har konverteringstabellen mellan CPV och CPA 96 i bilaga II till förordning (EG) nr 2195/2002 blivit inaktuell.
(12) Förordning (EG) nr 2195/2002 bör därför ändras.
Artikel 1
Bilaga II skall ersättas med texten i bilaga II till denna förordning.
Bilaga V skall ändras i enlighet med bilaga V till denna förordning.
Kommissionens förordning (EG) nr 317/2004
(Text av betydelse för EES)
med beaktande av Europaparlamentets och rådets förordning (EG) nr 2150/2002 av den 25 november 2002 om avfallsstatistik(1), särskilt artikel 4.1 i denna,
med beaktande av Luxemburgs begäran av den 25 juni 2003, och
(2) Efter begäran bör sådana undantag beviljas Österrike, Frankrike och Luxemburg.
Artikel 1
b) Frankrike beviljas undantag för redovisning av resultat avseende avsnitt 8.1.1, posterna 1 (jordbruk, jakt och skogsbruk), 2 (fiske) och 16 (tjänster) i bilaga I samt de som avser avsnitt 8.2 i bilaga II.
Efter övergångsperiodens utgång skall Österrike, Frankrike och Luxemburg redovisa uppgifter från referensåret 2006.
