RÅDETS FÖRSTA DIREKTIV av den 23 juli 1962 om fastställande av vissa gemensamma regler för internationella transporter (yrkesmässiga godstransporter på väg)
med beaktande av Europaparlamentets yttrande, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. De typer av transporter som är förtecknade i bilaga 1 skall vara undantagna från kvoterings- eller tillståndssystem.
Artikel 2
Detta direktiv skall inte påverka de villkor som en medlemsstat uppställer för sina egna medborgare för att bedriva sådan verksamhet som avses i detta direktiv.
KOMMISSIONENS FÖRORDNING (EEG) nr 1397/68 av den 6 september 1968 om ändring av förordning nr 474/67/EEG om förutfastställelse av exportbidraget för ris och brutet ris
med beaktande av rådets förordning nr 359/67/EEG av den 25 juli 1967 om den gemensamma organisationen av marknaden för ris(1), särskilt artikel 17.6 i denna, och
Det är därför nödvändigt att ändra förordning nr 474/67/EEG.
Artikel 1
- med tillägg av ett belopp som inte överstiger skillnaden mellan cif-priset och cif-priset för terminsköp, när det förstnämnda överstiger det sistnämnda med mer än 0,025 räkneenheter per 100 kg.
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
- från och med den 1 september 1972 för fordon som tas i bruk för första gången.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 3
Artikel 4
De ändringar som är nödvändiga för att anpassa kraven i bilaga 1 7 till tekniska framsteg skall beslutas enligt det förfarande som fastslås i artikel 13 i rådets direktiv av den 6 februari 1970 om typgodkännande av motorfordon och släpvagnar till dessa fordon.
2. Medlemsstaterna skall se till att till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
RÅDETS DIREKTIV av den 24 juli 1973 om åtgärder för att dämpa verkningarna av svårigheter vid försörjningen med råolja eller petroleumprodukter (73/238/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: Fastställandet av en gemensam energipolitik tillhör de mål som gemenskaperna har ställt upp.
Medlemsstaterna bör därför ges de nödvändiga befogenheterna för att, om så erfordras, omedelbart kunna vidta lämpliga åtgärder i enlighet med bestämmelserna i fördraget, särskilt artikel 103 i detta.
Det är nödvändigt att varje medlemsstat upprättar en plan som kan följas vid svårigheter i försörjningen med råolja eller petroleumprodukter.
Artikel 3
Medlemsstaterna skall senast den 30 juni 1974 sätta i kraft de rättsliga och administrativa bestämmelser som är nödvändiga för att följa detta direktiv.
RÅDETS FÖRORDNING (EKSG, EEG, Euratom) nr 559/73 av den 26 februari 1973 om ändring av rådets förordning (EEG, Euratom, EKSG) nr 260/68 om villkoren för och förfarandet vid skatt till Europeiska gemenskaperna
med beaktande av protokollet om immunitet och privilegier för Europeiska gemenskaperna, särskilt artikel 13 i detta,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
I artikel 3.3 a första strecksatsen skall "familjeförsörjartillägg" ersättas med "hushållstillägg".
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(1),
Dessa krav skiljer sig åt i de olika medlemsstaterna. Det är därför nödvändigt att alla medlemsstater antar samma krav, antingen som tillägg till eller i stället för sina nuvarande bestämmelser, särskilt för att det förfarande med EEG-typgodkännande, som behandlats i rådets direktiv av den 6 februari 1970(3) om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon, skall kunna tillämpas på alla fordonstyper.
När det gäller tekniska krav är det lämpligt att huvudsakligen tillämpa de som antagits av FNs ekonomiska kommission för Europa i reglemente nr 21 ("Enhetliga krav om godkännande av fordon med avseende på inredningar i dessa"), vilka återges i en bilaga till överenskommelsen av den 20 mars 1958 om antagande av enhetliga villkor för godkännande och ömsesidigt erkännande av utrustning och delar för motorfordon.
I detta direktiv avses med fordon varje motorfordon i kategori M1 (definieras i bilaga 1 till direktivet av den 6 februari 1970) som är avsett att användas på väg, har minst fyra hjul och är konstruerat för en högsta hastighet som överstiger 25 km/tim.
- passagerarutrymmets inre delar frånsett inre backspeglar, - manöverorganens utformning,
om dessa uppfyller kraven i bilagorna.
- manöverorganens utformning,
om dessa inredningsdetaljer uppfyller kraven i bilagorna.
Artikel 5
1. Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv inom 18 månader från dagen för anmälan och skall genast underrätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: I förordning (EEG) nr 922/72(2), ändrad genom förordning (EEG) nr 884/73(3), fastställer rådet allmänna tillämpningsföreskrifter för stöd till silkesmaskar för odlingsåren 1972/1973 och 1973/1974. Erfarenheten har visat att det är lämpligt att fortsätta att tillämpa förordningen under kommande odlingsår.
I artikel 1 i förordning (EEG) nr 922/72 skall orden "för odlingsåren 1972/1973 och 1973/1974" utgå.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av kommissionens förslag,
med beaktande av följande: Direktiv nr 64/221/EEG (3) samordnade särskilda åtgärder som gäller utländska medborgares rörlighet och bosättning och som är berättigade med hänsyn till allmän ordning, säkerhet eller hälsa, och direktiv nr 75/34/EEG (4) fastställde enligt vilka villkor medborgare i en medlemsstat skall ha rätt att stanna kvar inom en annan medlemsstats territorium efter att ha varit verksamma där som egna företagare.
Artikel 1
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
Med hänsyn till det tekniska kunnande som för närvarande har uppnåtts skall tillämpningsområdet för detta direktiv begränsas till aerosolbehållare av metall, glas och plast.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Den som svarar för att aerosolbehållare släpps ut på marknaden skall förse dessa med symbolen "3" (omvänt epsilon) som bevis för att de uppfyller kraven i detta direktiv och dess bilaga.
Artikel 6
Artikel 7
3. a) Kommissionen skall själv anta förslaget, om det har tillstyrkts av kommittén.
Artikel 8
c) Kodbeteckningar som gör det möjligt att identifiera varuparti.
2. Medlemsstaterna kan ställa som villkor för försäljning inom sitt territorium att nationalspråket eller -språken används för förpackningstexten.
Artikel 10
3. Om kommissionen anser att direktivet behöver bearbetas i tekniskt avseende, skall sådana bearbetningar godkännas av antingen kommissionen eller rådet i enlighet med det förfarande som anges i artikel 7. Om så är fallet kan den medlemsstat som infört säkerhetsåtgärder behålla dessa, tills de nya bestämmelserna trätt i kraft.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
RÅDETS DIREKTIV av den 26 juni 1975 om ändring av direktiven 66/400/EEG, 66/401/EEG, 66/402/EEG, 66/403/EEG och 69/208/EEG om saluföring av betutsäde, utsäde av foderväxter, utsäde av stråsäd, utsädespotatis och utsäde av olje- och spånadsväxter (75/444/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: Vissa direktiv om saluföring av utsäde bör ändras av nedan angivna skäl.
Det är i detta sammanhang lämpligt att, å ena sidan, underlätta saluföring och plombering av sådana små förpackningar och, å andra sidan, göra tillräcklig äkthetskontroll av utsädet obligatorisk.
Det är också nödvändigt att göra vissa ändringar av det sätt på vilket utsädeskvantiteterna anges.
Rådets direktiv 66/400/EEG(3) av den 14 juni 1966 om saluföring av betutsäde, senast ändrat genom direktiv 73/438/EEG(4) skall ändras på följande sätt: 1. Följande stycke skall läggas till artikel 2.1:
1. Medlemsstaterna skall kräva att förpackningar med basutsäde och certifikatutsäde, förutom då utsäde av den sistnämnda kategorin förpackas i EEG-småförpackningar, skall plomberas officiellt på sådant sätt att plomberingen skadas och inte kan anbringas på nytt när förpackningen öppnats.
4. Medlemsstaterna får anta bestämmelser om undantag från punkt 1 och 2 för småförpackningar med basutsäde."
5. Texten i artikel 11.2 b skall ersättas med följande:
Obligatoriska uppgifter 1. "EEG-småförpackning".
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 42 och 43 i detta,
med beaktande av följande. De grundläggande bestämmelserna om organisationen av marknaden för fjäderfäkött har ändrats ett flertal gånger sedan de antogs. Eftersom bestämmelserna är många och komplicerade och dessutom återfinns i ett antal olika nummer av Europeiska gemenskapernas officiella tidning, är de svåra att tillämpa och saknar följaktligen den klarhet som bör vara ett väsentligt drag i all lagstiftning. De bör därför sammanföras i en enda text.
Förverkligandet av en enhetlig marknad för fjäderfäkött inbegriper införandet av ett enhetligt system för handeln över gemenskapens yttre gränser, innefattande importavgifter och exportbidrag.
Gemenskapens deltagande i den internationella handeln med fjäderfäkött skulle säkras av möjligheten att vid export till tredje land bevilja ett exportbidrag som motsvarar skillnaden mellan priserna inom gemenskapen och priserna på världsmarknaden. För att garantera gemenskapens exportörer ett visst mått av trygghet med avseende på exportbidragens stabilitet, bör det göras möjligt att fastställa exportbidraget för fjäderfäkött på förhand.
Den gemensamma organisationen av marknaden för fjäderfäkött skall på lämpligt sätt och samtidigt ta hänsyn till de mål som fastställs i artikel 39 och artikel 110 i fördraget.
2. I denna förordning avses med: a) levande fjäderfä: levande höns, ankor, gäss, kalkoner och pärlhöns med en vikt på över 185 gram.
d) härledda produkter: 1. produkter enligt punkt 1 a utom kycklingar.
4. produkter enligt punkt 1 c,
e) kvartal: tremånadersperiod som börjar den 1 februari, den 1 maj, den 1 augusti eller den 1 november.
- Åtgärder för att möjliggöra kort- och långsiktiga prognoser på grundval av de produktionsmedel som används.
2. Handelsnormer - skall antas för en eller flera av de produkter som anges i artikel 1.1 b,
På förslag av kommissionen skall rådet med kvalificerad majoritet fastställa normerna och deras användningsområde samt allmänna tillämpningsföreskrifter för dem.
Artikel 4
Världsmarknadspriserna på foderspannmål skall fastställas kvartalsvis på basis av priserna på sådan spannmål under de sex månader som föregår det kvartal under vilket nämnda del beräknas.
3. På förslag av kommissionen skall rådet med kvalificerad majoritet - fastställa den kvantitet foderspannmål, differentierad med hänsyn till art av fjäderfä, som åtgår till att producera 1 kg slaktat fjäderfä och den kvantitet foderspannmål som åtgår till att producera en kyckling, samt procentsatserna av de olika slag av foderspannmål som ingår i dessa kvantiteter,
1. För de produkter som anges i artikel 1.2 d skall importavgiften härledas från importavgiften för slaktat fjäderfä, på basis av viktförhållandet mellan dessa olika produkter och slaktat fjäderfä och, vid behov, det genomsnittliga förhållandet mellan deras marknadsvärden.
Artikel 6
Artikel 7
b) Ett standardbelopp som representerar övriga foderkostnader och omkostnader för produktion och försäljning, differentierad med hänsyn till art av fjäderfä.
3. Slusspriset på kycklingar skall beräknas på samma sätt som slusspriset på slaktat fjäderfä. Dock skall världsmarknadspriset på kvantiteten foderspannmål vara priset på den kvantitet som åtgår till att i tredje land producera en kyckling och standardbeloppet skall vara det belopp som representerar övriga foderkostnader och omkostnader för produktion och försäljning för en kyckling. Mängden foderspannmål och standardbeloppet skall inte variera beroende på art.
Artikel 8
3. Anbudspriset fritt gränsen skall fastställas för all import från tredje land.
Då tilläggsavgifter krävs, skall dessa fastställas i enlighet med samma förfarande.
2. Exportbidraget skall vara detsamma för hela gemenskapen. Det får variera beroende på användning och bestämmande.
På förslag av kommissionen skall rådet med kvalificerad majoritet fastställa allmänna bestämmelser om beviljande av och förutfastställelse av exportbidrag och kriterier för fastställande av dessa belopp.
Artikel 10
1. De allmänna bestämmelserna om tolkningen av Gemensamma tulltaxan och de särskilda tillämpningsföreskrifterna skall gälla tullklassificeringen av produkter som omfattas av denna förordning. Tullnomenklaturen som skapas genom tillämpningen av denna förordning skall ingå som del i Gemensamma tulltaxan.
- Tillämpning av någon kvantitativ restriktion eller åtgärd med motsvarande verkan. Varje åtgärd som begränsar utfärdandet av import- eller exportlicenser till en angiven personkategori skall betraktas som en åtgärd som har samma verkan som en kvantitativ restriktion.
På förslag av kommissionen skall rådet med kvalificerad majoritet fastställa närmare tillämpningsföreskrifter för denna punkt samt närmare ange under vilka omständigheter och inom vilka gränser medlemsstaterna får vidta skyddsåtgärder.
Artikel 13
För att ta hänsyn till eventuella begränsningar av den fria omsättningen till följd av åtgärder för att förhindra spridning av djursjukdomar, får extraordinära åtgärder för att stödja marknader som påverkas av sådana begränsningar vidtas i enlighet med det förfarande som föreskrivs i artikel 17. Sådana åtgärder får endast vidtas i den mån och under den tid som det är absolut nödvändigt för att stödja denna marknad.
Artikel 16
Artikel 17
3. Kommissionen skall besluta med omedelbar verkan. Om beslutet inte är förenligt med kommitténs yttrande skall kommissionen emellertid genast underrätta rådet. I sådana fall får kommissionen uppskjuta verkställandet av de beslutade åtgärderna under en tid som inte överstiger en månad från dagen då rådet underrättats.
Kommittén får överväga varje annan fråga som dess ordförande hänskjuter till kommittén på eget initiativ eller på begäran av en medlemsstats företrädare.
Artikel 20
Om Italien åberopar bestämmelserna i artikel 23 i rådets förordning (EEG) nr 2727/75(4) av den 29 oktober 1975 om den gemensamma organisationen av marknaden för spannmål, skall rådet, på förslag av kommissionen, med kvalificerad majoritet besluta om de åtgärder som krävs för att undvika en snedvridning av konkurrensen.
2. Alla hänvisningar till den förordning som upphävs i punkt 1 skall betraktas som hänvisningar till den här förordningen.
Denna förordning träder i kraft den 1 november 1975.
med beaktande av kommissionens förslag,
med beaktande av följande: De tekniska krav som motorfordon måste uppfylla enligt nationell lagstiftning gäller bl.a. föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Ingen medlemsstat får vägra att registrera ett fordon eller förbjuda att det säljs, tas i bruk eller används av skäl som hänför sig till de föreskrivna skyltarna och märkningarna eller deras placering och fastsättningsmetod om de uppfyller kraven i bilagan till detta direktiv.
Artikel 5
RÅDETS DIREKTIV av den 8 december 1975 om kvaliteten på badvatten (76/160/EEG)
med beaktande av kommissionens förslag,
med beaktande av följande: För att skydda miljön och människors hälsa är det nödvändigt att minska föroreningen av badvatten och att skydda sådant vatten mot ytterligare försämring.
Enligt Europeiska gemenskapernas åtgärdsprogram för miljön(3) skall gemensamma kvalitetsmål uppställas med avseende på miljökvaliteten, bl.a. angivande av parametervärden för vatten, inklusive badvatten.
För att uppnå ett visst mått av flexibilitet vid tillämpningen av detta direktiv måste medlemsstaterna ha befogenhet att föreskriva undantag. Sådana undantag får emellertid inte bortse från krav som är väsentliga för skyddet av människors hälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
b) "badplats": varje plats där badvatten finns,
Fysikaliska, kemiska och mikrobiologiska parametrar som gäller för badvatten anges i bilagan, som utgör en integrerad del av detta direktiv.
Artikel 4
- i 90 % av proverna i alla andra fall med undantag av parametrarna för "kolibakterier, totalt" och "fekala kolibakterier" där procentsatsen får vara 80 %,
Artikel 6
Bestämmelserna i detta direktiv får åsidosättas a) i fråga om vissa parametrar märkta (0) i bilagan vid exceptionella meteorologiska eller geografiska förhållanden,
De undantag som föreskrivs i denna artikel får inte i något fall medföra att krav som är väsentliga för att skydda människors hälsa åsidosätts.
Sådana ändringar som är nödvändiga för att anpassa detta direktiv till den tekniska utvecklingen skall avse - analysmetoderna,
Artikel 10
b) Om förslaget inte är förenligt med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv inom två år efter dagen för anmälan. De skall genast underrätta kommissionen om detta.
Medlemsstaterna skall fyra år efter anmälan av detta direktiv och därefter regelbundet till kommissionen överlämna en utförlig rapport om sitt badvatten och dess mest betydelsefulla egenskaper.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(2), och
Rådets direktiv 71/316/EEG av den 26 juli 1971 om tillnärmning av medlemsstaternas lagstiftning om gemensamma föreskrifter för både mätdon och metrologiska kontrollmetoder(3) har fastställt förfaranden för EEG-typgodkännande och första EEG-verifikation. Enligt det direktivet är det nödvändigt att fastställa de tekniska krav som skall gälla för konstruktion och funktion av alkoholmätare och alkoholaerometrar för att de efter föreskriven kontroll och märkning fritt skall få importeras, marknadsföras och användas.
Artikel 1
Artikel 3
Bestämmelserna skall börja tillämpas senast den 1 januari 1980.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 75 i detta,
med beaktande av Europaparlamentets yttrande(),
Vid fastställande av miniminivån för sådan utbildning bör man särskilt ta hänsyn till de olika förutsättningar som råder för gods- respektive persontransporter på väg.
1. Den som innehar gällande nationellt körkort och som har genomgått yrkesutbildning som omfattar åtminstone de ämnen som är uppräknade i bilagan till detta direktiv, skall anses ha uppfyllt minimikravet på utbildning för förare av fordon avsedda för godstransporter på väg enligt artikel 5.1 b andra strecksatsen i förordning (EEG) nr 543/69 eller för förare av fordon avsedda för persontransporter på väg enligt punkt 2 c av nämnda artikel.
Artikel 2
Artikel 3
Artikel 4
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Avtalets text ingår i bilaga till denna förordning.
Artikel 3
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande (1),
För att aktieägarna och borgenärerna skall kunna garanteras ett minimum av likvärdigt skydd är det särskilt viktigt att samordna de nationella bestämmelserna om att bilda ett aktiebolag samt om att bevara, öka och sätta ned dess kapital.
Med hänsyn till ändamålet med artikel 54.3 i fördraget måste medlemsstaternas lagstiftning om ökning och nedsättning av kapitalet säkerställa att de principer beaktas och harmoniseras som syftar till en lika behandling av aktieägare med samma ställning och till ett skydd för borgenärer med fordringar som har uppkommit före en kapitalnedsättning,
1. De samordningsåtgärder som detta direktiv föreskriver skall vidtas i fråga om bestämmelserna i medlemsstaternas lagar eller andra författningar om följande bolagsformer: - I Belgien: la société anonyme/de naamloze vennootschap.
2. Medlemsstaterna behöver inte tillämpa detta direktiv på förvaltningsbolag med rörligt kapital eller på kooperativa företag som är organiserade i någon av de i punkt 1 angivna bolagsformerna. Om lagstiftningen i en medlemsstat utnyttjar denna möjlighet, skall den föreskriva att dessa bolag skall ta in orden "förvaltningsbolag med rörligt kapital" eller "kooperativt företag" i samtliga de handlingar som nämns i artikel 4 i direktiv 68/151/EEG.
- vars bolagsordning anger att bolaget inom gränserna för ett minimikapital och ett maximikapital alltid får ge ut, lösa in eller avyttra sina aktier.
b) föremålet för bolagets verksamhet;
d) bestämmelser som anger antalet ledamöter och hur dessa skall utses i de organ som företräder bolaget mot tredje man och svarar för förvaltning, ledning, övervakning eller kontroll av bolaget samt bestämmelser om kompetensfördelningen mellan organen, allt i den mån föreskrifter inte finns i lag eller annan författning;
Minst följande uppgifter skall finnas antingen i bolagsordningen eller stiftelseurkunden eller i en särskild handling som skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG: a) bolagets säte;
d) i förekommande fall de särskilda villkor som begränsar aktiernas överlåtbarhet;
g) hur stor del av det tecknade kapitalet som är betalt då bolaget bildas eller då det får tillstånd att börja sin verksamhet;
j) åtminstone uppskattningsvis summan av alla kostnader som har uppkommit för bolaget eller påförts detta med anledning av bolagsbildningen och, i förekommande fall, innan bolaget får tillstånd att börja sin verksamhet;
1. Om enligt lagstiftningen i en medlemsstat ett bolag inte får börja sin verksamhet utan tillstånd, skall denna lagstiftning även innehålla bestämmelser om ansvaret för förbindelser som har ingåtts av bolaget eller för dettas räkning innan ansökningen om tillstånd beviljades eller avslogs.
1. Om lagstiftningen i en medlemsstat kräver att ett bolag skall bildas av flera bolagsmän, medför inte det förhållandet att därefter alla aktierna förenas på en hand eller antalet bolagsmän sjunker under det i lagstiftningen föreskrivna minimiantalet att bolaget utan vidare upplöses.
Artikel 6
3. Med hänsyn till den ekonomiska och monetära utvecklingen inom gemenskapen och till tendensen att tillåta endast större och medelstora företag att välja de i artikel 1.1 angivna bolagsformerna, skall rådet vart femte år på förslag av kommissionen överväga och vid behov ändra de i denna artikel i europeiska beräkningsenheter uttryckta beloppen.
Artikel 8
Artikel 9
Artikel 10
3. Sakkunnigutlåtandet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
c) de bolag som lämnar apportegendomen har reserver som enligt lag eller bolagsordning inte får delas ut och som uppgår till minst det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet hos de aktier som ges ut mot apportegendom;
f) de bolag som lämnar apportegendomen för över ett belopp som motsvarar det vid c angivna värdet till en reserv som får delas ut först tre år efter det att det mottagande bolagets årsredovisning har offentliggjorts för det räkenskapsår under vilket apportegendomen lämnades eller, i förekommande fall, först vid den senare tidpunkt då alla fordringar som omfattas av det vid d angivna ansvaret och som görs gällande under den nu angivna treårsperioden har tillgodosetts.
Medlemsstaterna får föreskriva att dessa bestämmelser även skall tillämpas när tillgångarna tillhör en aktieägare eller någon annan.
Aktieägarna får inte befrias från sin skyldighet att betala aktierna i andra fall än som kan följa av bestämmelserna om nedsättning av det tecknade kapitalet.
Artikel 14
1. a) Med undantag för det fallet att det tecknade kapitalet sätts ned får någon utdelning inte ske till aktieägarna, om enligt bolagets årsredovisning nettotillgångarna på bokslutsdagen för det senaste räkenskapsåret understiger eller till följd av utdelningen skulle komma att understiga det tecknade kapitalet och de reserver som enligt lag eller bolagsordning inte får delas ut.
d) Med "utdelning" avses i a och c särskilt utbetalning av vinst eller ränta som hänför sig till aktierna.
3. Punkterna 1 och 2 inkräktar inte på medlemsstaternas bestämmelser om ökning av det tecknade kapitalet genom överföring av reserver till detta.
- som vänder sig till allmänheten för att placera sina egna aktier.
c) skall denna föreskriva att ett nu avsett bolag, som delar ut medel till aktieägarna när nettotillgångarna understiger det i punkt 1 a angivna beloppet, skall upplysa om utdelningen i en not till årsredovisningen.
Artikel 17
Artikel 18
3. Aktier som har tecknats i strid med denna artikel skall betalas av de i artikel 3 i angivna personerna eller bolagen eller, vid ökning av det tecknade kapitalet, av medlemmarna i styrelsen eller direktionen.
1. Om lagstiftningen i en medlemsstat tillåter att ett bolag förvärvar egna aktier, antingen direkt eller genom någon som handlar i eget namn men för bolagets räkning, skall enligt den lagstiftningen minst följande villkor gälla för ett sådant förvärv: a) Tillstånd till förvärvet skall lämnas av bolagsstämman som skall ange de närmare förutsättningarna för detta och särskilt det högsta antal aktier som får förvärvas, den tid inom vilken tillståndet gäller, vilken tid inte får överstiga 18 månader, samt vid förvärv mot vederlag det lägsta och högsta vederlaget. Medlemmarna av styrelsen eller direktionen skall se till att de vid b, c och d angivna villkoren iakttas när förvärvet äger rum.
d) Förvärvet får endast omfatta helt betalda aktier.
Artikel 20
c) helt betalda aktier som förvärvas utan vederlag eller som utgör inköpsprovision för banker och andra finansinstitut;
f) aktier som förvärvas för att hålla minoritetsaktieägare i närstående bolag skadeslösa;
2. Aktier som har förvärvats enligt 1 b-g skall dock avyttras inom högst tre år, med mindre det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet av de förvärvade aktierna inräknat de aktier som bolaget har förvärvat genom någon som handlat i eget namn men för bolagets räkning, inte överstiger tio procent av det tecknade kapitalet.
Aktier som har förvärvats i strid med artiklarna 19 och 20 skall avyttras inom ett år från förvärvet. Om de inte avyttras inom denna tid tillämpas artikel 20.3.
a) av de rättigheter som är knutna till aktier får rösträtt aldrig utövas för de egna aktierna; b) om dessa aktier tas upp som en tillgång i balansräkningen skall ett motsvarande belopp, som bolaget inte får förfoga över, tas upp som en reserv bland skulderna;
c) vid förvärv eller avyttring mot vederlag, uppgift om vederlaget för aktierna;
1. Ett bolag får inte ge förskott, lämna lån eller ställa säkerhet i syfte att tredje man skall förvärva aktier i bolaget.
Artikel 24
Artikel 25
3. Om det finns flera slag av aktier, skall bolagsstämmans beslut om kapitalökning enligt punkt 1 eller om bemyndigande att öka kapitalet enligt punkt 2 bli föremål för en särskild omröstning minst för varje kategori av aktieägare vilkas rätt berörs av beslutet.
Om aktier ges ut mot vederlag som ett led i ökningen av det tecknade kapitalet, skall de betalas med minst 25 procent av aktiernas nominella värde eller, i avsaknad av sådant värde, av det bokförda parivärdet. Om en överkurs fastställs, skall denna betalas helt.
3. Medlemsstaterna behöver inte tillämpa punkt 2, om ökningen av det tecknade kapitalet sker för att genomföra en fusion eller ett offentligt erbjudande om köp eller byte och i syfte att ersätta aktieägarna i ett bolag som upplöses genom fusionen eller är föremål för det offentliga erbjudandet om köp eller byte.
Om en kapitalökning inte fulltecknas, skall kapitalet ökas med det tecknade beloppet endast om emissionsvillkoren uttryckligen har föreskrivit det.
2. Medlemsstaterna a) behöver inte tillämpa punkt 1 på aktier med en begränsad rätt till utdelning enligt artikel 15 och/eller vid utskiftning av bolagets förmögenhet i samband med likvidation; eller
4. Företrädesrätten får inte begränsas eller upphävas i bolagsordningen eller stiftelseurkunden. Detta får däremot ske genom ett beslut av bolagsstämman. Direktionen eller styrelsen skall i så fall lämna bolagsstämman en skriftlig redogörelse som anger skälen för att begränsa eller upphäva företrädesrätten och grunderna för den föreslagna emissionskursen. Bolagsstämmans beslut skall fattas enligt bestämmelserna i artikel 40 om beslutförhet och majoritet. Beslutet skall offentliggöras enligt varje medlemsstats lagstiftning i överensstämmelse med artikel 3 i direktiv 68/151/EEG.
7. Företrädesrätten anses inte utesluten enligt punkt 4 eller 5, om aktierna på grund av beslutet om ökning av det tecknade kapitalet ges ut till banker eller andra finansinstitut för att dessa skall erbjuda aktierna till bolagets aktieägare enligt punkterna 1 och 3.
Om det finns flera slag av aktier, skall bolagsstämmans beslut om nedsättning av det tecknade kapitalet bli föremål för en särskild omröstning minst för varje kategori av aktieägare vilkas rätt berörs av beslutet.
2. Medlemsstaternas lagstiftning skall vidare minst föreskriva att nedsättningen inte gäller eller att någon utbetalning inte får ske till förmån för aktieägarna, förrän borgenärerna har fått gottgörelse eller en domstol har beslutat att deras framställning därom inte behöver efterkommas.
1. Medlemsstaterna behöver inte tillämpa artikel 32 vid en nedsättning av det tecknade kapitalet som sker för att täcka en inträffad förlust eller för att föra över vissa belopp till en reserv, om reserven därefter inte överstiger tio procent av det nedsatta tecknade kapitalet. Utom vid nedsättning av det tecknade kapitalet får denna reserv inte delas ut till aktieägarna; den får endast användas för att täcka en inträffad förlust eller för att öka det tecknade kapitalet genom överföring av reserver, i den mån medlemsstaterna tillåter en sådan åtgärd.
Det tecknade kapitalet får inte sättas ned under det minimikapital som har fastställts i överensstämmelse med artikel 6. Medlemsstaterna får dock tillåta en sådan nedsättning, om de även föreskriver att beslutet om nedsättning får verkställas först sedan det tecknade kapitalet har ökats till minst det fastställda minimikapitalet.
b) Endast belopp som får delas ut enligt artikel 15.1 får användas för inlösen.
1. Om lagstiftningen i en medlemsstat tillåter bolagen att sätta ned det tecknade kapitalet genom att tvångsvis dra in aktier, skall lagstiftningen minst kräva att följande villkor är uppfyllda:
d) Artikel 32 tillämpas utom i fråga om helt betalda aktier som ställs till bolagets förfogande utan vederlag eller som dras in med utnyttjande av medel som får delas ut enligt artikel 15.1; i dessa fall skall ett belopp som motsvarar det nominella värdet eller, i avsaknad av sådant värde, det bokförda parivärdet för samtliga indragna aktier föras över till en reserv. Utom vid nedsättning av det tecknade kapitalet får denna reserv inte delas ut till aktieägarna; den får endast användas för att täcka en inträffad förlust eller för att öka det tecknade kapitalet genom överföring av reserver, i den mån medlemsstaterna tillåter en sådan åtgärd.
Artikel 37
3. Artiklarna 31, 33 och 40 tillämpas inte i de fall som avses i punkt 1.
Artikel 39
c) villkoren och sättet för återköpet skall vara bestämda i bolagsordningen eller stiftelseurkunden;
f) punkt e tillämpas inte, om återköpet har skett med intäkter från en nyemission som har ägt rum i och för återköpet;
Artikel 40
Artikel 41
Artikel 42
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som behövs för att följa detta direktiv inom två år efter dagen för anmälan. De skall genast underrätta kommissionen om detta.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 43 och 100 i detta,
med beaktande av följande: Produktionen av nötkreatur upptar en mycket viktig plats i gemenskapens jordbruk. Tillfredsställande resultat är till stor del beroende av användningen av renrasiga avelsdjur.
Medlemsstaterna måste få möjlighet att kräva att härstamningsintyg som är utformade enligt ett gemenskapsförfarande skall uppvisas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- som förs av en avelsorganisation eller avelsförening som är officiellt godkänd av den medlemsstat där organisationen eller föreningen bildats, och
Medlemsstaterna skall se till att följande inte får förbjudas, begränsas eller hindras på avelsmässiga grunder: - Handel med renrasiga avelsdjur av nötkreatur inom gemenskapen.
- Godkännande av organisationer eller föreningar som för stamböcker enligt artikel 6.
Rådet skall på förslag från kommissionen före den 1 juli 1980 anta gemenskapsbestämmelser för godkännande av renrasiga avelsdjur av nötkreatur för avelsändamål.
Avelsorganisationer eller avelsföreningar som är officiellt godkända av en medlemsstat får inte motsätta sig att renrasiga avelsdjur av nötkreatur från andra medlemsstater införs i deras stamböcker, förutsatt att djuren uppfyller de krav som fastställs enligt artikel 6.
Artikel 6
- Villkor för upprättande av stamböcker.
2. Till dess att bestämmelserna i punkt 1 första, andra och tredje strecksatserna träder i kraft a) skall de officiella kontroller som avses i punkt 1 första strecksatsen och som utförs i varje medlemsstat, samt de stamböcker som för närvarande finns, erkännas av övriga medlemsstater,
Artikel 7
Artikel 8
3. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med en majoritet av 41 röster.
Artikel 9
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(1), senast ändrad genom förordning (EEG) nr 1707/73(2),
med beaktande av följande: I artikel 2 i kommissionens förordning (EEG) nr 616/72 av den 27 mars 1972 om tillämpningsföreskrifter för exportbidrag och avgifter på olivolja(6), senast ändrad genom förordning (EEG) nr 503/76(7), föreskrivs att den rätt att importera med befrielse från avgift som anges i artikel 9 i förordning nr 171/67/EEG, skall beviljas för de kvaliteter av olivolja för vilka det finns ett kontantbidrag.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"Den rätt till avgiftsfri import som anges i artikel 9.1 i förordning nr 171/67/EEG, skall vara beroende av att exporten omfattar kvaliteter på olivoljan och i förekommande fall presentationsformer, för vilka ett kontantbidrag gäller den dag då ansökan om detta tillstånd lämnas in."
KOMMISSIONENS FÖRSTA DIREKTIV av den 18 april 1978 om ändring av bilagorna till direktiv 66/402/EEG om saluföring av utsäde av stråsäd (78/387/EEG)
med beaktande av rådets direktiv 66/402/EEG av den 14 juni 1966 om saluföring av utsäde av stråsäd(1), senast ändrat genom rådets direktiv 78/55/EEG(2), särskilt artikel 21a i detta, och
I syfte att förbättra kvaliteten på utsäde bör bestämmelser antas om villkoren för föregående skörd.
För att uppfylla villkoren för officiella undersökningar av utsäde som utförs i enlighet med gällande internationella metoder är det nödvändigt att ändra vissa bestämmelser.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av rådets direktiv 76/114/EEG av den 18 december 1975 om tillnärmning av medlemsstaternas lagstiftning om föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt på motorfordon och släpvagnar till dessa fordon(2), och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
om föreskrivna skyltar och märkningar samt deras placering och fastsättning på fordonstypen eller fordonet överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
3. Från den 1 oktober 1981 får medlemsstaterna förbjuda att fordon tas i bruk om deras föreskrivna skyltar och märkningar samt placering och fastsättning inte överensstämmer med bestämmelserna i direktiv 76/114/EEG, i dess lydelse enligt detta direktiv.
Artikel 4
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag,
För detta ändamål bör en förteckning utarbetas över de åtgärder som motsvarar begreppet intervention för stabilisering av marknaderna.
De olika utgifts- och intäktsslagen för varje sektor på grundval av dessa regler bör bli föremål för närmare bestämmelser. Under tiden bör finansieringsförordningarna för varje sektor fortsätta att gälla.
Artikel 1
När, inom ramen för den gemensamma organisationen av marknaden, ett belopp fastställs per enhet för en interventionsåtgärd skall utgifterna i samband med detta helt täckas av gemenskapsmedel.
Artikel 4
I fråga om medel som har sitt ursprung i medlemsstaterna och som används till interventionsköp av produkter, skall de räntekostnader som skall finansieras av garantisektionen vid EUGFJ beräknas enligt en metod och en räntesats som är enhetlig inom hela gemenskapen och som skall fastställas enligt det förfarande som avses i enlighet med artikel 13 i förordning (EEG) nr 729/70. Räntesatsen skall vara representativ för de faktiska räntesatser som tillämpas.
Artikel 7
I de årsräkenskaper som anges i artikel 4.1 skall de kvantiteter lagrade produkter som skall överföras till påföljande räkenskapsår som regel värderas till sina inköpspriser. För detta ändamål skall det pris som skall tillämpas för kvantiteter som överförs till påföljande räkenskapsår fastställas för de olika produkterna enligt förfarandet i artikel 13 i förordning (EEG) nr 729/70, på grundval av de inköpspriser som betalats av interventionsorganen under en referensperiod och med beaktande av den värdeminskning som anges i artikel 7.
Vid behov skall tillämpningsföreskrifter för denna förordning antas i enlighet med förfarandet i artikel 13 i förordning (EEG) nr 729/70.
Artikel 11
med beaktande av rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(1), senast ändrad genom direktiv 78/547/EEG(2), och särskilt artiklarna 11, 12 och 13 i detta,
Bestämmelserna i detta direktiv är i överenstämmelse med yttrandet från Kommittén för anpassning till teknisk utveckling av direktiv om avskaffande av tekniska handelshinder inom motorfordonssektorn.
1. Bilagorna 1, 2, 3, 4, 5, 6 och 9 till direktiv 71/320/EEG ändras härmed enligt bilagan till detta direktiv.
1. Från den 1 januari 1980 får ingen medlemsstat, av skäl som hänför sig till bromsutrustningen,
om bromsutrustningen på fordonstypen eller fordonen överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
- vägra att bevilja ett nationellt typgodkännande för en fordonstyp vars bromsutrustning inte överensstämmer med bestämmelserna i direktiv 71/320/EEG, i dess senaste lydelse enligt detta direktiv.
5. Före den 1 januari 1980 skall medlemsstaterna sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv och genast underrätta kommissionen om detta.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I artikel 6 i kommissionens förordning (EEG) nr 2960/77(3) föreskrivs att eventuella köpare får ta ett prov på de oljor som säljs av interventionsorganen.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för oljor och fetter.
Förordning (EEG) nr 2960/77 skall ändras på följande sätt: 1. Artikel 5.3 skall ersättas med följande:
"Detta prov skall placeras i två etiketterade flaskor, som skall plomberas i närvaro av både den som är ansvarig för lagret och den eventuelle köparen eller dennes vederbörligen bemyndigade företrädare. En flaska skall lämnas till den eventuelle köparen och den andra till den som är ansvarig för lagret."
"Innan plomberingen utförs får den vars anbud antagits begära ett prov på denna olja. Detta prov skall placeras i två etiketterade flaskor, som skall plomberas i närvaro av både den som är ansvarig för lagret och den vars anbud antagits eller dennes vederbörligen bemyndigade företrädare. En flaska skall lämnas till anbudsgivaren och den andra till den som är ansvarig för lagret så att det vid behov kan kontrolleras att den vara som ett prov togs på enligt artikel 6 och den vara som tilldelats stämmer överens."
2. Den kvantitet olja som levererats till köparen får avvika från den kvantitet för vilken anbudet lämnades, beroende på den faktiska kvantiteten i behållaren vid leveranstillfället."
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 99 och 100 i detta,
I överensstämmelse med domstolens dom av den 10 oktober 1978 i mål 148-77 tillämpas fördraget och härledd lagstifting på de franska utomeuropeiska departementen, såvida inte gemenskapens institutioner beslutar om särskilda åtgärder som är anpassade till de ekonomiska och sociala villkoren i dessa departement.
Följande strecksats skall läggas till i artikel 3.2 i direktiv 77/388/EEG"- Frankrike:
Detta direktiv skall tillämpas från och med den 1 januari 1979.
KOMMISSIONENS FÖRORDNING (EEG) nr 1698/80 av den 30 juni 1980 om tillägg till förordning (EEG) nr 797/80 om justering av förutfastställda exportavgifter och exportbidrag för socker
med beaktande av rådets förordning (EEG) nr 3330/74 av den 19 december 1974 om den gemensamma organisationen av marknaden för socker(), senast ändrad genom förordning (EEG) nr 1396/78(), särskilt artiklarna 17.5, 19.2 och 19.4 i denna, och
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för socker.
Artikel 1 i förordning (EEG) nr 797/80 skall ändras på följande sätt: 1. I punkt 1 skall "på begäran av berörd part" utgå.
Artikel 2
RÅDETS DIREKTIV av den 20 juli 1981 om ändring av rådets direktiv 77/541/EEG om tillnärmning av medlemsstaternas lagstiftning om bilbälten och fasthållningsanordningar i motorfordon (81/576/EEG)
med beaktande av kommissionens förslag(1),
med beaktande av följande: Rådets direktiv 77/541/EEG av den 28 juni 1977 om tillnärmning av medlemsstaternas lagstiftning om bilbälten och fasthållningsanordningar i motorfordon(4) uppställer bl.a. i bilaga 1 krav på montering av bilbälten och fasthållningsanordningar i fordon i kategori M1 enligt definition i bilaga 1 i rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(5), senast ändrat genom direktiv 80/1267/EEG(6).
Ändring av detta direktiv innebär anpassning till den tekniska utvecklingen av vissa krav i bilagorna till direktiv 77/541/EEG. Ikraftträdandet av bestämmelserna i det nuvarande direktivet bör fås att sammanfalla med ikraftträdandet av bestämmelserna som efter antagande av det nuvarande direktivet kommer att antas för anpassning av kraven i bilagorna till direktiv 77/541/EEG till den tekniska utvecklingen.
I detta direktiv avses med "fordon" varje motorfordon i kategorierna M och N enligt definition i bilaga 1 till direktiv 70/156/EEG som är avsett att användas på väg, som har minst fyra hjul och som är konstruerat för en högsta hastighet som överstiger 25 km/tim."
Varje fordon som omfattas av artikel 9 och tillhör kategorierna M1 eller N1 eller kategori M2 (utom fordon med en tillåten största vikt som överstiger 3 500 kg och fordon med utrymmen särskilt utformade för stående passagerare) skall vara utrustade med bilbälten eller fasthållningsanordningar som uppfyller kraven i detta direktiv och har följande bältesarrangemang (som varken medger att låsningsfria upprullningsdon [1.8.1] eller upprullningsdon med manuell upplåsning [1.8.2] kan användas).
"3.1.1 För främre yttre sittplatser, trepunktsbilbälte med nödlåsande upprullningsdon med flerfunktion (1.8.4). Följande skall dock gälla: 3.1.1.1 För passagerarsätet är automatiskt låsande upprullningsdon (1.8.3) tillåtna.
c) Avsnitt 3.1.3 skall ersättas med följande:
"3.1.5 Oavsett föregående bestämmelser får ett nödlåsande upprullningsdon av typ 4 N (1.8.5) tillåtas i stället för ett upprullningsdon av typ 4 (1.8.4) i fordon i kategorierna N1 och M2, där det på ett tillfredsställande sätt har visats för provningsorganet som ansvarar för provningarna att montering av ett upprullningsdon av typ 4 skulle besvära föraren."
Artikel 3
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(1), och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av följande: Genom rådets förordning (EEG) nr 3179/78() antog gemenskapen konventionen om framtida multilateralt samarbete om fisket i Nordvästatlanten.
Det är därför nödvändigt att förordning 3179/78 slutgiltigt ändras.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
För att få redovisningsresultat som är tillräckligt enhetliga på gemenskapsnivå bör de rapporterande företagen fördelas efter områden och de olika företagskategorierna genom att undersökningsområdet delas in enligt gemenskapens typologi för jordbruksföretag, fastställd genom beslut 78/463/EEG ().
Erfarenheten visar att det inte längre är önskvärt att införa tilläggsvillkor i det avtal som skall slutas mellan medlemsstaten och bokföringsbyråerna.
Följande fotnot skall läggas till längst ner på sidan:
"Artikel 4
a) ha en storlek som i ekonomiskt avseende är lika med eller större än ett tröskelvärde som fastställs enligt punkt 1,
3. Det högsta antalet rapporterande företag skall vara 45 000.
"Artikel 5
a) planen för val av rapporterande företag, särskilt hur de rapporterande företagen skall fördelas per företagskategori och tillämpningsföreskrifterna för val av företag,
Den nationella kommitténs beslut skall vara enhälliga. Om enighet inte kan uppnås skall beslut fattas av en myndighet som medlemsstaten utser.
5. Tillämpningsföreskrifterna till denna artikel skall antas enligt förfarandet i artikel 19."
1. Varje medlemsstat skall tillsätta ett samordningsorgan, vars uppgifter skall vara
P planen för val av rapporterande företag, vilken skall utarbetas med de senaste statistikuppgifterna som underlag, sammanställd enligt gemenskapens typologi för jordbruksföretag,
P förteckningen över rapporterande företag,
f) att till den nationella kommittén, de regionala kommittéerna och bokföringsbyråerna överlämna alla förfrågningar om information som avses i artikel 16 och att överlämna svaren på dessa till kommissionen.
6) Artikel 16.1 skall ersättas med följande:
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 75 i detta,
med beaktande av följande: Rådet har samrått med Ekonomiska och sociala kommittén om kommissionens förslag med stöd av artikel 198 första stycket i fördraget. Kommittén har inte kunnat inkomma med sitt yttrande inom den av rådet utsatta tiden. Artikel 198 andra stycket i fördraget tillåter rådet att vidta fortsatta åtgärder även utan sådant yttrande. Rådet anser att denna möjlighet måste utnyttjas med tanke på vikten av att erforderliga ändringar snabbt antas.
Artikel 1
P ¼ñãáíéóðüò Óéäçñïäñüìùí ¸ëëÜäïò A.E. (ÏÓÅ)."
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: Mot bakgrund av den vetenskapliga och tekniska kunskapsutvecklingen bör bilaga 1 och 2 till direktiv 66/401/EEG och 69/208/EEG ändras av nedan angivna skäl.
De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga kommittén för utsäde och uppförökningsmaterial för jordbruk, trädgårdsnäring och skogsbruk.
Bilaga 1 till direktiv 66/401/EEG ändras på följande sätt:
Artikel 2
Lägsta sortrenhet skall främst undersökas vid fältbesiktningar som utförs enligt de villkor som fastställts i bilaga 1."
Punkt 3 skall ersättas med följande:
Artikel 4
"Utsädet skall ha tillräcklig sortäkthet och sortrenhet. I synnerhet skall utsäde av nedan angivna arter motsvara följande standarder eller andra villkor:
Artikel 5
Artikel 7
- bestämmelserna i artikel 2 i fråga om Poa spp., med verkan från och med den 1 januari 1983,
Artikel 8
med beaktande av kommissionens förslag, och
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 84.2 i detta, och
Artikel 3
c) den typ av sjöfartstjänst som berörs (t.ex. linjefart),
f) motåtgärdens rimlighet i förhållande till skadan.
Artikel 5
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande (2),
Direktivet har kompletterats med direktiv 83/349/EEG (5) om sammanställd redovisning.
Medlemsstaterna måste ges rätt att godkänna personer som, utan att uppfylla alla de krav som ställs på teoretisk utbildning, ändå under lång tid genom yrkesmässig verksamhet har fått tillräcklig erfarenhet inom områdena ekonomi, juridik och redovisning samt har godkänts vid yrkesexamen.
Fysiska personer som utför lagstadgad revision av räkenskaper på ett sådant revisionsbolags vägnar måste uppfylla villkoren i detta direktiv.
Detta direktiv berör varken den etableringsfrihet eller den rätt att fritt tillhandahålla tjänster som tillkommer personer med uppgift att utföra lagstadgad revision av räkenskaper.
AVSNITT I
b) utföra lagstadgad granskning av sammanställda bokslut och verifiera att innehållet i de sammanställda förvaltningsberättelserna är förenligt med de sammanställda boksluten, förutsatt att sådan granskning och verifiering föreskrivs i gemenskapsrätten.
Artikel 2
ii) En majoritet av röstetalet skall tillkomma fysiska personer eller revisionsbolag som uppfyller minst de i artikel 3-19 uppställda villkoren, med undantag för artikel 11.1 b; medlemsstaterna får föreskriva att sådana fysiska personer och revisionsbolag även skall vara godkända. De medlemsstater som då detta direktiv antas inte kräver nu angiven majoritet behöver dock inte föreskriva sådan, förutsatt att alla aktier eller andra andelar i revisionsbolaget är ställda till viss man och kan överlåtas endast med samtycke av revisionsbolaget och/eller, om medlemsstaten föreskriver det, med godkännande av behörig myndighet.
2. Då bestämmelserna i detta direktiv tillämpas, får de uppgifter som ankommer på medlemsstaternas myndigheter utövas av yrkesföreningar, om dessa enligt nationell lagstiftning har befogenhet att lämna sådant godkännande som avses i direktivet.
Artikel 4
Det i examen ingående teoretiska kunskapsprovet måste särskilt omfatta följande ämnesområden: a) - räkenskapsrevision,
- sammanställd redovisning,
- föreskrifter om upprättande av års- och sammanställt bokslut samt föreskrifter om metoder för värdering av balansposter och beräkning av resultatposter,
- lagstiftning om konkurs och liknande förfaranden,
- lagstiftning om social trygghet och arbetsrätt,
- matematik och statistik,
1. Med avvikelse från bestämmelserna i artikel 5 och 6 får en medlemsstat föreskriva att personer med universitetsexamen eller annan likvärdig examen eller med likvärdiga betyg i ett eller flera av de i artikel 6 angivna ämnena, får befrias från att avlägga teoretiska kunskapsprov i de ämnen som täcks av denna examen eller dessa betyg.
1. För att garantera förmågan att praktiskt tillämpa de teoretiska kunskaperna, vilken förmåga även prövas i examen, skall under minst tre år en praktisk utbildning äga rum som bl.a. skall omfatta revision av årsbokslut och sammanställda bokslut eller liknande redovisningshandlingar. Denna praktiska utbildning måste till minst två tredjedelar fullgöras hos någon som enligt medlemsstatens lagstiftning är godkänd i överensstämmelse med detta direktiv; medlemsstaten får dock tillåta att den praktiska utbildningen fullgörs hos någon som enligt en annan medlemsstats lagstiftning är godkänd i överensstämmelse med detta direktiv.
Medlemsstaterna får tillåta personer att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna även om de inte uppfyller villkoren enligt artikel 4, under förutsättning att de kan visa a) att de under 15 år har utövat yrkesmässig verksamhet som har gett dem möjligheter att förvärva tillräcklig erfarenhet på ekonomi-, juridik- och redovisningsområdena samt har godkänts vid en sådan yrkesexamen som avses i artikel 4, eller
1. Medlemsstaterna får från de i artikel 9 angivna åren för yrkesmässig verksamhet räkna av tid för teoretisk utbildning inom de ämnesområden som anges i artikel 6, förutsatt att denna utbildning har avslutats med en statligt erkänd examen. Utbildningen får inte understiga ett år och får inte heller med mer än fyra år räknas av från tiden för yrkesmässig verksamhet.
1. Myndigheterna i en medlemsstat får godkänna personer som helt eller delvis har förvärvat sina kvalifikationer i någon annan stat, om dessa personer uppfyller följande två villkor: a) en behörig myndighet skall finna att deras kompetens är likvärdig med den som krävs enligt medlemsstatens lagstiftning i överensstämmelse med detta direktiv, och
Artikel 12
Artikel 13
1. En medlemsstat får anse sådana revisionsbolag som godkända enligt detta direktiv, vilka har godkänts genom förvaltningsbeslut av en behörig myndighet i den medlemsstaten innan de i artikel 30.2 avsedda bestämmelserna skall börja tillämpas.
Artikel 15
Artikel 18
Artikel 19
I avvaktan på en senare samordning av den lagstadgade revisionen av räkenskapshandlingar får en medlemsstat - som inte utnyttjar den i artikel 51.2 i direktiv 78/660/EEG angivna möjligheten och i vilken stat, då detta direktiv antas, flera kategorier fysiska personer enligt nationell lagstiftning är behöriga att utföra lagstadgad revision av de i artikel 1.1 a angivna handlingarna - särskilt godkänna fysiska personer som handlar i eget namn att utföra lagstadgad revision av de i artikel 1.1 a angivna handlingarna i bolag som inte överskrider gränserna för två av de tre kriterierna i artikel 27 i direktiv 78/660/EEG, om dessa personer: a) uppfyller de i artikel 3-19 i detta direktiv ställda villkoren, dock att nivån för yrkesexamen får vara lägre än vad som krävs enligt artikel 4, och
Artikel 21
En medlemsstat som tillämpar artikel 20 får i fråga om där avsedda personer tillåta att den i artikel 8 angivna praktiska utbildningen fullgörs hos någon som enligt den statens lagstiftning har godkänts att utföra sådan lagstadgad revision som avses i artikel 20.
Medlemsstaterna skall föreskriva att de personer som har godkänts att utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna skall utföra revisionen med yrkesmässig omsorg.
Artikel 25
Medlemsstaterna skall säkerställa att godkända personer blir föremål för lämpliga påföljder om de inte utför revisionen enligt artikel 23, 24 och 25.
AVSNITT IV Offentliggörande
2. Därutöver skall följande uppgifter om varje godkänt revisionsbolag vara offentligt tillgängliga: a) Namn och adress för de fysiska personer som anges i artikel 2.1 b i.
3. I de fall en fysisk person får utföra lagstadgad revision av de i artikel 1.1 angivna handlingarna under de förutsättningar som anges i artikel 20, 21 och 22 skall punkt 1 i denna artikel tillämpas. Därvid skall emellertid anges i vilka kategorier av bolag och företagsgrupper som en sådan revision får utföras.
Den kontaktkommitté som har tillsatts enligt artikel 52 i direktiv 78/660/EEG skall även: a) med förbehåll för artikel 169 och 170 i Romfördraget underlätta en enhetlig tillämpning av detta direktiv genom regelbundet samråd, särskilt om praktiska problem i samband med tillämpningen,
1. Medlemsstaterna skall före den 1 januari 1988 sätta i kraft de lagar och andra författningar som behövs för att följa detta direktiv. De skall genast underrätta kommissionen om det.
4. Medlemsstaterna skall även till kommissionen överlämna förteckningar över examina som har anordnats eller erkänts i överensstämmelse med artikel 4.
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter(), senast ändrad genom förordning nr (EEG) nr 2260/84(), särskilt artikel 5.4 till denna,
I avvaktan på upprättandet av ett register för olivodling, bör stödet till de berörda odlarna beräknas på grundval av den genomsnittliga avkastningen av olivträd.
De sammanslutningar av organisationer för olivoljeproducenter som avses i artikel 20c.2 i den förordningen bör bestå av ett minimiantal av grupper eller representera en minsta procentuella andel av den inhemska produktionen. Dessa minsta antal eller andelar bör fastställas på en nivå som gör det möjligt att utföra det speciella samordnings- och kontrollarbete som dessa sammanslutningar är skyldiga att utföra på ett effektivt sätt.
Enligt artikel 20d.1 i den förordningen får en del av stödbeloppet behållas för att täcka de utgifter som producentorganisationer och sammanslutningar av dessa ådrar sig för att utföra kontrollarbetet. Åtgärder bör vidtas för att säkerställa att dessa belopp endast används för att betala för de arbetsuppgifter som avses i artiklarna 20c.1 och 20c.2 i den förordningen.
Ifrågavarande stöd är till stor fördel för oljeproducenterna och utgör en finansiell börda för gemenskapen. För att säkerställa att stödet endast beviljas för olja som är berättigad till det, bör bestämmelser fastställas om inrättandet av ett lämpligt system för administrativa kontroller.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
3. Stödet skall beviljas efter ansökan från de berörda parterna till den medlemsstat i vilken oljan har framställts.
5. För regleringsåren 1984/85 och 1985/86 skall de producerande medlemsstaterna bestämma vilka olivodlare, med en genomsnittlig produktion av minst 100 kg olja per regleringsår, som är berättigade att erhålla stöd, beviljat efter den kvantitet av olja som verkligen har framställts, genom användning av avkastningen av oliver och olivolja fastställd enligt artikel 18, i förhållande till antalet olivträd i produktionen.
1. Varje olivodlare skall vid början av regleringsåret och före en fastställd dag till de behöriga myndigheterna i medlemsstaten i fråga inge en skördedeklaration, som vid första tillfället det inges skall innehålla:
2. Under de följande regleringsåren skall varje olivodlare, före en dag som skall fastställas, inge en kompletterande deklaration, i vilken odlaren uppger alla förändringar som har skett eller att den tidigare lämnade skördedeklarationen fortfarande är tillämplig.
Producentorganisationerna skall till den behöriga medlemsstaten anmäla namnen på de olivodlare som avses i andra stycket.
- upplysningar om den avsedda användningen av oliverna.
1. Med beaktande av de andra kraven i artikel 20c.1 i förordning nr 136/66/EEG får en producentorganisation inte godkännas enligt den förordningen om den inte
c) företräder minst 25 % av olivodlarna eller produktionen av olivolja i den ekonomiska region där den har upprättats.
3. I detta direktiv avses med ekonomisk region ett område som, enligt kännetecken som skall fastställas av den berörda medlemsstaten, har likartade produktionsvillkor med avseende på olivodling.
1. Producentorganisationer som önskar bli erkända från början av ett regleringsår skall ansöka hos den behöriga myndigheten i medlemsstaten i fråga senast den 30 juni under det föregående regleringsåret.
3. Godkända producentorganisationer skall senast den 30 juni varje år anmäla alla ändringar som skett i deras organisationer efter deras godkännande eller sedan den sista årliga deklarationen inlämnades och anmäla alla mottagna återkallelser av eller ansökningar om medlemskap till den behöriga myndigheten.
Artikel 6
- utföra kontroller på plats av de upplysningar som lämnats, i en viss del av dessa deklarationer, vilken skall fastställas,
2. Om en producentorganisation tillhör en sammanslutning av dessa organisationer, skall skördedeklarationerna och ansökningarna om stöd från de olivodlare som är medlemmar överlämnas av sammanslutningen.
- även har arrenderat olivodlingar för mindre än tre år,
Artikel 8
- att de uppgifter som lämnats av varje odlare i fråga om de kvantiteter av oliver som pressats och de kvantiteter av olja som erhållits stämmer överens med de kvantiteter av oliver och olja som uppgivits i bokföringen hos de godkända fabrikerna.
- Om de upplysningar som anges i punkt 1 andra strecksatsen inte förefaller att stämma överens.
1. Med beaktande av kraven i artikel 20c.2 i förordning nr 136/66/EEG får en sammanslutning inte godkännas om den inte består av minst 10 producentorganisationer, godkända enligt artikel 5, eller ett antal organisationer som svarar för minst 5 % av den olivolja som framställs i den berörda medlemsstaten.
De sammanslutningar som avses i artikel 20c.2 i förordning nr 136/66/EEG
- skall ta emot förskott av produktionsstödet, såsom anges i artikel 12, och saldot på stödbeloppen från den berörda medlemsstaten och skall snarast dela upp dem mellan de producenter som är medlemmar i de organisationer som tillhör dem.
a) Ett belopp som skall fastställas skall utbetalas till varje sammanslutning på grundval av antalet medlemmar i de producentorganisationer som tillhör den.
- kontroller som utförts enligt förfarandet för erhållande av stöd.
4. För att underlätta verksamheten i sammanslutningar och producentorganisationer är medlemsstaterna behöriga att i början av varje regleringsår betala dem ett förskott, som skall beräknas på grundval av en enhetstaxa för antalet medlemmar.
1. De producerande medlemsstaterna skall ha rätt att till sammanslutningar av producentorganisationer utbetala ett förskott på de yrkade stödbeloppen.
- 50 % av det belopp som erhålls vid beräkning av ett genomsnitt av de stödbelopp som betalats under de två föregående regleringsåren.
a) till medlemsstaten i fråga, enligt bestämmelser som skall fastställas, har överlämnat fullständiga upplysningar om fabrikens tekniska utrustning och nuvarande pressningskapacitet samt alla ändringar av dessa uppgifter,
- inte blivit föremål för åtgärder rörande oriktigheter som upptäckts vid kontroller gjorda för regleringsåret 1983/1984 enligt artikel 7 och 9 i förordning (EEG) nr 2959/82(), och
2. Medlemsstaterna skall innan de beviljar ett godkännande kontrollera om villkoren för ett godkännande är uppfyllda och skall särskilt på platsen kontrollera den tekniska utrustningen och den faktiska pressningskapaciteten i fabrikerna.
Om det visar sig att ett av de villkor som anges i punkt 1 inte är uppfyllt, skall det tillfälliga godkännandet återkallas.
- samma fysiska eller juridiska person som förestår fabriken i fråga,
1. Varje producerande medlemsstat skall tillämpa ett kontrollsystem för att säkerställa att den produkt för vilken stöd beviljas är berättigad till detta stöd.
De utvalda fabrikerna skall vara representativa för pressningskapaciteten i ett produktionsområde.
- att de skördade oliverna skall användas för att framställa olja och, om möjligt, att de faktiskt har bearbetats till olja.
Dessa register skall användas som stöd i den kontrollverksamhet som skall förekomma enligt punkt 1 4.
Den kvantitet olivolja som avses i punkt 4 i bilagan till förordning nr 136/66/EEG för vilken stöd får medges skall bestämmas på grundval av den typ av olja som anges i punkt 1 i den bilagan.
Artikel 16
a) För varje olivodlare och för varje regleringsår som en ansökan om stöd har inlämnats
- uppgifter som erhållits vid de kontroller på plats som gjorts hos olivodlaren.
d) De förväntade årliga skördarna för varje enhetligt produktionsområde.
Följande organ skall ha tillgång till dem:
- Producentorganisationer och sammanslutningar av dessa, i fråga om de aspekter som medlemsstaterna anser vara nödvändiga för att effektivt kontrollera sina respektive medlemmar.
De skördar av oliver och olja som anges i artikel 5.2 första stycket andra strecksatsen i förordning nr 136/66/EEG skall fastställas för enhetliga produktionsområden, senast den 31 maj varje år på grundval av uppgifter som de producerande medlemsstaterna lämnar senast den 30 april varje år.
Följande uppgifter skall fastställas enligt samma förfarande:
Artikel 20
Före slutet av det tredje året under vilket denna förordning tillämpas skall kommissionen överlämna en rapport till rådet om den verksamhet som fastställs i denna förordning tillsammans med förslag om hur rådet skall ändra verksamheten.
Artikel 23
med beaktande av kommissionens förslag(),
med beaktande av följande: I syfte att göra hälsoskyddsåtgärderna enhetliga för konsumenterna fastställs bestämmelser i direktiv 64/433/EEG(), senast ändrat genom direktiv 83/90/EEG() om hygienundersökningar och kontroller av färskt kött som kan komma att införas i handeln inom gemenskapen.
Rådets direktiv 71/118/EEG(), senast ändrat genom direktiv 84/642/EEG() föreskriver att hälsoundersökningar och kontroller skall ske av färskt fjäderfäkött.
Med hänsyn till nationella förvaltnings- och finansieringsbestämmelser och -förfaranden bör en ytterligare frist på två år beviljas för att göra det möjligt för Grekland att införa det nödvändiga systemet för att ta ut avgifter i samband med undersökningar och kontroller.
1. Medlemsstaterna skall säkerställa att man från och med den 1 januari 1986
P förbjuder varje form av direkt eller indirekt återbetalning av avgifter.
Artikel 3
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 januari 1986. De skall genast underätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Ekonomiska och sociala kommitténs yttrande(), och
Enligt artikel 54.3 h i fördraget får medlemsstaterna inte bevilja någon form av stödåtgärder som skulle kunna snedvrida etableringsvillkoren.
Då ett direktiv om ömsesidigt erkännande av examensbevis inte nödvändigtvis innebär likvärdighet när det gäller den utbildning som dessa examensbevis avser, bör rätten att använda yrkestitlar på grundval av utbildningen endast vara tillåten på språket i ursprungslandet eller det senaste hemvistlandet.
Det är svårt att bedöma i vad mån föreskrifter i syfte att underlätta farmaceuters frihet att tillhandahålla tjänster f.n. kan vara till nytta; under nuvarande omständigheter bör några föreskrifter därför inte antas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Varje medlemsstat skall erkänna de utbildnings-, examens- och andra behörighetsbevis som tilldelas medborgare i medlemsstaterna av övriga medlemsstater i enlighet med artikel 2 i direktiv 85/432/EEG och som finns uppräknade i artikel 4 genom att ge dessa bevis, när det gäller rätten att påbörja och utöva sådan verksamhet som avses i artikel 1, samma innebörd inom sitt territorium som dem som medlemsstaten själv utfärdar.
Artikel 3
2. Tio år efter utgången av den tidsfrist som fastställts i artikel 19 skall kommissionen föreslå rådet lämpliga åtgärder för att utvidga verkningarna av ett ömsesidigt erkännande av utbildnings-, examens- och andra behörighetsbevis i syfte att underlätta det faktiska utövandet av etableringsrätten mellan Grekland och de övriga medlemsstaterna. Rådet skall vidta åtgärder med anledning av dessa förslag i enlighet med det förfarande som fastställts i fördraget.
a) I Belgien:
Bevis for bestået farmaceutisk kandidateksamen (intyg över genomgången farmaceutisk universitetsexamen).
2) Intyg från de behöriga myndigheterna i Tyskland som visar att de examensbevis som utfärdats efter den 8 maj 1945 av de behöriga myndigheterna i Tyska Demokratiska Republiken erkänns som likvärdiga med dem som avses i punkt 1 ovan.
e) I Frankrike:
Intyg som Registered Pharmaceutical Chemist.
h) I Luxemburg:
Het getuigschrift van med goed gevolg afgelegd apothekersexamen (bevis över genomgången farmaceutexamen).
Artikel 5
Artikel 6
- om de åtföljs av ett intyg som visar att innehavarna av dessa examensbevis i en medlemsstat faktiskt på föreskrivet sätt har utövat någon av de former av verksamhet som avses i artikel 1.2 i direktiv 85/432/EEG i minst tre år i följd under en femårsperiod före dagen för utfärdandet av intyget, förutsatt att det landet utfärdat bestämmelser som reglerar denna verksamhet.
1. Utan att det påverkar tillämpningen av artikel 14 skall värdlandet se till att medborgare i medlemsstaterna som uppfyller villkoren i artikel 2, 5 och 6 får rätt att använda den erkända akademiska titeln eller en eventuell förkortning av denna i ursprungslandet eller det senaste hemvistlandet på det landets språk. Värdlandet får kräva att denna titel åtföljs av namnet på och platsen för den institution eller examensnämnd som utfärdat den.
1. Ett värdland som kräver bevis om god vandel eller bevis om gott anseende av de egna medborgare som vill påbörja sådan verksamhet som avses i artikel 1 skall när det gäller medborgare från andra medlemsstater som tillräckligt bevis godta ett intyg utfärdat av en behörig myndighet i ursprungslandet eller det senaste hemvistlandet, som visar att det landets krav på god vandel eller gott anseende för att påbörja verksamheten i fråga är uppfyllda.
Artikel 9
Ursprungslandet eller det senaste hemvistlandet skall kontrollera riktigheten av sakförhållandena, om de sannolikt kommer att påverka rätten att i den medlemsstaten utöva verksamheten i fråga. Myndigheterna i det landet skall avgöra vilket slags utredningar som skall göras och i vilken omfattning och skall underrätta värdlandet om eventuella åtgärder som de vidtar med avseende på de upplysningar som överlämnats i enlighet med punkt 1.
Om det i ursprungslandet eller det senaste hemvistlandet inte ställs några krav av detta slag för att påbörja eller utöva verksamheten i fråga, skall värdlandet godta intyg som utfärdats av behörig myndighet i det andra landet och som motsvarar de intyg som utfärdas i värdlandet.
Artikel 12
Det ursprungsland eller senaste hemvistland som rådfrågats skall avge svar inom tre månader.
Om ett värdland kräver att de egna medborgare som vill påbörja eller utöva den verksamhet som avses i artikel 1 avlägger ed eller avger en högtidlig försäkran och om formen för en sådan ed eller försäkran inte kan användas av medborgare i andra medlemsstater, skall värdlandet se till att en lämplig och likvärdig form av ed eller försäkran erbjuds personen i fråga.
Artikel 15
2. Medlemsstaterna får upprätta de kontor som avses i punkt 1 vid de behöriga myndigheterna och organen, som de måste utse inom den tidsfrist som fastställts i artikel 19.1.
Om det finns skälig grund till tvivel får värdlandet kräva att de behöriga myndigheterna i en annan medlemsstat styrker äktheten av utbildnings-, examens- och andra behörighetsbevis som utfärdats i den andra medlemsstaten och som avses i kapitel II och III samt styrker att personen i fråga har uppfyllt utbildningsvillkoren i direktiv 85/432/EEG.
Artikel 18
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
I mån av behov skall kommissionen föreslå rådet lämpliga åtgärder.
RÅDETS DIREKTIV av den 20 december 1985 om samordning av lagar och andra författningar som avser företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag) (85/611/EEG)
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
Sådana gemensamma regler ger en tillräcklig garanti för att medlemsstaternas företag för kollektiva investeringar, med iakttagande av vad som skall gälla beträffande kapitalrörelser, skall kunna utbjuda sina andelar i andra medlemsstater utan att dessa skall ha möjlighet att för företagen eller deras andelar tillämpa några andra bestämmelser än sådana som faller utanför direktivets tillämpningsområde. Ett företag för kollektiva investeringar som utbjuder sina andelar i en annan medlemsstat än där företaget hör hemma, skall dock vidta alla åtgärder som krävs för att andelsägarna där skall kunna utöva sina finansiella rättigheter utan svårighet och få tillgång till nödvändig information.
Hänsyn bör tas till de särskilda omständigheter som råder beträffande de finansiella marknaderna i Grekland och Portugal genom att dessa länder medges en förlängd frist för att genomföra detta direktiv.
3. Sådana företag kan bildas med stöd av lag, antingen på kontraktsrättslig grund (som värdepappersfonder förvaltade av förvaltningsföretag) eller enligt trustlagstiftning (som "unit trusts") eller på bolagsrättslig grund (som investeringsbolag).
5. Medlemsstaterna skall förbjuda fondföretag för vilka detta direktiv gäller att ombilda sig till sådant företag för kollektiva investeringar som inte omfattas av direktivets bestämmelser.
Artikel 2
2. Senast fem år efter genomförandet av detta direktiv skall kommissionen överlämna en rapport till rådet över tillämpningen av bestämmelserna i punkt 1, särskilt dess fjärde strecksats. Om så erfordras skall kommissionen föreslå lämpliga åtgärder för att utöka bestämmelsernas tillämpningsområde.
AVSNITT II Auktorisation av fondföretag
Auktorisationen skall gälla i samtliga medlemsstater.
Med den verkställande ledningen avses de personer som, i enlighet med lag eller annan författning eller bolagsordning, företräder förvaltningsbolaget, investeringsbolaget eller förvaringsinstitutet eller som faktiskt bestämmer verksamhetsinriktningen för sådana företag.
Artikel 5
Ett förvaltningsbolag får inte ägna sig åt annan verksamhet än förvaltning av värdepappersfonder och investeringsbolag.
2. Ett förvaringsinstituts ansvarighet enligt artikel 9 skall gälla oberoende av om institutet anförtrott förvaringen av samtliga eller vissa tillgångar till någon annan.
Artikel 8
3. Medlemsstaterna skall bestämma vilka av de kategorier av institut som avses i punkt 2 som skall kunna utses till förvaringsinstitut.
Artikel 10
Artikel 11
Artikel 12
Ett investeringsbolag får inte bedriva andra verksamheter än de som anges i artikel 1.2.
2. Ett förvaringsinstituts ansvarighet enligt artikel 16 skall gälla oberoende av om institutet anförtrott förvaringen av samtliga eller vissa tillgångar till någon annan.
c) tillse att ett bolags intäkter används i enlighet med lag eller annan författning och med bolagsordningen.
5. En medlemsstat får bestämma att investeringsbolag som hör hemma i den staten och som utbjuder minst 80% av sina andelar på en eller flera fondbörser, vilka finns angivna i deras bolagsordningar, inte skall vara skyldiga att ha förvaringsinstitut som avses i detta direktiv, förutsatt att deras andelar noteras officiellt på fondbörserna i de medlemsstater där andelarna utbjuds, och att varje transaktion som ett sådant investeringsbolag kan komma att göra utanför fondbörserna sker uteslutande till börskurs. I ett investeringsbolags bolagsordning skall anges en fondbörs i varje land där andelar utbjuds och vars kursnotering skall vara bestämmande för de priser som skall gälla vid transaktioner som bolaget genomför utanför fondbörser i det landet.
c) fastställa andelarnas nettovärde, lämna uppgift om nettovärdet till de behöriga myndigheterna minst två gånger per vecka och offentliggöra uppgifter om nettovärdet två gånger per månad.
Kommissionen skall senast inom fem år från det att detta direktiv genomförts underrätta kontaktkommittén om tillämpningen av bestämmelserna i punkterna 4 och 5. När kontaktkommitténs yttrande erhållits skall kommissionen, om det behövs, föreslå lämpliga åtgärder.
2. Ett förvaringsinstitut skall stå under offentlig tillsyn. Det skall också kunna ställa erforderliga ekonomiska garantier samt besitta tillfredsställande sakkunskap och kompetens för att kunna effektivt bedriva verksamhet som förvaringsinstitut och uppfylla därmed förenade åtaganden.
Ett förvaringsinstitut skall i enlighet med den nationella lagstiftningen i den stat där investeringsbolaget har sitt stadgeenliga säte vara ansvarigt mot investeringsbolaget och andelsägarna för förluster som drabbar dem som följd av att institutet allvarligt försummat sina förpliktelser eller fullgjort dem på ett oriktigt sätt.
2. Ett förvaringsinstitut skall vid utförande av sina uppgifter handla uteslutande i andelsägarnas intresse.
AVSNITT V Placeringsbestämmelser för fondföretag
c) överlåtbara värdepapper som är officiellt noterade på en fondbörs i en icke-medlemsstat eller som är föremål för handel på någon annan reglerad marknadsplats i en icke-medlemsstat och vilken marknadsplats fungerar fortlöpande och är erkänd och öppen för allmänheten, förutsatt att valet av fondbörs eller annan marknadsplats godkänts av de behöriga myndigheterna eller är reglerat i lag eller annan författning eller i fondbestämmelserna eller i investeringsbolagets bolagsordning, och/eller
c) ett investeringsbolag får förvärva lös och fast egendom som det behöver för sin verksamhet,
4. Värdepappersfonder och investeringsbolag får ha kompletterande likvida tillgångar.
1. Medlemsstaterna får ge fondföretag tillstånd att använda sig av sådan teknik och sådana instrument som hänför sig till överlåtbara värdepapper under de villkor och inom de ramar staterna föreskriver, förutsatt att sådan teknik och sådana instrument används i syfte att åstadkomma en effektiv förvaltning av värdepappersportföljen.
1. Ett fondföretag får placera högst 5% av fondtillgångarna i överlåtbara värdepapper med samme utgivare.
Artikel 23
Ett sådant fondföretag skall inneha värdepapper från minst sex olika emissioner, varvid dock skall gälla att värdepapper från en och samma emission inte får motsvara mer än 30% av de samlade fondtillgångarna.
Artikel 24
3. Placeringar i andelar i en värdepappersfond som förvaltas av samma förvaltningsbolag eller av ett annat företag med vilket förvaltningsbolaget är anknutet via gemensam företagsledning eller ägarkontroll eller genom ett betydande direkt eller indirekt ägande får tillåtas endast om det rör sig om en fond som, i enlighet med sina fondbestämmelser, har specialiserat sig på placeringar inom ett visst geografiskt område eller en viss ekonomisk sektor och förutsatt att sådana placeringar medges av de behöriga myndigheterna. Tillstånd skall ges endast om fonden har meddelat sin avsikt att utnyttja denna möjlighet och möjligheten uttryckligen angivits i dess fondbestämmelser.
1. Ett investeringsbolag eller ett förvaltningsbolag får, såvitt gäller handhavandet av alla de värdepappersfonder som står under bolagets förvaltning och som omfattas av bestämmelserna i detta direktiv, inte förvärva aktier med sådan rösträtt som skulle göra det möjligt för bolaget att utöva ett väsentligt inflytande över ledningen hos en emittent.
- 10% av andelarna i ett sådant företag för kollektiva investeringar som avses i första och andra strecksatserna i artikel 1.2.
e) Ett investeringsbolags aktieinnehav i dotterbolag vars verksamhet består i förvaltning, rådgivning eller avsättning uteslutande för investeringsbolagets räkning.
Medlemsstaterna får, med beaktande av principen om riskspridning, tillåta nyligen auktoriserade fondföretag att under en tid av högst sex månader från auktorisationsdagen avvika från vad som föreskrivits i artiklarna 22 och 23.
Artikel 27
Artikel 28
3. Halvårsrapporten skall innehålla minst den information som anges i kapitel I-IV i lista B i bilagan till detta direktiv; om ett fondföretag har utbetalat eller föreslår utbetalning av interimsutdelning, skall i redovisningen anges resultatet efter skatt för halvårsperioden i fråga samt den interimsutdelning som utbetalats eller föreslås.
2. De handlingar som avses i punkt 1 behöver dock inte bifogas prospektet om andelsägarna informerats om att de på begäran kommer att tillställas dessa handlingar eller få upplysning om var i varje medlemsstat, där andelarna finns på marknaden, de kan ta del av handlingarna.
Artikel 31
Ett fondföretag skall till de behöriga myndigheterna ge in sina prospekt och eventuella ändringar och tillägg i dessa, liksom årsrapporter och halvårsrapporter.
2. Årsrapporterna och halvårsrapporterna skall finnas tillgängliga för allmänheten på i prospektet angivna platser.
Artikel 34
Vid all marknadsföring av ett fondföretags andelar skall anges att ett prospekt finns och uppges var allmänheten kan få tillgång till prospektet. AVSNITT VII
2. Trots bestämmelserna i punkt 1 får en medlemsstat ge fondföretag tillstånd att låna
b) upp till 10% av tillgångarna, i fråga om ett investeringsbolag, förutsatt att upplåningen har till syfte att möjliggöra förvärv av fast egendom som det behöver för verksamheten; i detta fall får summan av denna upplåning och den som avses i a inte överstiga 15% av låntagarens tillgångar.
b) Medlemsstaterna får tillåta de behöriga myndigheterna att kräva att återköp eller inlösen av andelar senareläggs med hänsyn till andelsägarnas eller allmänhetens intresse.
Reglerna för värdering av tillgångar och för beräkning av försäljnings- eller emissionspris samt återköps- eller inlösenpris på ett fondföretags andelar skall vara föreskrivna i lag eller annan författning, i fondbestämmelserna eller i investeringsbolagets bolagsordning.
Artikel 40
1. Med undantag för sådana fall som avses i artiklarna 19 och 21 gäller att varken
Artikel 42
I lag eller annan författning eller i ett investeringsbolags bolagsordning skall det anges vilka kostnader som skall bäras av bolaget.
1. Ett fondföretag som utbjuder sina andelar i en annan medlemsstat måste följa de lagar och andra författningar som gäller i den staten, och som inte faller inom tillämpningsområdet för detta direktiv.
Artikel 45
- sina fondbestämmelser eller sin bolagsordning,
Om ett fondföretag utbjuder sina andelar i en annan medlemsstat än den där företaget är beläget, skall det i den andra medlemsstaten, på minst ett av den andra medlemsstatens officiella språk, tillhandahålla de handlingar och den information som skall offentliggöras i den medlemsstat där det är hemmahörande, i den ordning som föreskrivs i den sistnämnda staten.
AVSNITT IX Bestämmelser om de myndigheter som svarar för auktorisation och tillsyn
2. De myndigheter som avses i punkt 1 skall vara offentliga myndigheter eller institutioner utsedda av offentliga myndigheter.
Artikel 50
3. Bestämmelserna i punkt 2 skall emellertid inte utesluta utbyte av information mellan de i artikel 49 angivna myndigheterna i olika medlemsstater i enlighet med bestämmelserna i detta direktiv. Beträffande sålunda utväxlad information skall anställda eller tidigare anställda hos myndigheter som erhåller information enligt ovan iaktta tystnadsplikt.
1. Myndigheter som avses i artikel 49 skall uppge skälen för såväl beslut att vägra auktorisation som de övriga beslut med negativ innebörd som fattas i samband med införande av föreskrifter för tillämpning av detta direktiv, samt underrätta sökandena om skälen.
1. Endast myndigheterna i den medlemsstat där ett fondföretag är beläget skall ha behörighet att vidta åtgärder mot företaget om det bryter mot lag eller annan författning eller fondbestämmelserna eller investeringsbolagets bolagsordning.
AVSNITT X Kontaktkommitté
a) att, så långt det inte strider mot artiklarna 169 och 170 i fördraget, underlätta ett samordnat genomförande av detta direktiv genom regelbundna samråd om praktiska problem som kan uppkomma vid dess tillämpning och beträffande vilka en diskussion bedöms ändamålsenlig,
2. Det skall inte ankomma på kommittén att pröva beslut som fattats i enskilda fall av de myndigheter som avses i artikel 49.
AVSNITT XI Övergångsbestämmelser, undantag och avslutande bestämmelser
Artikel 55
1. Trots bestämmelserna i artikel 6 får medlemsstaterna tillåta förvaltningsbolag att emittera innehavarbevis avseende andra företags registrerade värdepapper.
1. Medlemsstaterna skall senast den 1 oktober 1989 sätta i kraft de beslut som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
Ett år före detta datum skall kommissionen rapportera till rådet om hur genomförandet av direktivet fortgår och om eventuella svårigheter som kan uppkomma för Grekland eller Portugal att genomföra direktivet per det datum som anges i föregående stycke.
Medlemsstaterna skall se till att kommissionen erhåller uppgift om texterna till de viktigaste föreskrifterna som de antar inom det område som omfattas av detta direktiv.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 235 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
Fördraget innehåller inte tillräckliga bestämmelser för ett sådant rättsligt instrument.
Fysiska personer, bolag och andra rättsliga enheter bör enligt förordningens syfte i största möjliga utsträckning ha tillträde till denna företagsform. Förordningen hindrar dock inte att det på det nationella planet tillämpas rättsregler och/eller etiska regler som gäller utövningen av en verksamhet eller ett yrke.
För att en gruppering skall kunna fylla sitt ändamål skall den ha rättskapacitet. Ett organ som är rättsligt skilt från grupperingens medlemmar skall representera grupperingen mot tredje man.
Regler bör ges om särskilda grunder för upplösning av grupperingen, dock bör hänvisning ske till nationella rättsregler om likvidation och avslutning av denna.
I frågor som inte omfattas av denna förordning tillämpas medlemsstaternas rättsregler och gemenskapsrätten, t.ex. när det gäller
- immaterialrätt.
Denna förordning skall i sin helhet omedelbart träda i kraft. Tillämpningen av vissa bestämmelser skall dock senareläggas för att ge medlemsstaterna möjlighet att inrätta den administration inom sina respektive områden som behövs för registrering av grupperingarna och för att säkerställa att handlingar angående dessa blir offentliga. Från den dag förordningen tillämpas skall de grupperingar som bildas kunna verka utan territoriella inskränkningar.
1. Syftet med en grupperings verksamhet är att underlätta eller utveckla medlemmarnas ekonomiska verksamhet och att förbättra resultatet av denna verksamhet; en gruppering har inte till syfte att skapa vinst för egen del. En grupperings verksamhet skall knyta an till medlemmarnas ekonomiska verksamhet och får endast vara av understödjande karaktär i förhållande till den senare verksamheten.
b) under några omständigheter, varken direkt eller indirekt, inneha andelar eller aktier av något slag i ett företag som är medlem i grupperingen; innehav av andelar eller aktier i andra företag tillåts endast i den mån det är nödvändigt för att syftet med grupperingen skall uppnås och om det sker för medlemmarnas räkning,
e) vara medlem av någon annan europeisk ekonomisk intressegruppering.
a) Bolag som avses i artikel 58 andra stycket i fördraget och andra rättsliga enheter av offentligrättsligt eller privaträttsligt slag, som har bildats enligt en medlemsstats lagstiftning och som har sitt registrerade eller i lag bestämda säte samt sitt huvudkontor inom gemenskapen; om ett bolag eller en annan rättslig enhet enligt en medlemsstats lagstiftning inte behöver ha ett registrerat eller i lag bestämt säte, räcker det att bolaget eller den rättsliga enheten har sitt huvudkontor inom gemenskapen.
a) två bolag eller andra rättsliga enheter som avses i punkt 1 och som har sina huvudkontor i olika medlemsstater, eller
3. En medlemsstat kan bestämma att grupperingar som enligt artikel 6 är intagna i den statens register inte får ha mer än 20 medlemmar. Med hänsyn därtill får en sådan medlemsstat även bestämma att enligt dess lagstiftning varje medlem i en rättslig enhet, som har bildats enligt den lagstiftningen och som inte är ett registrerat bolag, skall behandlas som en särskild medlem när det gäller medlemskap i en gruppering.
Ett avtal om att bilda en gruppering skall innehålla minst följande uppgifter:
c) Föremålet för grupperingens verksamhet.
Artikel 6
Avtalet om att bilda en gruppering skall ges in till det register som anges i artikel 6.
c) Ett rättsligt avgörande som enligt artikel 15 fastställer eller tillkännager att grupperingen är ogiltig.
f) Ett beslut av medlemmarna varigenom grupperingen förklaras upplöst enligt artikel 31 eller ett rättsligt avgörande om upplösning enligt artikel 31 eller 32.
i) Förslag till byte av säte enligt artikel 14.1.
Följande skall offentliggöras enligt artikel 39 i den tidning som där anges i punkt 1:
c) I artikel 7 b-j avsedda handlingar och uppgifter.
1. De handlingar och uppgifter som skall offentliggöras på grund av denna förordning kan åberopas av en gruppering mot tredje man enligt vad som har bestämts i tillämplig nationell lagstiftning med stöd av artikel 3.5 och 3.7 i rådets direktiv 68/151/EEG av den 9 mars 1968 om samordning av de skyddsåtgärder som krävs i medlemsstaterna av de i artikel 58 andra stycket i Romfördraget avsedda bolagen i bolagsmännens och tredje mans intressen, i syfte att göra skyddsåtgärderna likvärdiga inom gemenskapen (4).
Ett huvudkontor eller avdelningskontor i någon annan medlemsstat än den där grupperingen har sitt säte skall registreras i den stat där kontoret är beläget. För detta ändamål skall grupperingen till den sistnämnda statens register ge in kopior av de handlingar som måste ges in till registret i den medlemsstat där grupperingen har sitt säte och, om det behövs, en översättning som uppfyller kraven vid det register där kontoret skall registreras.
Artikel 12
a) i den ort där grupperingen har sitt huvudkontor, eller
En gruppering får byta säte inom gemenskapen.
1. Om byte av säte medför att enligt artikel 2 någon annan lagstiftning blir tillämplig, skall förslag till bytet upprättas samt ges in och offentliggöras enligt föreskrifterna i artiklarna 7 och 8.
3. Sedan den nya registreringen har offentliggjorts kan det nya sätet åberopas mot tredje man enligt artikel 9.1; innan grupperingens avförande ur det tidigare registret har offentliggjorts får dock tredje man fortfarande åberopa det tidigare sätet, om grupperingen inte visar att tredje man kände till det nya.
1. Om en gruppering är ogiltig på grund av den lagstiftning som enligt artikel 2 är tillämplig, skall ogiltigheten fastställas eller tillkännages genom avgörande av en domstol. Den domstol som handlägger saken skall dock bestämma en frist inom vilken rättelse får ske, om grupperingens förhållanden kan bringas i överensstämmelse med gällande rätt.
Ett sådant avgörande enbart inverkar inte på giltigheten av de förpliktelser som grupperingen har ådragit sig eller som gäller till förmån för denna, om förpliktelserna har uppkommit innan avgörandet enligt föregående stycke kan göras gällande mot tredje man.
Avtalet om att bilda grupperingen kan innehålla bestämmelser om andra organ; i så fall skall avtalet ange dessas befogenheter.
1. Varje medlem har en röst. Avtalet om att bilda grupperingen kan dock tilldela vissa medlemmar flera röster förutsatt att ingen medlem får röstmajoritet.
b) ändra det antal röster som varje medlem har tilldelats,
e) ändra det belopp med vilket varje medlem eller vissa medlemmar skall bidra till grupperingens finansiering,
Artikel 18
1. En gruppering leds av en eller flera fysiska personer som utses i avtalet om att bilda grupperingen eller genom beslut av medlemmarna.
- enligt den interna lagstiftningen i den stat där grupperingen har sitt säte, eller
2. En medlemsstat kan för grupperingar som enligt artikel 6 är intagna i den statens register föreskriva att en juridisk person får vara företagsledare, under förutsättning att denne till sina representanter utser en eller flera fysiska personer för vilka bestämmelserna i artikel 7 d skall gälla.
3. Förutsättningarna för att utse och entlediga företagsledarna samt dessas befogenheter skall bestämmas i avtalet om att bilda grupperingen eller genom enhälligt beslut av medlemmarna.
När en företagsledare handlar på grupperingens vägnar förpliktar han denna mot tredje man även om hans handlingar faller utanför föremålet för grupperingens verksamhet, såvida inte grupperingen visar att tredje man kände till eller med hänsyn till omständigheterna inte kunde vara obekant med att handlingen föll utanför föremålet för grupperingens verksamhet; enbart offentliggörandet av den i artikel 5 c angivna uppgiften skall därvid inte anses tillräckligt som bevis.
Artikel 21
Artikel 22
Artikel 23
2. Innan likvidationen av en gruppering är avslutad får grupperingens borgenärer inte väcka talan mot en medlem för att få betalt enligt punkt 1, om de inte först har anmodat grupperingen att betala och betalning inte har erlagts inom skälig tid.
a) Grupperingens namn föregånget eller följt av orden "europeisk ekonomisk intressegruppering" eller förkortningen "EEIG", om inte orden eller förkortningen redan ingår i namnet.
d) I förekommande fall att företagsledarna endast får handla i förening.
Artikel 26
En medlem kan dock genom en bestämmelse i avtalet om att bilda grupperingen eller i inträdeshandlingen fritas från ansvar för förbindelser som har uppkommit före inträdet. En sådan bestämmelse kan göras gällande enligt artikel 9.1 mot tredje man, om den har offentliggjorts enligt artikel 8.
En sådan uteslutning får ske endast genom ett domstolsavgörande efter gemensam ansökan av en majoritet av de övriga medlemmarna, om inte något annat är bestämt i avtalet om att bilda grupperingen.
Dessutom kan en medlemsstat med hänsyn till sin lagstiftning om upplösning, likvidation, obestånd och betalningsinställelse bestämma att ett medlemskap skall upphöra vid tidpunkter som anges i den nämnda lagstiftningen.
Så snart någon upphör att vara medlem skall företagsledarna underrätta de övriga medlemmarna om det; företagsledarna skall dessutom vidta de åtgärder som krävs enligt artiklarna 7 och 8. De sistnämnda åtgärderna får även vidtas av var och en som saken angår.
Artikel 31
b) ändamålet med grupperingen har uppnåtts eller inte längre kan uppnås.
4. Efter upplösning av en gruppering genom beslut av medlemmarna skall företagsledarna vidta de åtgärder som krävs enligt artiklarna 7 och 8. Dessa åtgärder får även vidtas av var och en som saken angår.
2. På ansökan av en medlem får rätten förordna att en gruppering skall upplösas, om det föreligger en riktig grund för det.
Om någon upphör att vara medlem i en gruppering på annan grund än överlåtelse av rättigheter enligt artikel 22.1, skall värdet av den avgående medlemmens rättigheter och skyldigheter bestämmas med hänsyn till grupperingens förmögenhetsförhållanden vid tidpunkten för medlemskapets upphörande.
Med den begränsning som anges i artikel 37.1 svarar en avgången medlem enligt artikel 24 för de förbindelser som har uppkommit genom grupperingens verksamhet före avgången.
2. Likvidationen och avslutningen av denna skall ske enligt nationell rätt.
Artikel 36
1. En preskriptionstid på fem år räknat från offentliggörandet enligt artikel 8 av en medlems avgång gäller i stället för längre preskriptionstider i nationell lagstiftning i fråga om åtgärder mot den avgångne medlemmen med anledning av förbindelser som har uppkommit genom grupperingens verksamhet före avgången.
En behörig myndighet i en medlemsstat får förbjuda en gruppering att utöva verksamhet varigenom grupperingen åsidosätter allmänna intressen i den staten. Förbudet skall kunna prövas av domstol. Artikel 39
Medlemsstaterna får bestämma att avgifter skall erläggas för den verksamhet som avses i de två föregående styckena; avgifterna får dock inte överstiga de administrativa kostnaderna för verksamheten.
Artikel 40
1. Medlemsstaterna skall före den 1 juli 1989 vidta de åtgärder som krävs av dem enligt artikel 39. De skall underrätta kommissionen så snart åtgärderna har vidtagits.
1. När denna förordning har antagits skall en kontaktkommitté tillsättas under kommissionens överinseende. Kontaktkommitténs uppgift skall vara att
2. Kontaktkommittén skall bestå av representanter för medlemsstaterna och kommissionen. En representant för kommissionen skall vara ordförande. Kommissionen skall tillhandahålla ett sekretariat.
med beaktande av rådets förordning (EEG) nr 449/69 av den 11 mars 1969 om återbetalning av stöd som medlemsstaterna har beviljat frukt- och grönsaksproducenters organisationer(3), särskilt artikel 7.3 i denna, och
Det åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för Europeiska utvecklings- och garantifonden för jordbruket.
Bilagorna 1 och 2 i rådets förordning (EEG) nr 2264/69(6) skall ersättas med bilagorna 1 och 2 till denna förordning.
med beaktande av Anslutningsakten för Spanien och Portugal, särskilt artiklarna 171 och 358 i denna,
Detta program måste tillämpas på de kategorier av sardiner som kan förutses vara lättast att avsätta på marknaden efter beredning.
När det gäller de kvantiteter som berättigar till bidrag bör närmare bestämmelser införas för hur ansökningarna om utbetalning av bidraget skall lämnas in.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fiskeriprodukter.
- sålts till en beredare för fullständig och slutlig beredning i enlighet med de hygienföreskrifter och tekniska bestämmelser som gäller för livsmedelsprodukter i den medlemsstat där beredaren är etablerad.
b) framställning av konserver enligt nr 16.04 i gemensamma tulltaxan,
För varje parti av samma kommersiella kategori som säljs skall bidragets storlek bestämmas i enlighet med artikel 2.4 i förordning (EEG) nr 3117/85.
Av kontrollformuläret skall följande uppgifter framgå:
"VERARBEITUNG, FÜR DIE EINE AUSGLEICHS- ENTSCHÄDIGUNG GEWÄHRT WIRD
3. Producentorganisationen skall lämna in ansökan om utbetalning av bidraget till de behöriga myndigheterna i den berörda medlemsstaten före slutet av den första månaden efter det att försäljningsavtalet ingåtts.
2. De närmare bestämmelserna för hur kontrollen skall gå till skall utarbetas av medlemsstaten och omfatta minst följande krav:
- Närmare angivande av de uppgifter som skall ingå i den ansökan om bidrag som anges i artikel 5.
1. De berörda medlemsstaterna skall senast två månader efter ikraftträdandet av denna förordning anmäla till kommissionen vilka kontrollåtgärder som införts i enlighet med artikel 6.1.
Artikel 8
Denna förordning träder i kraft den 1 mars 1986, förutsatt att Anslutningsfördraget för Spanien och Portugal då trätt i kraft. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"- burro concentrato".
RÅDETS BESLUT av den 22 december 1986 om införande av en ordning för samråd och samarbete på turistområdet (86/664/EEG)
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
Samråd är ett bra medel för att underlätta samarbetet mellan medlemsstaterna och kommissionen i avsikt att uppnå fördragets mål.
Sådant samråd bör inte upprepa det arbete som utförts inom andra gemenskapsorgan.
En rådgivande turistkommitté, härefter kallad "kommittén", skall inrättas hos kommissionen. Den skall bestå av medlemmar utsedda av varje medlemsstat.
Artikel 3
Artikel 4
Artikel 5
med beaktande av Anslutningsakten för Spanien och Portugal, särskilt artikel 396 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
med beaktande av rådets förordning (EEG) nr 426/86 av den 24 februari 1986 om den gemensamma organisationen av marknaden för bearbetade produkter av frukt och grönsaker (), särskilt artikel 6.4 i denna, och
Med tanke på genomförandet av systemet med produktionsstöd måste denna förordning tillämpas tillsammans med kommissionens förordning (EEG) nr 1599/84 av den 5 juni 1984 om tillämpningsföreskrifter för produktionsstödet för bearbetade produkter av frukt och grönsaker (), senast ändrad genom förordning (EEG) nr 1155/86 (), särskilt vad gäller undersökning av de bearbetade produkterna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
P hela tomater eller tomater i bitar, skalade och konserverade enligt definitionen i artikel 1.2 h, ij, k och l i förordning (EEG) nr 1599/84.
P vatten,
P vanligt salt (natriumklorid),
2. Den totala tillsatsen av vanligt salt får inte överstiga 3 % av nettovikten och vid tillsättning av kalciumklorid får det totala kalciuminnehållet inte överstiga 0,045 % i hela tomater och 0,080 % i tomater i bitar. Vid bestämningen av tillsatsen vanligt salt skall det naturliga kloridinnehållet anses vara lika med 2 % av torrsubstansen.
1. Skalade tomater skall vara fria från främmande smaker och lukter och färgen skall vara karakteristisk för den sort som används och för korrekt bearbetade skalade tomater.
Artikel 6
P skal:
De fastställda gränsvärdena gäller per 10 kg nettovikt.
b) skal: både skal som sitter fast på tomatköttet och skal som påträffas löst i behållaren.
2. Den avrunna nettovikten för hela skalade tomater skall i genomsnitt vara lika med minst 56 % av behållarens volym uttryckt i gram.
I denna avdelning skall "tomatsaft" och "tomatkoncentrat" avse de produkter som definieras i artikel 1.2 n och o i förordning (EEG) nr 1599/84.
P vanligt salt (natriumklorid),
P tomatsaft med ett torrsubstansinnehåll på mindre än 7 %, får askorbinsyra (E 300) användas. Innehållet av askorbinsyra skall dock inte överstiga 0,03 % av den färdiga produktens vikt,
a) 15 viktprocent av torrsubstansinnehållet i tomatkoncentrat med ett torrrsubstansinnehåll som överstiger 20 %, och
Artikel 10
b) en god smak som är karakteristisk för en korrekt bearbetad produkt.
b) praktiskt taget fria från oorganiska orenheter.
b) halten av oorganiska orenheter inte överstiger 0,1 % av torrsubstansinnehållet, reducerat med eventuell tillsats av vanligt salt och vad avser tomatkoncentrat i pulverform, eventuell tillsats av kiseldioxid.
b) en sockerhalt uttryckt som invertsocker på minst 42 viktprocent av torrsubstansinnehållet minskat med eventuell tillsats av vanligt salt,
e) ett pH-värde på högst 4,5.
I denna avdelning skall "tomatflingor" avse den produkt som definieras i artikel 1.2 m i förordning (EEG) nr 1599/84.
a) ha en karakteristisk röd färg, och
2. Tomatflingors torrsubstanshalt skall vara minst 93 %.
Artikel 13
3. Märkningen som avses i denna artikel kan vara i form av en kod och skall godkännas av de behöriga myndigheterna i den medlemsstat där framställningen sker. Dessa myndigheter får fastställa ytterligare föreskrifter angående själva märkningen.
1. I bilagan fastställs analysmetoderna för att bestämma
c) saltinnehållet,
f) innehållet av flyktiga syror,
i) innehållet av kalciumjoner, och
Denna förordning träder i kraft den 1 juli 1986.
Enligt dessa regler är krav på importlicens eller liknande förfarande, även om de är rent formella, förbjudna i handeln mellan medlemsstaterna.
Genomförandet av en gemensam handelspolitik är ännu inte slutfört. Åtgärder från medlemsstaters sida för vissa varor från tredje land har ännu inte ersatts av enhetliga, gemensamma regler.
Enligt Europeiska enhetsakten kommer den 1 januari 1993 ett område utan inre gränser att upprättas inom vilket varor, tjänster och kapital fritt kan röra sig. Detta innebär å ena sidan att de kvarstående skillnaderna i medlemsstaternas handelspolitik gradvis kommer att försvinna eller minska, och å andra sidan att kommissionen måste vara fullt medveten om dessa mål när den bedömer behovet av att tillåta åtgärder enligt artikel 115 i fördraget. Genom kommissionens beslut 80/47/EEG av den 20 december 1979 om övervaknings- och skyddsåtgärder som medlemsstater kan tillåtas vidta för import av vissa varor med ursprung i tredje land och som har övergått till fri omsättning i någon medlemsstat(1) fastställdes vissa kriterier och förfaranden vid tillämpning av artikel 115 i fördraget.
Om en medlemsstat begär att få tillämpa skyddsåtgärder, måste fristen för utfärdande av importhandlingar förlängas om den volym som omfattas av ansökningar under prövning når en viss nivå.
Eftersom de skyddsåtgärder som har beslutats enligt artikel 115 i fördraget, inte bara utgör undantag från bestämmelserna i artiklarna 9 och 30 i fördraget, utan också hindrar upprättandet av en gemensam handelspolitik i enlighet med artikel 113 i fördraget, måste de tolkas och tillämpas strikt. Med hänsyn till detta och till de mål som har fastställts i som har fastställts i Europeiska enhetsakten bör sådana åtgärder bara tillämpas under en begränsad tid och när lägets allvar så kräver.
Artikel 1
Artikel 2
2. I regel skall kommissionen inte ge sådant tillstånd som avses i punkt 1 om
3. Utan att det påverkar tillämpningen av artikel 3, skall importhandlingen utfärdas av medlemsstaten i fråga, för varje begärd kvantitet och utan avgift, inom högst fem arbetsdagar från dagen för importörens ansökan, oberoende av var hans företag är beläget inom gemenskapen.
b) De regler som gäller för direkt import gentemot ursprungslandet och andra tredje länder, däribland i förekommande fall tullregler, importmöjligheternas storlek eller volym samt de ekonomiska överväganden på vilka reglerna är grundade.
- i alla tredje länder,
De uppgifter som krävs enligt punkterna c och d skall omfatta de två närmast föregående åren och det aktuella året. Om dessa uppgifter inte kan tillhandahållas i tid eller med den noggrannhet som krävs, skall medlemsstatens ansökan innehålla de uppgifter som finns tillgängliga.
b) Uppgift om ursprungslandet och den exporterande medlemsstaten.
- dess nummer i Gemensamma tulltaxan samt dess NIMEXE-nummer.
f) Uppgifter som styrker att varorna är i fri omsättning. Om varorna ännu inte är i fri omsättning den dag då ansökan om import görs eller om det vid den tidpunkten inte går att styrka att de är i fri omsättning, skall en importhandling utfärdas, men giltigheten begränsas till en månad efter den tidpunkt då den sökande tar emot handlingen.
1. I de fall då import till en medlemsstat av en vara som avses i artikel 1 medför ekonomiska svårigheter får medlemsstaten i fråga vidta skyddsåtgärder efter att ha fått tillstånd från kommissionen, som skall bestämma villkor och närmare regler för sådana åtgärder.
a) Den exporterande medlemsstaten.
- när den har sitt ursprung i tredje landet i fråga, med fördelning på direkt import och import av varor i fri omsättning,
- med ursprung i gemenskapen.
f) Om kommissionen begär det, de åtgärder som har vidtagits eller föreslagits för att avhjälpa situationen för den berörda sektorn.
- Fristen för utfärdande av importhandlingar skall ökas till tio arbetsdagar från den dag då importören lämnade in sin ansökan.
7. Kommissionen skall ta ställning till medlemsstatens begäran inom fem arbetsdagar efter mottagandet.
1. Som ett led i uppfyllandet av formaliteterna i samband med import av varor som är föremål för övervaknings- eller skyddsåtgärder inom gemenskapen får medlemsstatens behöriga myndigheter anmoda importören att ange ursprunget av de varor som är upptagna i tulldeklarationen eller i ansökan om en importhandling.
Artikel 6
Artikel 7
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100 i detta,
med beaktande av följande: Direktiv 70/156/EEG(3), senast ändrat genom Anslutningsakten för Spanien och Portugal, fastställde gemenskapens förfarande för typgodkännande av fordon som tillverkas i enlighet med de tekniska krav som specificerats i särdirektiv, och även förteckningen över fordonsdelar och egenskaper som ingår i dessa direktiv.
För att tillämpa förfarandet för typgodkännande på ett riktigt sätt bör kontroller av produktionens överensstämmelse även avse åtgärder som vidtagits av tillverkaren i syfte att säkerställa att fordon, särskilda tekniska enheter eller komponenter i serietillverkning överensstämmer med den godkända typen.
I de fall där det i särdirektiven föreskrivs att en särskild teknisk enhet måste förses med typgodkännandenummer behöver varje enhet inte nödvändigtvis åtföljas av ett intyg om överensstämmelse. Tillverkaren av en särskild teknisk enhet måste i varje enskilt fall tillhandahålla upplysningar om begränsningar i användningen av enheten och villkoren för dess montering.
Direktiv 70/156/EEG ändras på följande sätt:
- särskild teknisk enhet: en anordning för vilken det fastställs krav i ett särdirektiv, som är avsedd att vara en del av ett fordon och som kan vara typgodkänt särskilt men endast i samband med en eller flera, specificerade fordonstyper,
I detta direktiv avses med:
- "standardtypegodkendelse" i dansk lagstiftning,
- "homologacion de tipo" i spansk lagstiftning,
- "omologazione" eller "approvazione del tipo" i italiensk lagstiftning,
- "aprovaço de marca e modelo" i portugisisk lagstiftning,
2. Artiklarna 4 och 5 skall ersättas med följande:
a) Fordonstypen måste överensstämma med specifikationerna i det tekniska underlaget.
3. En medlemsstat som har beviljat typgodkännande skall i nödvändig utsträckning och vid behov i samarbete med behöriga myndigheter i andra medlemsstater, vidta nödvändiga åtgärder för att kontrollera att de åtgärder som avses i punkt 2 även fortsättningsvis är tillräckliga och att serietillverkade fordon överensstämmer med den godkända typen. Kontroll av att serietillverkade fordon överensstämmer med den godkända typen skall begränsas till stickprovskontroller, såvida inte annat anges i särdirektiven.
1. De behöriga myndigheterna i varje medlemsstat skall inom en månad sända en kopia av typgodkännandeintyget för varje fordonstyp som har godkänts eller vägrats godkännande till de behöriga myndigheterna i de andra medlemsstaterna.
4. Artikel 7.2 skall ersättas med följande:
5. Artikel 8 skall ersättas med följande:
Om bristande överensstämmelse konstateras skall de behöriga myndigheterna i den medlemsstat som utfärdade typgodkännandet vidta de åtgärder som beskrivs under punkt 1.
Kommissionen skall hållas informerad och, den skall vid behov, hålla erforderliga överläggningar i syfte att nå en överenskommelse."
1. EEG-typgodkännande kan, när detta uttryckligen föreskrivs i särdirektiven, även utfärdas för typer av system eller fordonsdelar som utgör en särskild teknisk enhet och för komponenter i överensstämmelse med artiklarna 3 till 9 och 14.
4. Innehavaren av ett EEG-typgodkännandeintyg, vilket, i enlighet med bestämmelserna i punkt 2, innehåller uppgifter om begränsningar i fråga om användning, skall för varje tillverkad enhet eller komponent tillhandahålla detaljerade upplysningar om dessa begränsningar och varje villkor för montering."
Artikel 2
1. Medlemsstaterna skall till den 1 oktober 1988 sätta i kraft de författningar som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
Det finns skäl att upphäva vissa av de tillfälliga undantagen från förbuden i direktivet, eftersom mindre farliga behandlingsmetoder nu finns att tillgå.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"Tillfälligt tillstånd får beviljas för en fabrik som börjar sin verksamhet enligt det program för produktionsstöd som fastställs i denna förordning. Tillståndet skall beviljas så snart en ansökan om godkännande har lämnats in enligt de i punkt 1 angivna villkoren. Giltighetstiden för det tillfälliga tillståndet får inte vara längre än till slutet av det regleringsår då det beviljades. Giltighetstiden för tillfälliga tillstånd som beviljades under regleringsåren 1984/85, 1985/86 och 1986/87 skall upphöra vid utgången av regleringsåret 1986/87."
RÅDETS FÖRORDNING (EEG) nr 678/87 av den 26 januari 1987 om tillämpningen av systemet med ursprungscertifikat som föreskrivs enligt Internationella kaffeavtalet 1983 när kvoterna är tillfälligt upphävda
med beaktande av rådets förordning (EEG) nr 288/82 av den 5 februari 1982 om gemenskapsregler för import(1), senast ändrad genom förordning (EEG) nr 899/83(2), särskilt artikel 16.1 b i denna,
Förordning (EEG) nr 3761/83(4) införde det system med ursprungsintyg som föreskrivs i Internationella kaffeavtalet 1983 när kvoterna tillämpas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
med beaktande av rådets förordning (EEG) nr 170/83 av den 25 januari 1983 om ett gemenskapssystem för bevarande och förvaltning av fiskeresurserna(),
Om en förstärkande nätkasse med denna maskstorlek används på nätredskap med en maskstorlek som är mindre än 40 millimeter har det visat sig att det bildas nätfickor, som leder till skador på fångsten beroende på tekniska problem med att få ut denna ur lyftet, vilket leder till att lyftet slits ut och rivs sönder.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fiskeresurser.
Förordning (EEG) nr 3440/84 ändras på följande sätt:
2. Artikel 6 skall ändras enligt följande:
- Punkt 3 skall ersättas med följande:
"6. En förstärkande nätkasse som är fastsatt på en trål med en maskstorlek på över 60 mm får sträcka sig högst två meter framför den bakre lyftstoppen."
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (), ändrad genom förordning (EEG) nr 3985/87 (), särskilt artikel 15.1 andra stycket i denna, och med beaktande av följande: I enlighet med artikel 15.1 andra stycket i förordning (EEG) nr 2658/87 skall kommissionen göra anpassningar av teknisk art av gemenskapens rättsakter som hänvisar till tulltaxe- eller statistiknomenklaturen. Rådets förordning (EEG) nr 2771/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för ägg () har ändrats genom kommissionens förordning (EEG) nr 4000/87 (), varvid varubeskrivningarna och de tulltaxenummer som anges i dessa anpassades i enlighet med Kombinerade nomenklaturen. Många andra förordningar om äggsektorn måste bli föremål för en teknisk anpassning varvid hänsyn skall tas till nya Kombinerade nomenklaturen som är baserad på systemet för harmoniserad varubeskrivning- och kodifiering som skall ersätta konventionen av den 15 december 1950 om nomenklaturen för klassificering av handelsvaror i tulltaxor. På grund av antalet och innehållet i de texter där en anpassning är nödvändig, bör alla förordningar som skall anpassas samlas i en ändringsförordning. I samband med denna anpassning av kommissionens förordning 164/67/EEG () bör vissa faktorer som används vid beräkningen av slusspriserna och som i nämnda förordning fortfarande anges i beräkningsenheter, uttryckas i ecu med användning av den koefficient på 1,208 953 som avses i artikel 13 i rådets förordning (EEG) nr 1676/85 (), senast ändrad genom förordning (EEG) nr 1636/87 (). HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Bilagan till kommissionens förordning nr 164/67/EEG av den 26 juni 1967 om fastställande av faktorerna för beräkning av importavgifter och slusspriser för härledda äggprodukter, senast ändrad genom förordning (EEG) nr 1775/74 (), skall ersättas med bilaga 1 till den här förordningen.
Artikel 5
Artikel 6
Bilagorna 1 och 2 till rådets förordning (EEG) nr 2773/75 av den 29 oktober 1975 om fastställande av bestämmelser för beräkning av importavgiften och slusspriset för ägg (), senast ändrad genom förordning (EEG) nr 3232/86 (), skall ersättas med bilaga 2 och 3 till denna förordning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater. ()()()
med beaktande av följande: Genom förordning (EEG) nr 1898/87 fastställs principen att beteckningarna mjölk och mjölkprodukter inte får användas för andra produkter än de som upptas i förordningens artikel 2. Ett undantag från denna princip är beteckningen på produkter vars beskaffenhet är känd genom traditionellt bruk eller beteckningar som uppenbarligen används för att beskriva en karakteristisk egenskap hos produkten.
med beaktande av rådets direktiv 71/127/EEG av den 1 mars 1971 om tillnärmning av medlemsstaternas lagstiftning om backspeglar för motorfordon(1), i dess lydelse enligt kommissionens direktiv 86/562/EEG(2), särskilt artikel 9 i detta, och
För fordon i kategori N2 med en massa över 7,5 ton har nuvarande krav även visat sig otillräckliga vad avser siktfältet längs den sida av förarhytten som är längst bort från föraren. För att råda bot på denna brist är det nödvändigt att möjliggöra montering av en närzonsbackpegel.
Artikel 1
1. Från och med den 1 januari 1989 får medlemsstaterna inte, av skäl som hänför sig till backspeglar
om backspeglarna på denna fordonstyp eller dessa fordonstyper överensstämmer med bestämmelserna i detta direktiv.
- Medlemsstaterna får vägra nationellt typgodkännande för en fordonstyp, vars backspeglar inte överensstämmer med bestämmelserna i detta direktiv.
Medlemsstaterna skall senast den 1 januari 1989 sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 99 i detta,
Direktiv 83/181/EEG bestämmer inte bara räckvidden av artikel 14.1 d i direktiv 77/388/EEG(), senast ändrat genom direktiv 84/386/EEG(), utan syftar även till upprättandet av gemenskapsregler för momsbefrielse vid slutlig införsel av varor som går utöver räckvidden av den nämnda artikeln. Dessa regler bör ändras eller kompletteras på ett sådant sätt att de åstadkommer en mer enhetlig tillämpning av detta på gemenskapsnivå.
Artikel 1
"2. Befrielse skall också beviljas när det gäller sedvanliga bröllopsgåvor som ges till en person som uppfyller de villkor som fastställs i punkt 1 av personer som har sin normala bosättningsort i ett land utanför gemenskapen. Befrielsen skall tillämpas på gåvor med ett värde av högst 200 ecu per styck. Medlemsstater får dock bevilja befrielse för mer än 200 ecu, om värdet av varje skattebefriad gåva inte överstiger 1 000 ecu."
3. I artikel 35.1 b andra strecksatsen skall orden "artikel 60.1 b" ersättas med "artikel 60".
Referenssubstanser för kvalitetskontroll av läkemedel
5. Följande tillfogas till artikel 56:
"Artikel 62
b) tjänster som erbjuds av en person som är etablerad i en annan medlemsstat, eller
Den befrielse som avses i artikel 62 skall begränsas till reklamtrycksaker som uppfyller följande villkor:
c) Trycksakerna får inte vara skickade som gruppförsändelser från samma avsändare till samma mottagare.
"s) Införsel av officiella publikationer som utgör språkrör för utförsellandet, internationella institutioner, regionala eller lokala myndigheter eller offentligrättsliga organ, som är etablerade i utförsellandet liksom av trycksaker som distribueras inför val till Europaparlamentet eller nationella val i det land från vilket trycksakerna härrör av utländska politiska organisationer som är officiellt erkända i medlemsstaterna, försåvitt publikationerna och trycksakerna har beskattats i utförsellandet och inte åtnjutit restitution av skatt vid utförsel."
1. Om inte annat sägs i artikel 83 85 skall följande varor vara skattebefriade vid införsel:
2. I punkt 1 används nedan angivna beteckningar med de betydelser som här anges:
eller vägfordon för annat särskilt ändamål än transport.
d) specialcontainer: container som är försedd med en särskilt utformad anordning för kylsystem, syrsättningssystem, system för termisk isolering eller andra system."
- Efter punkt b tillfogas följande:
"c) skattebefrielser i samband med överenskommelser som med hänsyn till principen om reciprocitet ingås med icke-medlemsländer som är avtalsslutande parter till konventionen om internationell civil luftfart (Chicago 1944) i syfte att genomföra rekommenderade praxis enligt 4.42 och 4.44 i bilaga 9 till konventionen (åttonde upplagan, juli 1980)."
Artikel 3
I artikel 2.1 i förordning (EEG) nr 3878/87 fastställs vilka morfologiska kännetecken rissorterna skall ha för att berättiga till produktionsstöd. I punkt 2 i samma artikel föreskrivs att från och med regleringsåret 1988/89 skall ingen sort berättiga till produktionsstöd som inte också har vissa kvalitativa kännetecken med avseende på klibbighet, konsistens och amylosinnehåll.
Förfarandet vid ändring av den sortlista som anges i bilaga B till förordning (EEG) nr 3878/87 bör inbegripa årliga kontroller som omfattar provtagning som gör det möjligt att genomföra de nödvändiga sortanalyserna.
Artikel 1
- En konsistens på minst 0,85 kg/cm².
Artikel 3
Artikel 4
3. Kommissionens tjänstemän skall före den 31 mars varje år meddela medlemsstaterna om analysresultaten.
med beaktande av rådets förordning (EEG) nr 2658/87(1) av den 23 juli 1978, om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan, senast ändrad genom förordning (EEG) nr 1315/88(2), särskilt artikel 9, och
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt de tillämpliga KN-nummer som anges i kolumn 2 av de skäl som anges i kolumn 3.
Artikel 1
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(2), och
Organen i de fyra producerande medlemsstaterna befinner sig inte i samma läge. På grund av administrativa och juridiska svårigheter har upprättandet av organen och organens verksamhet försenats i vissa medlemsstater. Dessa medlemsstater utnyttjade inte i tillräcklig grad de högsta belopp som var reserverade för dem under inledningsfasen, när utgifterna helt kunde debiteras gemenskapen. Den tid som denna fas omfattar bör därför förlängas med ett år utan höjning av de högsta belopp som redan är tilldelade enligt nuvarande bestämmelser.
Artikel 1.5 i förordning (EEG) nr 2262/84 skall ersättas med följande:
- För Grekland 100 % upp till högst 7 miljoner ecu.
Medlemsstaterna får, enligt villkor som skall bestämmas i enlighet med det förfarande som anges i artikel 38 i förordning nr 136/66/EEG, täcka en del av de utgifter som de själva skall bära genom avdrag från det beviljade gemenskapsstödet för olivolja.
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 118a i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
Kommissionens meddelande om dess program arbetarskyddsfrågor(4) förutsätter att direktiv antas i syfte att säkerställa arbetstagarnas säkerhet och hälsa.
Det åligger medlemsstaterna att inom sina territorier verka för förbättringar av arbetstagarnas säkerhet och hälsa; åtgärder, som vidtas för att skydda arbetstagarnas säkerhet och hälsa i arbetet bidrar även, i vissa fall, till att bibehålla hälsan och möjligen säkerheten hos personer i arbetstagarens hushåll.
För att säkerställa en förbättrad skyddsnivå måste arbetstagarna och/eller deras representanter informeras om de risker som föreligger för deras säkerhet och hälsa och om de åtgärder, som krävs för att minska eller eliminera dessa risker; de måste ha förutsättningar att medverka till att tillräckliga skyddsåtgärder vidtas genom avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis.
Arbetsgivare skall vara skyldiga att hålla sig à jour med de senaste tekniska och vetenskapliga framstegen vad gäller arbetsplatsens utformning med beaktande av de risker som är förbundna med deras verksamhet och att informera de arbetstagarrepresentanter, som enligt detta direktiv har rätt att ta del av sådan information, på ett sådant sätt att en högre skyddsnivå kan säkerställas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
2. Detta direktiv skall inte tillämpas på sådana offentliga verksamheter, där det inte kan undvikas att förhållanden som är speciella för dessa verksamheter kommer i konflikt med direktivet, exempelvis försvaret eller polisen eller viss specifik verksamhet inom civilförsvaret.
Definitioner
b) arbetsgivare, varje fysisk eller juridisk person som står i ett arbetsgivarförhållande till arbetstagare och har ansvar för företaget och/eller verksamheten,
Artikel 4
AVSNITT II ARBETSGIVARNAS SKYLDIGHETER
1. Arbetsgivaren är skyldig att svara för att arbetstagarens säkerhet och hälsa tryggas i alla avseenden som är förbundna med arbetet.
Artikel 6
Arbetsgivaren skall vara uppmärksam på behovet av att avpassa dessa åtgärder med hänsyn till ändrade omständigheter och sträva efter att förbättra de rådande förhållandena.
a) Arbetsgivaren skall utvärdera riskerna för arbetstagarnas säkerhet och hälsa, bland annat vid val av arbetsutrustning, de kemiska ämnen och preparat som används samt arbetsplatsernas utformning.
- integreras i all verksamhet och på alla nivåer inom företaget och/eller verksamheten.
d) Arbetsgivaren skall vidta lämpliga åtgärder för att säkerställa att endast de arbetstagare, som fått tillräckliga instruktioner, får tillträde till särskilt riskfyllda och farliga områden.
Artikel 7
2. De utsedda arbetstagarna skall inte på något sätt missgynnas på grund av sin verksamhet med avseende på skyddsfrågor och förebyggande arbete.
5. Under alla omständigheter skall
6. Ansvaret för åtgärder till skydd mot och förebyggande av de risker för säkerhet och hälsa, som avses i denna artikel, skall åligga en eller flera arbetstagare eller en eller flera enheter inom eller utanför företaget och/eller verksamheten.
8. Medlemsstaterna skall definiera de erforderliga färdigheter och kvalifikationer som avses i punkt 5.
Första hjälpen, brandbekämpning, utrymning, allvarlig och överhängande fara
2. I överensstämmelse med punkt 1 skall arbetsgivaren framför allt ifråga om första hjälpen och utrymning avdela de arbetstagare som behövs för att genomföra sådana åtgärder.
a) så snart som möjligt informera alla arbetstagare, som utsätts eller kan utsättas för allvarlig och överhängande fara, om risken i fråga och om vidtagna eller planerade skyddsåtgärder,
4. Arbetstagare som vid en allvarlig, överhängande och oundviklig fara lämnar sin arbetsplats och/eller ett farligt område skall inte på något sätt missgynnas på grund av detta utan skall skyddas mot alla skadliga och orättfärdiga följdverkningar i enlighet med nationell lagstiftning och/eller praxis.
Artikel 9
a) se till att det finns en riskvärdering av miljöfaktorer på arbetsplatsen, inbegripet faktorer för sådana grupper som är utsatta för speciella risker,
d) i enlighet med nationell lagstiftning och/eller praxis upprätta rapporter över arbetsolycksfall, som drabbat arbetstagarna.
Information till arbetstagarna
b) de åtgärder som vidtas i enlighet med artikel 8.2.
a) den riskvärdering samt information om de skyddsåtgärder som avses i artikel 9.1 a och b,
Artikel 11
Detta förutsätter
- avvägd medverkan i enlighet med nationell lagstiftning och/eller praxis.
b) utseende av arbetstagare enligt artikel 7.1 eller 8.2 och den verksamhet som avses i artikel 7.1,
e) den planering och uppläggning av utbildningen som avses i artikel 12.
6. I överensstämmelse med nationell lagstiftning och/eller praxis har arbetstagare och/eller arbetstagarrepresentanter rätt att vända sig till den arbetsmiljöansvariga myndigheten med klagomål, om de anser att de åtgärder som arbetsgivaren vidtagit inte är tillräckliga för att uppnå säkerhet och hälsa på arbetsplatsen.
Utbildning av arbetstagare
- förflyttning eller byte av arbete,
Utbildningen skall
2. Arbetsgivaren skall säkerställa att anställda i utomstående företag och/eller verksamheter som utför arbete för arbetsgivarens räkning har fått tillräckliga instruktioner ifråga om arbetsmiljörisker som gäller deras arbete i arbetsgivarens företag och/eller verksamhet.
Den utbildning som åsyftas i punkt 1 skall förläggas till arbetstid.
Artikel 13
Hälsokontroll
3. Hälsokontrollen kan ingå som en del av den allmänna sjukvården.
Särskilt utsatta riskgrupper skall skyddas mot de faror som speciellt berör dem.
2. Utan att det inskränker det förfarande som avses i artikel 17 i fråga om tekniska justeringar får detta direktiv och särdirektiven ändras i enlighet med artikel 118a i fördraget.
Kommitté
- den tekniska utvecklingen, ändringar i internationella regler eller specifikationer och nya rön,
Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande ärendet är.
3. Kommissionen skall anta förslaget, om det har tillstyrkts av kommittén.
Artikel 18
3. Medlemsstaterna skall vart femte år rapportera till kommissionen om den praktiska tillämpningen av bestämmelserna i detta direktiv, och om arbetsgivarnas och arbetstagarnas synpunkter.
Artikel 19
med beaktande av kommissionens förslag(),
och med beaktande av följande: När rådet antog direktiv 83/183/EEG(), förband sig rådet att enhälligt på kommissionens förslag införa bestämmelser som tillåter en avsevärd lättnad i eller rent av avlägsnande av formaliteterna för beviljande av skattebefrielser vid permanent införsel från en medlemsstat av enskildas personliga egendom. Särskilda kommittén för ett Medborgarnas Europa inbjöd i sin första rapport, som bekräftades av Europeiska rådet i Bryssel av den 29 och 30 mars 1985, kommissionen att presentera ett sådant förslag.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 2.2 b skall ersättas med följande:
- tolv månader då det gäller motorfordon (inklusive tillhörande släpvagnar), husvagnar och husbilar, nöjesbåtar och privatflygplan,
a) Punkt 1 blir punkt 1 a,
a) Orden "under en tid av minst tolv månader" i slutet av första stycket skall ersättas med "före inrättandet av andrabostaden".
a) Början av punkt 1 skall ersättas med följande:
"2. Skattebefrielse skall också beviljas för sedvanliga bröllopsgåvor till någon som uppfyller de villkor som fastställs i punkt 1 från personer som har sin normala hemvist i en annan medlemsstat än den dit införsel sker. Befrielsen skall gälla för gåvor med ett enhetsvärde av högst 350 ecu. Medlemsstaterna får dock bevilja skattebefrielse då gränsen 350 ecu överskrids förutsatt att värdet av varje skattebefriad gåva inte överstiger 1 400 ecu".
b) I punkt 2 skall hänvisningen till "artikel 2.2" ersättas med hänvisning till "artikel 2.2a".
RÅDETS DIREKTIV av den 11 december 1989 om veterinära kontroller vid handeln inom gemenskapen i syfte att fullborda den inre marknaden (89/662/EEG)
med beaktande av kommissionens förslag(1),
med beaktande av följande: Gemenskapen kommer att vidta åtgärder för att stegvis upprätta den inre marknaden under tiden fram till den 31 december 1992.
Det slutliga målet är att de veterinära kontrollerna skall utföras enbart vid avsändningsstället. För att uppnå detta krävs en harmonisering av de grundläggande krav som rör hälsoskyddet för människor och djur.
I destinationslandet skulle veterinära stickprovskontroller kunna utföras hos mottagarna. Vid allvarlig misstanke om felaktigheter skulle dock den veterinära kontrollen kunna utföras medan varorna är på väg.
Behovet av skyddsåtgärder måste uppmärksammas. Inom detta område, måste, inte minst med hänsyn till effektiviteten, ansvaret i första hand falla på den avsändande medlemsstaten. Kommissionen måste kunna vidta snabba åtgärder, särskilt genom att göra besök på platsen och vidta de åtgärder som läget kräver.
Bestämmelserna i gällande direktiv bör anpassas till de nya regler som fastställs i detta direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
2. handel: handel mellan medlemsstater med varor som avses i artikel 9.2 i fördraget,
5. officiell veterinär: den veterinär som förordnats av den behöriga centrala myndigheten i medlemsstaten.
De anläggningar som produkterna härrör ifrån skall genom kontinuerlig egenkontroll säkerställa att produkterna uppfyller de krav som uppställts i föregående stycke.
2. När transporten innefattar flera destinationer skall produkterna sammanföras till ett antal partier som svarar mot antalet destinationer. Varje parti skall åtföljas av det ovannämnda certifikatet eller dokumentet.
När produkterna förs in till gemenskapens territorium via en annan medlemsstat än någon av dem som avses ovan skall denna medlemsstat verkställa en kontroll i handlingarna av ursprunget och varornas destination i enlighet med artikel 6.1.
1. Medlemsstater från vilka varorna avsänds skall vidta de åtgärder som krävs för att säkerställa att de berörda parterna uppfyller de veterinära kraven i samtliga led av produktion, lagring, saluföring och transport av de produkter som avses i artikel 1. De skall särskilt säkerställa att
Artikel 5
När den behöriga myndigheten i den medlemsstat genom vilken varorna transiteras eller den medlemsstat till vilken varorna avsänts har fått uppgifter som ger anledning till misstanke om att gällande bestämmelser överträtts, får kontroller som innefattar kontroll av transportsättet också utföras under transporten av varor till medlemsstatens territorium.
- för en godkänd distributör som delar upp partierna eller för ett handelsföretag med många filialer, eller någon verksamhet som inte är underkastad ständig tillsyn skall den senare, innan partiet delas upp eller saluföras, kontrollera att varorna märkts och att de intyg eller dokument som avses i den första strecksatsen finns tillgängliga samt anmäla varje felaktighet eller avvikelse till den behöriga myndigheten.
2. Om gemensamma varustandarder inte fastställts genom gemenskapsregler och i det fall som avses i artikel 14 kan den mottagande medlemsstaten, utan att det påverkar tillämpningen av artikel 4 och med vederbörlig hänsyn till de allmänna bestämmelserna i fördraget, kräva att ursprungsanläggningen skall följa de regler som gäller enligt den ifrågavarande medlemsstatens nationella lagstiftning. Den medlemsstat från vilken produkterna härrör skall se till att den ifrågavarande produkten uppfyller dessa normer.
b) de skall föra ett register i vilket sådana leveranser noteras,
4. Närmare bestämmelser för tillämpning av denna artikel skall utformas i enlighet med det förfarande som fastställs i artikel 18.
1. I samband med den kontroll som företas på de platser där produkter kan införas till gemenskapens territorium från tredje land, däribland hamnar, flygplatser och gränsstationer mot tredje land, skall medlemsstaterna se till att följande åtgärder vidtas:
De produkter som avses i bilaga A får inte godkännas vid tullklarering annat än om dessa kontroller har visat att de uppfyller gemenskapens bestämmelser.
- efter enbart visuell besiktning för att fastställa att dokument och produkter stämmer överens, vidarebefordras under tullövervakning till destinationsorten, där veterinär besiktning skall utföras.
Artikel 7
Kostnader i samband med förstöring av partiet skall betalas av avsändaren eller dennes ombud.
Utöver detta får kommissionen på begäran av en medlemsstat och i enlighet med det förfarande som fastställs i artikel 17, när det uppkommer situationer som inte förutsetts av gemenskapens lagstiftning, vidta varje åtgärd som är nödvändig för att uppnå samstämmighet i medlemsstaternas handlande.
- använda dem för något annat ändamål, däribland att sända tillbaka dem efter att att ha inhämtat medgivande från den behöriga myndigheten i ursprungslandet.
Artikel 8
Om de kontroller som avses i artikel 7 visar upprepade oegentligheter, skall den behöriga myndigheten i den mottagande medlemsstaten underrätta kommissionen och de veterinära myndigheterna i de övriga medlemsstaterna.
- uppdra åt en officiell veterinär, vars namn skall finnas med på en av kommissionen på förslag av medlemsstaterna upprättad förteckning och som kan godkännas av de olika berörda parterna, för att kontrollera fakta vid den berörda anläggningen,
När dessa åtgärder vidtagits för att komma tillrätta med upprepade oegentligheter vid någon anläggning skall kommissionen debitera den berörda anläggningen alla utgifter som uppkommit genom tillämpning av strecksatserna i föregående stycke.
På begäran av någon av de två berörda medlemsstaterna - om oegentligheterna har bekräftats av experternas utlåtanden - skall kommissionen i enlighet med det förfarande som fastställs i artikel 17, vidta lämpliga åtgärder som får utsträckas till att bemyndiga medlemsstaterna att införa ett tillfälligt förbud mot införsel till sina territorier av produkter som härrör från den berörda anläggningen. Dessa åtgärder skall bekräftas eller omprövas snarast möjligt i enlighet med det förfarande som fastställs i artikel 17.
Beslut som fattats av den behöriga myndigheten i den mottagande staten skall tillsammans med en motivering delges avsändaren eller hans ombud och den behöriga myndigheten i den medlemsstat från vilken partiet avsänts.
Dessa experter skall yttra sig inom högst 72 timmar. Parterna skall avvakta expertens yttrande med vederbörlig hänsyn tagen till gemenskapens veterinära lagstiftning.
Den medlemsstat från vilken sändningen utgått skall omedelbart vidta de kontroll- och försiktighetsåtgärder som fastställs i gemenskapsreglerna, däribland särskilt fastställande av buffertzoner som avses i dessa regler eller vidta varje annan åtgärd som den finner lämplig.
De åtgärder som vidtagits av medlemsstaterna skall utan dröjsmål anmälas till kommissionen och till de övriga medlemsstaterna.
4. Kommissionen skall i samtliga fall vid första lämpliga tillfälle ta ställning till situationen på nytt i Ständiga veterinärmedicinska kommittén. Den skall besluta om vilka åtgärder som behöver tillgripas för de produkter som avses i artikel 1 och, om situationen så kräver, för de ursprungliga produkterna eller de produkter som härletts från dessa produkter i enlighet med förfarandet i artikel 17. Kommissionen skall följa läget och i enlighet med samma förfarande ändra eller upphäva de beslut som fattats alltefter vad situationen kräver.
Varje medlemsstat och kommissionen skall utse den eller de veterinärmyndigheter som skall svara för de veterinära kontrollerna och samarbetet med de andra medlemsstaternas inspektionsmyndigheter.
- verkställa inspektioner av lokaler, kontor, laboratorier, installationer, transportmedel, anläggningar och utrustning, rengörings- och underhållsmedel och de rutiner som används vid framställning, bearbetning, kontrollmärkning, märkning och presentation av dessa produkter,
- granska skriftligt eller datoriserat material som är av betydelse för de kontroller som verkställs utöver de åtgärder som vidtagits med stöd av artikel 3.1.
1. Artikel 8.3 och artiklarna 10 och 11 i direktiv 64/433/EEG(8), senast ändrat genom direktiv 88/657/EEG(9), utgår.
i) skall artiklarna 5.2, 5.3, 5.4 och 5.5 och artiklarna 6 och 8, utgå, och
5. I direktiv 80/215/EEG
6. Artikel 5.3 och 5.4 och artiklarna 7, 8 och 12 i direktiv 85/397/EEG(15), ändrat genom förordning (EEG) nr 3768/85(16), utgår.
9. I bilaga B till direktiv 72/462/EEG(18) skall följande läggas till i intyget: "Första mottagarens namn och adress".
"Artikel 19
3. Följande artikel läggs till direktiv 77/99/EEG:
"Artikel 18
Artikel 14
Rådet skall, efter förslag från kommissionen, före den 31 december 1991 fastställa de slutliga reglerna vad gäller handel med de produkter som räknas upp i bilaga B.
"2 a En eller flera kommissionsledamöter får, på begäran av en medlemsstat eller på initiativ av kommissionen själv, genast bege sig till den berörda platsen för att, i samarbete med de behöriga myndigheterna, granska de åtgärder som vidtagits och avge ett yttrande om dessa åtgärder."
2. Kommissionen skall granska de program som överlämnats av medlemsstaterna i enlighet med punkt 1.
3. Kommissionen skall själv anta förslaget om det är förenligt med yttrandet från kommittén.
Om rådet inte har fattat något beslut inom 15 dagar från det att förslaget kommit det till handa, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas, såvida inte rådet med enkel majoritet har avvisat förslaget.
2. Företrädaren för kommissionen skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. De röster som avgivits av företrädarna för medlemsstaterna skall vägas enligt samma artikel i fördraget. Ordföranden får inte rösta.
Rådet skall fatta sitt beslut med kvalificerad majoritet.
Före det datum som nämns i första stycket skall rådet med kvalificerad majoritet fatta beslut, efter förslag från kommissionen, om de regler och allmänna principer som skall gälla vid de kontroller av införsel från länder utanför gemenskapen av varor som omfattas av detta direktiv. Före detta datum skall på samma sätt kontrollstationer vid de yttre gränserna inrättas och de krav fastställas som dessa gränsstationer skall uppfylla.
Fram till den 31 december 1992 får medlemsstaterna för att tillåta gradvis införande av de kontrollarrangemang som fastställs i detta direktiv, utan hinder av artikel 5.1
Artikel 21
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv vid ett datum som skall fastställas genom det beslut som skall fattas före den 31 december 1990, i enlighet med andra stycket i artikel 19.1, dock senast den 31 december 1991.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
Då man öppnar det offentliga upphandlingsområdet för konkurrens mellan medlemsstaterna, krävs en väsentligt större garanti för insyn och icke-diskriminering. För att detta skall ha påtaglig verkan, måste snabba och effektiva rättsmedel stå till buds i händelse av överträdelse av gemenskapsrättens regler för offentlig upphandling eller av nationell lagstiftning om genomförandet av sådana regler.
Om företagen inte begär prövning, torde rättelse i vissa fall aldrig komma till stånd, såvida man inte inrättar en särskild ordning för ändamålet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Medlemsstaterna skall förhindra diskriminering mellan företag, vilka vid upphandling gör gällande skada till följd av den åtskillnad som görs i detta direktiv mellan nationella bestämmelser om införande av gemenskapsrätten och andra nationella bestämmelser.
1. Medlemsstaterna skall se till att införda bestämmelser om prövning enligt artikel 1 innefattar behörighet att
c) ge ersättning åt en person, som skadats av överträdelse.
5. Medlemsstaterna får bestämma att, i de fall skada görs gällande på grund av att beslut tillkommit i strid mot lag, det överklagade beslutet först skall upphävas av ett organ med nödvändig behörighet för detta.
7. Medlemsstaterna skall se till att införa bestämmelser, som garanterar, att granskningsorganens beslut verkligen åtlyds.
Artikel 3
3. Inom 21 dagar från mottagandet av underrättelsen enligt punkt 2 skall medlemsstaten till kommissionen avge
c) uppgift om att upphandlingsförfarandet har avbrutits, antingen på upphandlingsmyndighetens eget initiativ, eller på grundval av maktbefogenheter som givits i artikel 2.1 a.
Artikel 4
Medlemsstaterna skall före den 1 december 1991 införa de bestämmelser som är nödvändiga för att följa detta direktiv. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning och andra författningar som de antar inom det område som omfattas av detta direktiv.
med beaktande av rådets förordning (EEG) nr 2658/87(1) av den 23 juli 1987, om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan, senast ändrad genom förordning (EEG) nr 20/89(2), särskilt artikel 9 i denna, och
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt de tillämpliga KN-nummer som anges i kolumn 2 av de skäl som anges i kolumn 3.
Artikel 1
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Dessa klädesplagg är av det slag som i allmänhet bärs utanpå andra kläder och som skyddar mot vind, kyla och regn.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
med beaktande av Fördraget om upprättandet av Europeiska atomenergigemenskapen, särskilt artikel 31 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
Kommissionen framlade två meddelanden till rådet, den 14 juni respektive den 9 december 1988. De var avsedda som tillägg till bilagan till förordningen och hade utarbetats efter samråd med expertgruppen som avses i artikel 31 i fördraget.
Därför verkar det lämpligt att sammanföra gränsvärdena och andra uppgifter i denna bilaga i en enda tabell.
Artikel 1
Artikel 7 i förordning (Euratom) nr 3954/87 skall ersättas med följande:
Artikel 3
med beaktande av rådets direktiv 64/433/EEG av den 26 juni 1964 om hygienproblem som påverkar handeln med färskt kött inom gemenskapen(1), senast ändrat genom direktiv 86/587/EEG((2), särskilt artikel 13 i detta, och
De hygienkrav som föreslås a
med beaktande av följande: I enlighet med artikel 13 i direktiv 64/433/EEG och i enlighet med förfarandet i artikel 16 får på begäran undantag från punkt 45 c i bilaga 1 beviljas varje medlemsstat som lämnar liknande garantier. Vid sådana undantag skall hygienkrav som lägst motsvarar kraven i nämnda bilaga fastställas.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till förordning (EEG) nr 2658/87, är det nödvändigt att fastställa bestämmelser för klassificering av de varor som anges i bilagan till den här förordningen.
Nomenklaturkommittén har inte yttrat sig inom den tid som ordföranden bestämt vad gäller produkt nr 4 i tabellen i bilagan.
Artikel 1
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Det framgår av officiella uppgifter som Australien har tillhandahållit att den ovan nämnda skadegöraren inte förekommer där och att landet länge har upprätthållit ett strängt förbud mot import av växter och växtprodukter som kan föra med sig denna skadegörare.
Kommissionen kommer att säkerställa att Australien årligen tillhandahåller alla de tekniska uppgifter som är nödvändiga för att bedöma den ovan nämnda situationen.
Härmed förklaras att Australien erkänns vara fritt från Erwinia amylovora (Burr.) Winsl. et al. Artikel 2
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
i samarbete med Europaparlamentet(2),
Både pentaklorfenol (CAS nr 87-86-5) och dess föreningar är farliga för människan och miljön, särskilt vattenmiljön. Användningen av dessa ämnen bör regleras.
Den gällande gemenskapslagstiftning som avser medlemsstaternas rätt att besluta om mer långtgående begränsningar för användningen av de aktuella ämnena och preparaten i arbetsmiljön berörs inte av detta direktiv.
Artikel 1
Om inte annat följer av bestämmelserna i artikel 3.5 skall båtförarcertifikat för navigering på Rhen, som utfärdas i överensstämmelse med den reviderade konventionen om sjöfarten på Rhen, gälla för alla vattenvägar inom gemenskapen.
2. Medlemsstaterna skall ömsesidigt erkänna de båtförarcertifikat som fortfarande är giltiga och som är upptagna i grupp B i bilaga 1 som giltiga för navigering på deras inre vattenvägar, bortsett från dem för vilka behörighetsbeviset för navigering på Rhen erfordras eller sådana som är upptagna i bilaga 2, som om de själva hade utfärdat ifrågavarande båtförarcertifikat.
Medlemsstaterna skall erkänna det certifikat som utfärdas i enlighet med nummer 10 170 i ADNR (förordningen om transport av farligt gods på Rhen) som bevis på dessa kunskaper.
Artikel 5
Artikel 7
Kommissionen skall själv anta ändringen av bilaga 1 om den är förenlig med kommitténs yttrande.
Artikel 8
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Den definition av toleransen som fastställs i artikel 4 i förordning (EEG) nr 3492/90 för förvaring av jordbruksprodukter i offentliga interventionslager och beräkningsmetoden för bestämning av de finansiella följderna av lagring måste anges närmare.
För vissa produkter som bearbetas mellan uppköp och lagring skall särskilda toleranser fastställas för svinn i samband med bearbetning.
För vissa jordbruksprodukter har beräkningsmetoden för procentsatsen för normalt svinn i samband med lagring genomgått grundläggande förändringar. Dessa procentsatser bör därför revideras mot bakgrund av erfarenheten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE. Artikel 1
Den faktiska vikten vid inlagring och utlagring skall beräknas genom att från den registrerade vikten dra den standardvikt för förpackningen som fastställts i uppköpsvillkoren eller, i avsaknad av sådan, den genomsnittliga förpackningsvikt som används av myndigheten.
- bearbetning av tobak i blad 19 %.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: I förordning (EEG) nr 1208/81(2) fastställs gemenskapens skala för klassificering av slaktkroppar av vuxna nötkreatur.
Förordning (EEG) 1208/81 ändras på följande sätt:
1. Slaktkroppar av vuxna nötkreatur skall indelas i följande kategorier:
C. Slaktkroppar av kastrerade djur av hankön.
Utan att det påverkar gällande interventionsbestämmeler skall bokstäverna A, B, C, D och E användas för att identifiera slaktkroppar från och med den 1 januari 1992.
a) konformation,
Den konformationsklass som betecknas med bokstaven S i bilaga 1 får användas av medlemsstaterna om de vid frivilligt införande av en konformationsklass över de existerande klasserna (djur med dubbelmuskulatur) önskar att ta hänsyn till egenskaperna hos eller den förväntade utvecklingen av en viss produktion.
2. Bilaga 1 skall ersättas med den bilaga som finns i bilagan till denna förordning.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
I kommissionens förordning (EEG) nr 1014/90(2) fastställs en första omgång tillämpningsföreskrifter. Dessa behöver kompletteras.
"Artikel 7b
solbaerrom, även kallad blackcurrant rum.
KOMMISSIONENS FÖRORDNING (EEG) nr 2988/91 av den 11 oktober 1991 om ändring av förordning (EEG) nr 1538/91 om tillämpningsföreskrifter till förordning (EEG) nr 1906/90 om vissa handelsnormer för fjäderfäkött
med beaktande av rådets förordning (EEG) nr 1906/90 av den 26 juni 1990 om vissa handelsnormer för fjäderfäkött(1), särskilt artikel 9 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
RÅDETS BESLUT av den 13 juli 1992 om datorisering av veterinära förfaranden vid import (Shift-projektet), om ändring av direktiven 90/675/EEG, 91/496/EEG, 91/628/EEG och beslut 90/424/EEG och om upphävande av beslut 88/192/EEG (92/438/EEG)
med beaktande av kommissionens förslag,
Dessa nya bestämmelser skall bidra till att skydda människors och djurs hälsa samtidigt som de gör det möjligt att genomföra den inre marknaden för djur och animaliska produkter.
Direktiv 90/675/EEG, 91/496/EEG och 91/628/EEG bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Organisation och drift av databaser som innehåller import till gemenskapen av djur och produkter.
I detta beslut skall vid behov de definitioner tillämpas som återfinns i direktiv 90/675/EEG, 91/496/EEG och 91/628/EEG.
2. Det informationssystem som avses i artikel 1.1 första strecksatsen skall fungera enligt principerna i bilaga 1.
2. De databaser som avses i artikel 1.1 andra strecksatsen skall organiseras och fungera enligt principerna i bilaga 2.
2. De databaser som avses i artikel 1 tredje strecksatsen skall organiseras och fungera enligt principerna i bilaga 3.
Artikel 7
Direktiv 90/675/EEG skall ändras på följande sätt:
"d) konsultera de databaser som avses i artikel 1, andra strecksatsen i beslut 92/438/EEG."
4. Artikel 11.4 b första strecksatsen skall ersättas med följande:
"I så fall skall den behöriga myndigheten informeras via det datoriserade nätverket som länkar samman veterinärmyndigheter (Animo)."
7. I artikel 16.1 a skall den tredje strecksatsen utgå.
Artikel 9
"Kontrollen skall göras efter att man har konsulterat de databaser som avses i artikel 1 andra strecksatsen i beslut 92/438/EEG."
4. I artikel 9.1 d skall orden "som avses i artikel 12.4 andra stycket" ersättas med "som avses i artikel 20 i direktiv 90/425/EEG".
6. I artikel 12.1 c skall tredje strecksatsen utgå.
8. I artikel 30.2 första stycket skall orden "andra stycket" utgå.
Artikel 11
1. Ekonomiskt bidrag från gemenskapen kan beviljas för datorisering av veterinärförfarandena vid import enligt beslut 92/438/EEG(*).
Artikel 13
3. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande ärendet är. Kommittén skall fatta sitt beslut med en majoritet på 54 röster, varvid medlemsstaternas röster skall vägas enligt fördragets artikel 148.2. Ordföranden får inte rösta.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas och tillämpa dem omedelbart.
Artikel 15
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Kommissionen antog den 19 juli 1991 beslut 91/398/EEG om ett datoriserat system som länkar samman veterinärmyndigheterna (Animo)(3) och den 2 juli 1992 beslut 92/373/EEG om utnämnande av datacentret Animo(4).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Samordningsmyndigheten skall förhandla fram ett kontrakt med Eurokom om användning av det gemensamma datacentret. Kontraktet skall undertecknas i enlighet med nationella bestämmelser.
- gäller till den 1 juli 1995,
- innehåller en förpliktelse från Eurokom att uppfylla alla de tekniska krav som fastställs i bilagan till kommissionens beslut 91/638/EEG(5), baserade på den tekniska lösning som Eurokom föreslog i sitt anbud. Avtal om ytterligare uppgifter för Eurokom, inklusive uppgifter i samband med införande av systemet i varje medlemsstat och projektets förvaltning, skall ingås i form av separata överenskommelser,
b) Överföringskostnader som skall variera med hänsyn till tillgång eller frånvaro av ett nationellt datacentrum och som motsvarar det fördelaktigaste pris som Eurokom har kunnat erhålla från leverantören av kommunikationsutrustning.
Artikel 4
Om det under införandet av systemet uppstår en situation som, särskilt vad gäller de ekonomiska aspekterna, inte ligger i linje med detta besluts mål, skall kommissionen vidta nödvändiga åtgärder i enlighet med förfarandet i artikel 42 i rådets beslut 90/424/EEG(7).
KOMMISSIONENS DIREKTIV 92/4/EEG av den 10 februari 1992 om ändring i rådets direktiv 78/663/EEG om särskilda renhetskriterier för emulgerings-, stabiliserings-, förtjocknings- och geleringsmedel för användning i livsmedel
med beaktande av rådets direktiv 89/107/EEG av den 21 december 1988 om tillnärmning av medlemsstaternas lagstiftning om tillsatser som är godkända för användning i livsmedel(1), särskilt artikel 3.3 i detta, och med beaktande av följande:
De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga livsmedelskommittén.
Bilagan till direktiv 78/663/EEG ändras på det sätt som visas av bilagan till det här direktivet.
När en medlemsstat antar bestämmelser till följd av detta direktiv skall dessa innehålla en hänvisning till direktivet eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
RÅDETS DIREKTIV 92/32/EEG av den 30 april 1992 om ändring för sjunde gången i rådets direktiv 67/548/EEG om tillnärmning av lagar och andra författningar om klassificering, förpackning och märkning av farliga ämnen
med beaktande av kommissionens förslag(1),
med beaktande av följande: Olikheter mellan lagar och andra författningar om klassificering, förpackning och etikettering av farliga ämnen och anmälan av nya ämnen i medlemsstaterna kan leda till handelshinder mellan medlemsstater och skapa ojämlika konkurrensvillkor. Sådana skillnader mellan bestämmelserna i de olika medlemsstaterna påverkar direkt den inre marknadens funktion och har som följd att hälsa och miljö inte garanteras skydd på samma nivå.
Alla nya ämnen som släpps ut på marknaden bör anmälas till de behöriga myndigheterna, varvid vissa uppgifter lämnas. Vad beträffar ämnen som släpps ut på marknaden i mindre kvantiteter än ett ton per år och tillverkare kan lägre krav ställas. Om å andra sidan ett ämne släpps ut på marknaden i kvantiteter som överstiger vissa gränser bör kompletterande undersökningar genomföras.
Dessutom är det viktigt att noga följa utvecklingen och användningen av nya ämnen som släpps ut på marknaden. Det är därför nödvändigt att införa ett system varigenom alla nya ämnen tas upp i en förteckning.
I rådets direktiv 87/18/EEG av den 18 december 1986 om harmonisering av lagar och andra författningar om tillämpningen av principerna för god laboratoriesed och kontrollen av och tillämpningen vid prov med kemiska ämnen(9) anges gemenskapens principer för god laboratoriesed, som skall följas vid tester av kemikalier.
För att säkerställa en tillräckligt hög skyddsnivå för människan och miljön är det nödvändigt att vidta åtgärder som avser förpackning och provisorisk märkning av sådana farliga ämnen som inte finns upptagna i bilaga 1 till direktiv 67/548/EEG. Av samma anledning är det nödvändigt att göra tillhandahållandet av skyddsanvisningar obligatoriskt.
Sekretess bör garanteras för vissa uppgifter om affärs- och driftförhållanden.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) anmälan av ämnen,
2. Direktivet skall inte gälla följande preparat i bruksfärdigt skick, avsedda för slutanvändaren:
c) Ämnesblandningar som i form av avfall omfattas av direktiv 75/442/EEG(5) och 78/319/EEG(6).
f) Bekämpningsmedel.
Kommissionen skall senast 12 månader efter anmälan av detta direktiv enligt förfarandet i artikel 29.4 a upprätta en förteckning över ovan nämnda ämnen och preparat. Förteckningen skall ses över regelbundet och vid behov ändras i enlighet med nämnda förfarande.
Artikel 2
a) ämnen: kemiska grundämnen och deras föreningar i naturlig eller framställd form, inklusive eventuella tillsatser nödvändiga för att bevara produkternas stabilitet och eventuella föroreningar som härrör från tillverkningsprocessen, men exklusive eventuella lösningsmedel som kan avskiljas utan att detta påverkar ämnets stabilitet eller ändrar dess sammansättning.
d) anmälan: de handlingar med föreskrivna uppgifter som lämnats till den behöriga myndigheten i en medlemsstat enligt följande:
f) vetenskaplig forskning och utveckling: vetenskapliga experiment, analyser eller kemisk forskning som utförs under kontrollerade förhållanden. Häri innefattas fastställandet av inneboende egenskaper, verkan och effektivitet såväl som vetenskapliga undersökningar i samband med produktutveckling.
2. Med farliga avses i detta direktiv följande ämnen och preparat:
c) synnerligen brandfarliga ämnen och preparat: flytande ämnen och preparat som har ytterst låg flampunkt eller låg kokpunkt samt gasformiga ämnen och preparat som är antändbara i kontakt med luft av rumstemperatur och normalt lufttryck.
- fasta ämnen och preparat som lätt fattar eld även vid kortvarig kontakt med en antändningskälla och som fortsätter att brinna eller förbrukas även sedan kontakten med antändningskällan upphört, eller
e) Brandfarliga ämnen och preparat: flytande ämnen och preparat med låg flampunkt.
h) Hälsoskadliga ämnen och preparat: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan leda till döden eller ge akuta eller kroniska skador.
k) Sensibiliserande ämnen och preparat: ämnen och preparat som vid inandning eller upptagning genom huden kan framkalla överkänslighet, så att karakteristiska symptom uppstår vid förnyad exponering för ämnet eller preparatet.
n) Ämnen och preparat skadliga för fortplantningen: ämnen och preparat som vid inandning, förtäring eller upptagning genom huden kan orsaka eller öka förekomsten av icke ärftliga skador på avkomman eller på den manliga eller kvinnliga fortplantningsfunktionen eller -förmågan.
Tester och bedömning av ämnenas egenskaper
Laboratorieförsök skall utföras i enlighet med principerna för god laboratoriesed i direktiv 87/18/EEG och bestämmelserna i direktiv 86/609/EEG.
Klassificering
3. I bilaga 1(2) finns en förteckning över ämnen som klassificerats enligt principerna i punkt 1 och 2, med uppgift om deras harmoniserade klassificering och märkning. Beslutet att ta upp ett ämne i bilaga 1 med harmoniserad klassificering och märkning skall fattas enligt förfarandet i artikel 29.
1. Om inte annat följer av artikel 13 skall medlemsstaterna vidta alla nödvändiga åtgärder för att säkerställa att ämnen inte kan släppas ut på marknaden, som sådana eller ingående i preparat, om de inte
Dessutom skall medlemsstaterna vidta alla nödvändiga åtgärder för att säkerställa att bestämmelserna om säkerhetsdatablad i artikel 27 följs.
Undersökningsplikt
Fullständig anmälan
- En redovisning av ämnets negativa effekter inom olika tänkbara användningsområden.
- Om tillverkaren befinner sig utanför gemenskapen skall anmälaren, i enlighet med artikel 2.1 d andra strecksatsen, vid behov bifoga en förklaring från tillverkaren att anmälaren har utsetts att ensam företräda tillverkaren när det gäller att inge anmälan för ämnet i fråga.
2. Om inte annat följer av artikel 14 skall varje anmälare av ett redan anmält ämne underrätta den behöriga myndigheten
- när den mängd av ämnet som släppts ut på marknaden uppnår 1000 ton per år och tillverkare, eller när den totala mängd av ämnet som släppts ut på marknaden uppnår 5000 ton per tillverkare, varvid den behöriga myndigheten skall lägga upp ett program för tester/undersökningar enligt bilaga 8 nivå 2, som skall genomföras av anmälaren inom den tid som den behöriga myndigheten bestämmer.
Begränsade anmälningskrav för ämnen som släpps ut på marknaden i mängder under ett ton per år och tillverkare
- Alla övriga uppgifter enligt artikel 7.1.
4. Likaledes skall en anmälare som har lämnat en begränsad anmälan enligt kraven i punkt 1, lämna en fullständig anmälan enligt kraven i artikel 7 innan den mängd av ämnet som släpps ut på marknaden uppnår ett ton per år per tillverkare eller den totala mängd som släpps ut på marknaden per tillverkare uppnår fem ton
Redan anmälda ämnen (tioårsregeln)
Utsläppande på marknaden av anmälda ämnen
2. Om inte annat anges av den behöriga myndigheten, får ämnen som anmälts enligt artikel 8.1 eller 8.2 släppas ut på marknaden tidigast 30 dagar efter det att myndigheten mottagit en dokumentation som överensstämmer med kraven i detta direktiv.
Ämnen som framställs utanför gemenskapen
Polymerer
Undantagsbestämmelser
- Tillsatser och ämnen som endast används i djurfoder och omfattas av direktiv 70/524/EEG och 82/471/EEG(1).
- Ämnen som endast används i vissa andra produktkategorier för vilka gemenskapen tillämpar anmälnings- eller godkännandeförfaranden och för vilka kraven i fråga om uppgiftslämnande är likvärdiga med dem som föreskrivs i detta direktiv. Senast 12 månader efter anmälan av detta direktiv skall kommissionen i enlighet med förfarandet i artikel 29.4 a upprätta en förteckning över sådana gemenskapsregler. Denna förteckning skall regelbundet ses över och vid behov ändras enligt samma förfarande.
- Ämnen som släpps ut på marknaden i mindre mängder än 10 kg per år och tillverkare, förutsatt att tillverkaren/importören uppfyller de krav som uppställs av de medlemsstater där ämnet släpps ut på marknaden. Dessa krav får inte gå utöver vad som föreskrivs i bilaga 7 C, punkt 1 och 2.
- Ämnen som säljs till ett begränsat antal registrerade kunder för användning vid processinriktad forskning och utveckling i mängder som är begränsade till vad som krävs för den processinriktade forskningen och utvecklingen. Dessa ämnen får undantas i ett år, under förutsättning dels att tillverkaren eller importören till den behöriga myndigheten i varje medlemsstat där tillverkning, import eller processinriktad forskning och utveckling sker lämnar uppgifter om ämnenas identitet, märkningsinformation, mängder, skälen varför dessa mängder behövs samt en förteckning över kunderna och deras forsknings- och utvecklingsprogram, dels att han rättar sig efter krav som dessa myndigheter eller medlemsstaterna uppställer för sådan forskning och utveckling. De krav som medlemsstaterna uppställer får inte gå utöver vad som föreskrivs i artikel 8. Efter ett år skall anmälningsskyldighet normalt gälla för dessa ämnen. Tillverkaren eller importören skall också försäkra att ämnet eller preparatet det ingår i endast kommer att hanteras av kundens personal under kontrollerade förhållanden och inte vid något tillfälle kommer att göras tillgängligt för allmänheten, som sådant eller i ett preparat. Om den behöriga myndigheten anser att en oacceptabel risk föreligger för människan eller miljön kan myndigheten vidare föreskriva att detsamma skall gälla för produkter som innehåller de nya ämnen som framställts under den processinriktade forskningen och utvecklingen.
Om det inte är möjligt att märka ämnena fullständigt och i enlighet med principerna i artikel 23 på grund av att resultaten från testerna enligt bilaga 7 A inte är tillgängliga, bör utöver märkningen från de utförda testerna på etiketten anges "Varning - ämnet ännu inte fullständigt testat".
1. En anmälare av ett ämne som redan anmälts i enlighet med artikel 7.1 eller 8.1 skall vara skyldig att på eget initiativ skriftligen underrätta den behöriga myndighet till vilken anmälan ursprungligen lämnades om:
- nya användningsområden för vilka ämnet släpps ut på marknaden och som han rimligen kan förväntas känna till,
2. Varje importör av ett ämne framställt av en tillverkare utanför gemenskapen som importerar ämnet inom ramen för en anmälan som tidigare lämnats av en ensam företrädare i enlighet med artikel 2.1 d, skall vara skyldig att tillse att denne förses med aktuell information angående de mängder av ämnet som han släpper ut på marknaden inom gemenskapen.
1. För ett ämne som redan har anmälts i enlighet med artikel 7.1 eller 8.1, kan den behöriga myndigheten medge att den som därefter anmäler ämnet vid tillämpningen av avsnitt 3-5 i bilaga 7 A och B och avsnitt 3 och 4 i bilaga 7 c åberopar de testresultat som lämnats av den förste anmälaren, förutsatt att den andre anmälaren kan visa att det nyanmälda ämnet är identiskt med det redan anmälda, också vad beträffar renhetsgrad och föroreningar. Den förste anmälaren måste ge skriftligt tillstånd till att hans testresultat får åberopas.
b) om den första anmälarens namn och adress.
c) Den första anmälaren har inte begärt och beviljats ett tidsbegränsat undantag från denna artikel.
4. Om en anmälare och en ny anmälare av ett och samma ämne trots bestämmelserna i punkt 2 och 3 inte kan nå en överenskommelse om utbyte av information, får medlemsstaterna, i syfte att förhindra tester på ryggradsdjur, i fråga om anmälare inom deras territorier tillämpa nationella bestämmelser, som innebär att gamla och nya anmälare är skyldiga att dela på uppgiftslämnandet, och fastställa förfarandet för användningen av uppgifterna. Bestämmelserna får omfatta regler om det tidsbegränsade undantag som avses i artikel 7.1 sista strecksatsen och om en rimlig avvägning mellan berörda parters intressen.
1. Medlemsstaterna skall utse en eller flera behöriga myndigheter som skall ansvara för mottagandet av uppgifter enligt artikel 7-14 och för bedömningen av huruvida uppgifterna överensstämmer med kraven i detta direktiv.
- i kontrollsyfte ta nödvändiga prover,
I fråga om ämnen som anmälts i enlighet med artikel 7.1, 8.1 och 8.2 skall den behöriga myndighet som mottar anmälan göra en riskbedömning i enlighet med de allmänna principer som avses i artikel 3.2. Bedömningen skall omfatta rekommendationer om den lämpligaste metoden för att testa ämnet och, där så är lämpligt, rekommendationer om åtgärder i syfte att minska riskerna för människan och miljön i samband med att ämnet släpps ut på marknaden. Riskbedömningen skall regelbundet ses över med hänsyn till kompletterande uppgifter som lämnas i enlighet med denna artikel eller artikel 7.2, 8.3 och 14.1.
3. I fråga om anmälningar som lämnats i enlighet med artikel 8 skall de behöriga myndigheterna senast 30 dagar efter det att anmälan kommit in avgöra om den överensstämmer med detta direktiv och, i fall då anmälan bedöms inte överensstämma med detta direktiv, upplysa anmälaren om vilka kompletterande uppgifter som krävs för att dokumentationen skall överensstämma med direktivet. Om anmälan överensstämmer med detta direktiv skall myndigheten inom samma tid meddela anmälaren det officiella nummer som tilldelats hans anmälan.
6. Om inte annat följer av artikel 19.1 skall medlemsstaterna och kommissionen tillse att sekretess gäller för uppgifter om kommersiell utveckling och tillverkning.
När en medlemsstat mottagit den dokumentation som avses i artikel 7.1 och 8.1 eller uppgifter från kompletterande tester som utförts enligt artikel 7.2 och 8.3 eller kompletterande uppgifter som lämnats i enlighet med artikel 14, skall den till kommissionen snarast möjligt sända en kopia av dokumentationen eller av de kompletterande uppgifterna eller en sammanfattning därav.
Artikel 18
2. En behörig myndighet i en annan medlemsstat kan direkt samråda med den behöriga myndighet som mottog den ursprungliga anmälan eller med kommissionen om vissa punkter i de uppgifter som ingår i den dokumentation som föreskrivs i detta direktiv eller om den riskbedömning som avses i artikel 16.1. Den kan också föreslå att ytterligare tester eller uppgifter begärs eller att riskbedömningen omprövas. Om den behöriga myndighet som mottog den ursprungliga anmälan inte tillmötesgår de andra myndigheternas önskemål rörande kompletterande uppgifter, bekräftande tester eller ändringar av de undersökningsprogram som avses i bilaga 8, eller rörande riskbedömningen, skall den motivera sitt beslut för de berörda myndigheterna. Om myndigheterna inte kan enas och någon av myndigheterna med stöd av utförligt angivna skäl finner att kompletterande uppgifter, bekräftande tester, ändringar av undersökningsprogrammen eller en omprövning av riskerna verkligen krävs för att skydda människan och miljön, kan den begära att kommissionen fattar ett beslut i enlighet med förfarandet i artikel 29.4 b.
1. Om anmälaren anser att det finns ett sekretessproblem, kan han ange vilka uppgifter enligt artikel 7, 8 och 14 som enligt hans bedömning är kommersiellt känsliga och kan medföra skada industriellt eller kommersiellt om de lämnas ut, och som därför bör hållas hemliga för alla utom för de behöriga myndigheterna och kommissionen. En fullständig motivering måste lämnas i sådana fall.
b) tillverkarens eller anmälarens namn,
e) sammanfattningen av resultaten från toxikologiska och ekotoxikologiska tester,
Om anmälaren, tillverkaren eller importören själv senare offentliggör tidigare sekretessbelagda uppgifter, skall han meddela den behöriga myndigheten detta.
3. Ämnen som finns upptagna i förteckningen enligt artikel 21.1 och som inte är klassificerade som farliga i detta direktivs mening kan, om den behöriga myndighet som mottagit anmälan så begär, upptas under sitt handelsnamn. Normalt får sådana ämnen upptas under handelsnamnet i högst tre år. Om den behöriga myndighet som mottog anmälan anser att ett offentliggörande av det kemiska namnet i dess IUPAC-form i sig självt skulle avslöja information angående kommersiellt utnyttjande eller kommersiell framställning, kan ämnet emellertid upptas under sitt handelsnamn så länge den behöriga myndigheten anser det lämpligt.
I samtliga fall gäller att sådana uppgifter
Artikel 20
I sådana fall skall de behöriga myndigheterna i en medlemsstat och kommissionen för tillämpningen av artikel 18.2 alltid kunna ta del av anmälningshandlingarna och de kompletterande uppgifterna.
Förteckningar över existerande och nya ämnen
Förpackning
b) Materialet i förpackningen och förslutningen skall inte kunna angripas av innehållet eller bilda farliga föreningar med detta.
e) Behållare som innehåller ämnen som säljs till eller tillhandahålls allmänheten och är märkta "mycket giftigt", "giftigt" eller "frätande" enligt detta direktiv skall, oberoende av storleken, vara försedda med barnsäkra förslutningsanordningar och en varningsmärkning som kan uppfattas vid beröring.
3. Ändringar i de kategorier av ämnen vilkas förpackningar skall vara utrustade enligt punkt 1 e och 1 f skall beslutas enligt förfarandet i artikel 29.
Märkning
a) Namnet på ämnet enligt en av de benämningar som anges i bilaga 1. Om ämnet ännu inte är upptaget i bilaga 1 skall namnet anges med den internationellt vedertagna nomenklaturen.
Om mer än en farosymbol tilldelas ett ämne gäller följande:
- Om symbolen E är obligatorisk behöver inte symbolerna F och O anges.
f) EEG-nummer, när sådant tilldelats. EEG-numret erhålls från EINECS eller från den förteckning som avses i artikel 21.1.
4. Information av typen "inte giftig", "inte hälsoskadlig" eller annan liknande upplysning får inte förekomma på etiketter eller förpackningar till ämnen som omfattas av detta direktiv.
Dessa mått är endast avsedda för den information som krävs enligt detta direktiv och vid behov för kompletterande hälso- och säkerhetsinformation.
4. De i artikel 23 föreskrivna upplysningarna på etiketten skall framträda tydligt mot bakgrunden och skall vara tryckta i så stor stil och med så stora mellanrum att de är lätta att läsa.
6. Vid tillämpningen av detta direktiv skall märkningskraven anses vara uppfyllda i följande fall:
- och denna förpackning är märkt i enlighet med internationella regler om transport av farliga ämnen och enligt artikel 23.2 a, b och d-f, och
Artikel 25
Ovannämnda artiklar skall inte heller gälla bestämmelser som avser butan, propan eller gasol förrän den 30 april 1997.
b) trots bestämmelserna i artikel 23 och 24 tillåta att förpackningen för farliga ämnen som inte är explosiva, mycket giftiga eller giftiga förpackas omärkta eller märks på något annat sätt, om de innehåller så små mängder att det inte finns någon anledning anta att de som hanterar ämnet eller andra kan utsättas för fara,
3. Om en medlemsstat tillämpar något av undantagen i punkt 2 skall den genast underrätta kommissionen.
Reklam för ett ämne som tillhör en eller flera av kategorierna i artikel 2.2 skall vara förbjuden om inte de aktuella kategorierna anges i reklamen.
1. För att särskilt yrkesmässiga användare skall kunna vidta nödvändiga åtgärder till skydd för miljön samt hälsan och säkerheten på arbetsplatsen skall tillverkaren, importören eller distributören i samband med eller före den första leveransen lämna ett säkerhetsdatablad till mottagaren. Detta blad skall innehålla den information som krävs för att skydda människan och miljön.
Artikel 28
Artikel 29
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Yttrandet skall beslutas med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Rösterna från medlemsstaternas företrädare i kommittén skall vägas på det sätt som föreskrivs i artikeln. Ordföranden får inte rösta.
4. a) Utom i de fall som avses i b) skall kommissionen om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits själv besluta att de föreslagna åtgärderna skall vidtas. I det fall som avses i artikel 31.2 skall tidsfristen vara sex veckor.
Klausul om fri rörelse
Skyddsklausul
3. Om kommissionen sedan beslut fattats i enlighet med punkt 2 anser att tekniska anpassningar av bilagorna till detta direktiv krävs för fall som avses i punkt 1 ovan, skall den fatta ett beslut i frågan i enlighet med förfarandet i artikel 29.
1. Vart tredje år skall medlemsstaterna till kommissionen lämna en rapport om genomförandet av detta direktiv inom sina respektive territorier. Den första rapporten skall lämnas tre år efter genomförandet av detta direktiv.
3. Bilaga 2, 6, 7 och 8 ändras härmed enligt följande:
- Bilaga 7 ersätts av bilaga 3 till detta direktiv.
3. Direktiv 78/631/EEG:
4. Direktiv 88/379/EEG:
- I artikel 3.5 ersätts "artikel 8.2 i direktiv 67/548/EEG" med "artikel 13.3 i direktiv 67/548/EEG".
- antingen de koncentrationer som anges i bilaga 1 till direktiv 67/548/EEG för ämnet i fråga, eller
"p) Preparat skall anses behöva behandlas som skadliga för fortplantningen och tilldelas minst farosymbolen och faroangivelsen "giftigt" om de innehåller ett ämne som har sådana verkningar och som tilldelas minst en av de R-fraser enligt bilaga 6 till direktiv 67/548/EEG som betecknar ämnen som är skadliga för fortplantningen enligt kategori 2, i koncentrationer som motsvarar eller överstiger
- Artikel 3.5 q skall ha följande lydelse:
- den koncentration som anges i punkt 6 i bilaga 1 (tabell VI) till detta direktiv, om ämnet inte är upptaget i bilaga 1 till direktiv 67/548/EEG eller förekommer där, men utan angivelse av koncentrationsgränser."
- I artikel 7.1 c ii ersätts "artikel 11.4" av "artikel 19.4".
"3a De i artikel 7 föreskrivna uppgifterna på etiketten skall framträda tydligt mot bakgrunden och skall vara tryckta i så stor stil och med så stora mellanrum att de är lätta att läsa.
- I rubriken till bilaga 1, del 6 ersätts "teratogena verkningar" med "verkningar på fortplantningen".
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 oktober 1993. De skall genast underrätta kommissionen om detta.
Artikel 4
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande(),
För att snedvridningar skall undvikas förutsätter avskaffandet av dessa kontroller vad gäller mervärdesskatt inte endast en enhetlig skattebas utan även att ett flertal skattesatser och skattenivåer ligger tillräckligt nära varandra mellan medlemsstaterna. Det är därför nödvändigt att ändra direktiv 77/388/EEG().
Artikel 1
"3. a) Från och med den 1 januari 1993 skall medlemsstaterna tillämpa en normalskattesats, vilken till och med den 31 december 1996 inte får vara lägre än 15%.
b) Medlemsstaterna får tillämpa en reducerad skattesats på tillhandahållande av naturgas och elektricitet, under förutsättning att ingen risk för snedvridande verkningar på konkurrensen föreligger. En medlemsstat som avser att tillämpa en sådan skattesats skall underrätta kommissionen innan så sker. Kommissionen skall fatta beslut beträffande förekomsten av risk för snedvridning av konkurrensen. Om kommissionen inte har gjort detta inom tre månader efter mottagandet av sådan underrättelse, anses någon risk för snedvridning av konkurrensen inte föreligga.
Intill dess kan de medlemsstater som för närvarande tillämpar reducerad skattesats fortsätta att göra det; de som för närvarande tillämpar normalskattesats kan däremot inte tillämpa reducerad skattesats. Detta medger ett tvåårigt uppskov med införandet av normalskattesatsen.
2. Första meningen i artikel 12.4 skall utgå.
4. Artikel 28.2 ersätts med följande:
Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa bestämningen av egna resurser i samband med dessa operationer.
c) Medlemsstater som enligt villkoren i artikel 12.3 måste höja den normalskattesats som gällde den 1 januari 1991 med mer än 2 %, får tillämpa en reducerad skattesats som är lägre än det minimum som fastlagts i artikel 12.3 vad gäller den reducerade skattesatsen på sådana kategorier av varor och tjänster som specificeras i bilaga H. Vidare får dessa medlemsstater tillämpa en sådan skattesats på restaurangtjänster, barnkläder, barnskor och bostäder. Medlemsstaterna får inte med stöd av detta stycke införa regler om undantag med återbetalning av skatten i föregående led.
f) Grekland får tillämpa mervärdesskattesatser som är intill 30 % lägre än motsvarande skattesatser på det grekiska fastlandet i departementen Lesbos, Chios, Samos, Dodekaneserna och Cykladerna, liksom på följande öar i Egeiska havet: Thasos, Norra Sporaderna, Samothrake och Skiros.
Artikel 2
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
KOMMISSIONENS FÖRORDNING (EEG) nr 305/92 av den 7 februari 1992 om ändring av förordning (EEG) nr 410/90 om fastställande av kvalitetsnormer för kiwifrukt
med beaktande av rådets förordning (EEG) nr 1035/72 av den 18 maj 1972 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom förordning (EEG) nr 1623/91(2), särskilt artikel 2.2 andra stycket i denna, och med beaktande av följande:
För att anpassa kvalitetsnormerna för kiwifrukt till de övriga EEG-normerna för frukt och grönsaker bör det göras ändringar vad avser "hållbarhet", "storlek" och "storlekssortering".
b) Det tredje stycket under "ii) Klass I" skall i alla språkversioner ha följande lydelse:
- Ett mindre färgfel.
c) Under "iii) Klass II" skall tredje stycket fjärde strecksatsen angående "Haywardmärken ha följande lydelse:
"Storleken bestäms av fruktens vikt."
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
Det är nödvändigt att ändra bilaga V i förordning (EEG) nr 2377/90 för att beakta de ändringar som gjorts ifråga om kraven vid prövning av veterinärmedicinska produkter vilka infördes genom kommissionens direktiv 92/18/EEG av den 20 mars 1992 om ändring av bilaga till rådets direktiv 81/852/EEG om tillnärmning av medlemsstaternas lagstiftning om analytiska, farmakologiska, toxikologiska och kliniska normer och prövningsplaner för veterinärmedicinska läkemedel.
RÅDETS FÖRORDNING (EEG) nr 1764/92 av den 29 juni 1992 om ändring av ordningen för import till gemenskapen av vissa jordbruksprodukter som har sitt ursprung i Algeriet, Cypern, Egypten, Israel, Jordanien, Libanon, Malta, Marocko, Syrien och Tunisien
med beaktande av kommissionens förslag, och
För att kunna göra detta är det nödvändigt att ändra ordningen för import till gemenskapen, som omfattas av bestämmelserna i protokollen till associerings- eller samarbetsavtal med Algeriet, Cypern, Egypten, Israel, Jordanien, Libanon, Malta, Marocko, Syrien och Tunisien.
1. De tullar som gäller den 31 december i gemenskapen i dess sammansättning den 31 december 1985 för de produkter som förtecknas i bilaga II till fördraget och som har sitt ursprung i de berörda icke-medlemsländerna i medelhavsområdet och för vilka tullavveckling utsträcks till tiden efter den 1 januari 1993 enligt de protokoll till associerings- eller samarbetsavtal som finns i bilaga 1 till denna förordning skall upphävas i två lika steg från och med den 1 januari 1992 och från och med den 1 januari 1993.
RÅDETS FÖRORDNING (EEG) nr 2077/92 av den 30 juni 1992 om branschorganisationer och branschavtal inom tobakssektorn
med beaktande av kommissionens förslag(1),
med beaktande av följande: Utvecklingen på medellång och lång sikt av gemenskapens och världens jordbruksmarknader gör det nödvändigt att ompröva vissa instrument inom den gemensamma jordbrukspolitiken för att återskapa balans på marknaden. Dessa justeringar, som principiellt syftar till att skapa mera flexibla former för marknadsstödet, förutsätter att aktörerna på marknaden ändrar sitt ekonomiska beteende och tar större hänsyn till den faktiska situationen på marknaden.
För att stödja den del av branschorganisationernas verksamhet som är av särskilt intresse med tanke på de nuvarande reglerna om den gemensamma organisationen av marknaden inom tobakssektorn bör bestämmelser införas som gör det möjligt att på vissa villkor utvidga de regler som en branschorganisation antagit för sina medlemmar till att även omfatta alla producenter eller producentgrupper, även de som inte är medlemmar, i en eller flera regioner. Icke medlemmar bör också kunna vara skyldiga att betala hela eller del av den medlemsavgift som är avsedd att täcka de kostnader för nämnda verksamhet som inte avser administration. Denna ordning bör genomföras på ett sådant sätt att berörda socioekonomiska gruppers rättigheter garanteras, särskilt konsumentens rättigheter.
För att informera medlemsstaterna och andra intressenter bör det i början av varje år offentliggöras en lista över de organisationer som erkänts under det föregående året och en lista över de organisationer som fått sitt erkännande återkallat under samma period samt de bestämmelser som fått ett utvidgat tillämpningsområde med angivande av deras omfattning.
a) Medverkan till ökad samordning av avsättningen av tobak i blad och tobak i balar.
d) Ökning av produkternas förädlingsvärde, särskilt genom marknadsföringsåtgärder och forskning om nya användningsområden som inte utgör ett hot mot folkhälsan.
g) Utveckling av metoder och medel för förbättring av produktkvaliteten i produktions- och beredningsledet.
3. Medlemsstaten skall återkalla erkännandet om
c) branschorganisationen underlåter att uppfylla anmälningsplikten enligt artikel 7.2.
1. Kommissionen skall efter ansökan erkänna branschorganisationer som
c) uppfyller föreskrifterna i artikel 3.1 b d.
3. Kommissionen skall återkalla erkännandet av de organisationer som anges i punkt 1 i de fall som anges i artikel 3.3.
Artikel 6
1. Utan hinder av artikel 1 i förordning nr 26(4) skall artikel 85.1 i fördraget inte tillämpas på de avtal och samordnade förfaranden som de erkända branschorganisationerna ingått för genomförande av de åtgärder som anges i artikel 2.3.
- kommissionen inom tre månader efter det att den har erhållit alla de upplysningar som behövs inte har funnit att avtalen eller de samordnade förfarandena är oförenliga med gemenskapens bestämmelser.
- kan leda till någon form av uppdelning av marknaderna inom gemenskapen,
- innebär ett fastställande av priser eller kvoter, utan att det påverkar tillämpningen av åtgärder som branschorganisationerna vidtar till följd av särskilda bestämmelser som fastställts av gemenskapen,
Artikel 8
2. De bestämmelser, för vilka ett utvidgat tillämpningsområde begärs, skall ha tillämpats i minst ett år och avse ett av följande områden:
c) Användande av miljövänliga odlingsmetoder.
3. En utvidgad tillämpning av bestämmelserna skall godkännas av kommissionen i enlighet med det förfarande som anges i artikel 9.
De berörda intressenterna skall ha två månader på sig att lämna sina synpunkter.
4. Om de bestämmelser för vilka utvidgad tillämpning begärs är "tekniska föreskrifter" i den betydelse som anges i direktiv 83/189/EEG(5), skall de anmälas till kommissionen i enlighet med artikel 8 i det direktivet samtidigt med den i punkt 2 angivna anmälan.
Kommissionen skall under alla omständigheter avslå ansökan om den finner att den utvidgade tillämpningen
- äventyrar målen för den gemensamma jordbrukspolitiken eller andra delar av gemenskapslagstiftningen.
Artikel 10
- Forskning för att öka förädlingsvärdet på produkterna, särskilt genom nya användningsområden som inte utgör ett hot mot folkhälsan.
3. De berörda medlemsstaterna skall anmäla till kommissionen vilka beslut som de avser att fatta enligt punkt 1. Dessa beslut får träda i kraft tidigast tre månader efter tidpunkten för anmälan till kommissionen. Kommissionen får inom denna tid kräva att hela eller delar av förslaget till beslut förkastas, om det allmänna ekonomiska intresse som hävdas inte förefaller välgrundat.
Varje beslut som medlemsstaterna eller kommissionen fattar om åtgärder som innebär att enskilda eller grupper som inte är medlemmar i en branschorganisation skall betala avgift skall offentliggöras i Europeiska gemenskapernas officiella tidning. Beslutet får träda i kraft tidigast två månader efter tidpunkten för offentliggörandet.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Det har också på senare år iakttagits att konsumenterna tenderar att fästa större vikt vid livsmedlens kvalitet än kvantitet. Intresset för speciella produkter skapar en allt större efterfrågan på jordbruksprodukter och livsmedel med känt geografiskt ursprung.
Strävan att skydda jordbruksprodukter eller livsmedel som har ett känt geografiskt ursprung har gjort att vissa medlemsstater har infört registrerade ursprungsbeteckningar. Dessa har visat sig vara till gagn för producenterna som kunnat tillförsäkra sig större inkomster genom verkliga insatser för att förbättra kvaliteten, och för konsumenterna som får möjlighet att köpa högkvalitetsprodukter med garanti beträffande produktionsmetod och ursprung.
Denna förordnings räckvidd begränsas till vissa jordbruksprodukter och livsmedel där det finns ett samband mellan egenskaperna hos produkten eller livsmedlet och det geografiska ursprunget. Räckvidden kan sedermera ökas så att också andra produkter eller livsmedel omfattas.
För att en geografisk beteckning eller en ursprungsbeteckning skall åtnjuta skydd i varje medlemsstat måste den registreras på gemenskapsnivå. Registreringen skall också ge information om produkten eller livsmedlet till dem som sysslar med handel samt till konsumenterna.
Föreskrifter bör införas för handeln med tredje land som erbjuder likvärda garantier för utfärdande och kontroll av geografiska beteckningar och ursprungsbeteckningar på deras territorium.
Artikel 1
Bilaga 1 kan ändras enligt det förfarande som fastställs i artikel 15.
- som härstammar från ifrågavarande region, ort eller land,
- som härstammar från ifrågavarande region, ort eller land,
4. Trots punkt 2 a skall vissa geografiska beteckningar behandlas som ursprungsbeteckningar när råvarorna till produkterna kommer från ett vidare geografiskt område än det område där produkterna bearbetas eller från ett annat område, om
och - kontroll har ordnats av att dessa villkor iakttas.
7. För att en beteckning skall behandlas som ursprungsbeteckning enligt punkt 4, måste ansökan om registrering inges inom två år från det att denna förordning trätt i kraft.
I denna förordning avses med namn som har blivit generiskt ett namn på en jordbruksprodukt eller ett livsmedel som, visserligen har samband med den ort eller den region där produkten eller livsmedlet från början framställdes eller marknadsfördes men har blivit den allmänna benämningen på produkten eller livsmedlet i fråga.
- förhållandena i andra medlemsstater,
2. Ett namn får inte registreras som ursprungsbeteckning eller geografisk beteckning om det kommer i konflikt med namnet på en växtsort eller en djurras och därmed riskerar att vilseleda allmänheten om produktens verkliga ursprung.
1. För att en jordbruksprodukt eller ett livsmedel skall kunna få en skyddad ursprungsbeteckning (PDO) eller geografisk skyddad beteckning (PGI) måste produkten eller livsmedlet överensstämma med en produktspecifikation.
b) En beskrivning av jordbruksprodukten eller livsmedlet, med uppgift i förekommande fall om råvarorna och de viktigaste fysiska, kemiska, mikrobiologiska och/eller organoleptiska egenskaperna hos produkten eller livsmedlet.
e) En beskrivning av vilken metod som använts för framställning av jordbruksprodukten eller livsmedlet och i förekommande fall uppgift om den ursprungliga hävdvunna metoden i trakten.
h) Uppgifter om hur märkning sker med skyddad ursprungsbeteckning respektive geografisk beteckning eller jämbördiga traditionella nationella beteckningar.
2. En grupp eller en fysisk eller juridisk person får ansöka om registrering endast av jordbruksprodukter eller livsmedel som denne själv producerar eller förädlar i den mening som avses i artikel 2.2 a eller b.
5. Medlemsstaten i fråga skall kontrollera att ansökningen uppfyller de krav som uppställts i denna förordning och om den finner att så är fallet tillställa kommissionen ansökan inklusive den produktspecifikation som avses i artikel 4 jämte de övriga handlingar varpå den byggt sitt beslut.
Kommissionen skall underrätta den berörda medlemsstaten om vad den därvid har funnit.
4. Kommissionen skall i Europeiska gemenskapernas officiella tidning offentliggöra
5. Om kommissionen på basis av den granskning som föreskrivits i punkt 1 finner att namnet inte är skyddsberättigat, skall kommissionen i enlighet med det förfarande som föreskrivs i artikel 15 besluta att inte företa det offentliggörande som föreskrivs i punkt 2 i denna artikel.
1. Inom sex månader efter det offentliggörande i Europeiska gemenskapernas officiella tidning som avses i artikel 6.2, har varje medlemsstat rätt att framställa invändning mot registreringen.
4. En invändning skall upptas till behandling endast i något av följande fall:
- Invändningen visar att det namn som registreringsansökningen avser är av generisk beskaffenhet.
b) Om ingen förlikning har träffats, skall kommissionen fatta beslut i enlighet med det förfarande som föreskrivs i artikel 15, med beaktande av traditionell skälig praxis och av den faktiska risken för förväxling. Om kommissionen beslutar att fullfölja registreringsförfarandet, skall den genomföra offentliggörande i enlighet med artikel 6.4.
Artikel 9
Kommissionen får dock i enlighet med det förfarande som föreskrivs i artikel 15 besluta att vid mindre ändringar inte tillämpa det förfarande som avses i artikel 6.
2. Ett kontrollorgan kan bestå av en eller flera för uppgiften utsedda kontrollmyndigheter och/eller privata organ som har godkänts för ändamålet av medlemsstaten. Medlemsstaterna skall tillställa kommissionen förteckningar på dessa myndigheter och/eller privata organ och deras respektive befogenheter. Kommissionen skall offentliggöra dessa uppgifter i Europeiska gemenskapernas officiella tidning.
Fr. o. m. den 1 januari 1988 måste ett privat organ för att kunna godkännas av en medlemsstat för de ändamål denna förordning avser, uppfylla de krav som fastställs i standarden EN 45011 av den 26 juni 1989.
6. Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att se till, att en producent som följer denna förordning har tillgång till kontrollsystemet.
1. Varje medlemsstat har rätt att framföra anmärkning om att ett villkor som ingår i en beteckningsskyddad jordbruksprodukts eller ett beteckningsskyddat livsmedels produktspecifikation inte är uppfylld.
4. Kommissionen skall granska denna ansökan genom att rådfråga de berörda medlemsstaterna. Kommissionen skall när så är lämpligt höra den kommitté som avses i artikel 15. Kommissionen skall därefter vidta de åtgärder som är nödvändiga. Till dessa kan höra att registreringen avförs.
- Tredje land är berett att ge skydd likvärt det som är tillgängligt inom gemenskapen för motsvarande jordbruksprodukter eller livsmedel som härstammar från gemenskapen.
Artikel 13
b) Varje obehörigt bruk, imitation eller anspelning, även när produktens verkliga ursprung anges eller det skyddade namnet har översatts eller åtföljs av uttryck som "stil", "typ", "metod", "sådan som tillverkas i", "imitation" eller dylikt.
När det i en registrerad beteckning ingår en benämning på en jordbruksprodukt eller ett livsmedel och denna benämning anses generisk, skall det inte anses strida mot reglerna i punkt a eller b ovan att använda denna generiska benämning om jordbruksprodukten eller livsmedlet i fråga.
- att märkningen klart anger produktens verkliga ursprung.
Artikel 14
Denna punkt skall också tillämpas när ansökan om registrering av varumärke ingivits före dagen för offentliggörande av den registreringsansökan som föreskrivs i artikel 6.2 under förutsättning att detta offentliggörande skedde innan varumärket registrerades.
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen varvid medlemsstaternas röster skall vägas enligt nämnda artikel. Ordföranden får inte rösta.
Om rådet inte fattat något beslut inom tre månader från det att saken hänskjutits till rådet, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 17
3. Medlemsstaterna får bibehålla det nationella skyddet för de beteckningar som de har meddelat i enlighet med punkt 1 intill dess att beslut om registrering i enlighet med denna förordning har fattats.
KOMMISSIONENS FÖRORDNING (EEG) nr 2145/92 av den 29 juli 1992 om en omformulering vad avser de destinationszoner som skall användas vid fastställandet av exportbidrag, exportavgifter och vissa exportlicenser för spannmål och ris
med beaktande av rådets förordning (EEG) nr 2727/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för spannmål(1), senast ändrad genom förordning (EEG) nr 1738/92(2), särskilt artikel 16.6 i denna,
De politiska förändringarna i östblocket, dvs. upplösningen av Sovjetunionen och Jugoslavien i oberoende stater, gör det nödvändigt att aktualisera den förteckning över destinationszoner som anges i bilagan till förordning (EEG) nr 1124/77. I den bilagan bör "Sovjetunionen" och "Jugoslavien" ersättas med namnen på de nybildade stater som tidigare ingick i Sovjetunionen och Jugoslavien. Dessutom bör det ske en omgruppering av staterna i område I, II, III och VIII när möjligheten nu bjuds.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Förordning (EEG) nr 1124/77 skall upphöra att gälla.
KOMMISSIONENS FÖRORDNING (EEG) nr 2221/92 av den 31 juli 1992 om ändring av förordning (EEG) nr 1274/91 om tillämpningsföreskrifter för förordning (EEG) nr 1907/90 om vissa handelsnormer för ägg
med beaktande av rådets förordning (EEG) nr 1907/90 av den 2 juni 1990 om vissa handelsnormer för ägg(1), särskilt artiklarna 10.3, 20.1 och 22.2 i denna, och med beaktande av följande:
Det valfria angivandet av produktionssystem bör begränsas till de termer som anges i förordning (EEG) nr 1274/91, med undantag för organiska eller biologiska produktionssystem. För att underlätta kontroller i hela gemenskapen bör förteckningarna över registrerade producenter utväxlas mellan medlemsstaterna och förpackningsanläggningar bör föra veckoregister över lager med klassificerade ägg.
En positiv vikttolerans bör införas för att säkerställa en rättvis konkurrens mellan aktörerna.
- Artikel 1.6, andra strecksatsen, skall ersättas med följande text:
2. Aktören får vid förpackningstillfället ange värpdagen på förpackningen, varvid värpdagen även skall anges på de ägg som förpackningen innehåller. Värpdagen får emellertid även stämplas på äggen på produktionsföretaget.
- dagen, från 01 till 31
1 Förpackningsanläggningar skall föra separata register över
2 De producenter som avses i punkt 1 skall därefter kontrolleras regelbundet. De skall föra löpande register över
- antalet ägg eller vikten på de ägg som levererats och på vilka man avser ange värpdagen, eller på vilka produktionsföretaget redan har stämplat värpdagen, uppdelade efter köpare, och med angivande av deras namn och adress samt förpackningsanläggningens nummer.
- producentens namn, adress och nummer samt en kodad hänvisning till det hönshus från vilket äggen kommer,
5 För förpackningsanläggningar som får leveranser från egna produktionsenheter som är belägna på samma ställe och där äggen inte förpackats i slutna behållare, skall äggen
- levereras till andra förpackningsanläggningar eller industrin på värpdagen eller, om värpdagen infaller på en annan dag än arbetsdag, den första därpå följande arbetsdagen.
- de dagliga kvantiteter ägg som de mottar, uppdelade efter producenter och på vilka man avser ange värpdagen, eller på vilka produktionsföretaget redan har stämplat värpdagen, med angivande av producentens namn och adress samt registreringsnummer,
7 De produktionsenheter och förpackningsanläggningar som avses i punkt 1 skall kontrolleras minst en gång varannan månad."
"Inga andra termer än dem som anges här nedan får användas för att på ägg av klass 'A' och på små förpackningar innehållande sådana ägg ange de produktionssystem som avses i artikel 10.3 i förordning (EEG) nr 1907/90, med undantag för organiska och biologiska produktionssystem, och dessa termer får endast användas om de tillämpliga villkoren enligt bilaga 2 är uppfyllda."
"De förpackningsanläggningar som avses i punkt 2 skall föra separata register över den dagliga kvalitets- och viktklassificeringen samt försäljningen av ägg och små förpackningar som är märkta i enlighet med punkt 1, inbegripet köparens namn och adress, antalet förpackningar, antalet sålda ägg och/eller vikten på de ägg som sålts per viktklass och leveransdag, liksom veckoregister över lager med klassificerade ägg. I stället för att föra försäljningsregister kan de emellertid arkivera fakturor eller följesedlar på vilka finns angivet de uppgifter som avses i punkt 1."
6 Artikel 24 skall ersättas med följande:
Med undantag för det fall som avses i artikel 13.3 i förordning (EEG) nr 1907/90, skall vid kontroll av ett parti ägg av klass `A` en tolerans medges med hänsyn till vikten per ägg. Ett sådant parti får innehålla högst 12 % ägg vars vikt gränsar till den på förpackningen angivna vikten och högst 6 % ägg av närmast lägre viktklass.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Genom kommissionens förordning (EEG) nr 2342/92(3) skärptes kontrollbestämmelserna i fråga om import från tredje land och beviljande av exportbidrag för renrasiga nötkreatur och upphävdes förordning (EEG) nr 1544/79.
Artikel 1
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artiklarna 113 och 235 i detta,
Kommissionen, biträdd av företrädare för medlemsstaterna, skall företräda gemenskapen i den gemensamma kommitté som inrättas i enlighet med artikel 13 i avtalet.
RÅDETS DIREKTIV 93/35/EEG av den 14 juni 1993 om ändring för sjätte gången av direktiv 76/768/EEG om tillnärmning av medlemsstaternas lagstiftning om kosmetiska produkter
med beaktande av kommissionens förslag(1),
med beaktande av följande: De juridiska oklarheterna i direktiv 76/768/EEG(4), särskilt i artiklarna 1 och 2, bör undanröjas.
I fråga om färdiga kosmetiska produkter bör det fastställas vilka upplysningar som skall hållas tillgängliga för kontrollmyndigheterna på tillverkningsstället eller på den plats dit de först importerats inom gemenskapen. Dessa upplysningar skall innefatta alla nödvändiga uppgifter om identitet, kvalitet, säkerhet för människors hälsa och om de verkningar den kosmetiska produkten uppges ha.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Artikel 1.1 skall ersättas med följande:
Det faktum att varningstexter av detta slag förekommer skall dock inte befria någon från skyldigheten att iaktta de övriga kraven i detta direktiv."
Om inte tillräckliga framsteg har uppnåtts i utvecklingen av tillfredsställande metoder som kan ersätta djurförsök, särskilt i sådana fall då alternativa provningsmetoder, trots att alla rimliga ansträngningar har gjorts, inte har kunnat valideras vetenskapligt som likvärdiga i fråga om skyddsnivån för konsumenterna med beaktande av OECD:s riktlinjer för toxicitetstester, skall kommissionen senast den 1 januari 1997 lämna förslag till åtgärder för att uppskjuta det datum då denna bestämmelse skall träda i kraft under rimlig tid, och i vart fall minst två år, i enlighet med det förfarande som fastställs i artikel 10. Kommissionen skall rådfråga Vetenskapliga kommittén för kosmetologi, innan den lämnar sådana förslag.
"Artikel 5a
Denna inventering skall delas upp i två avdelningar: en för parfym och aromatiska råvaror och en för övriga ämnen.
- beståndsdelens normala funktion(er) i den färdiga produkten,
5. I artikel 6.1 skall den inledande meningen ersättas med följande:
"d) Särskilda försiktighetsåtgärder som skall iakttas vid användning, i synnerhet sådana som anges i spalten "Villkor för användning och varningstexter som skall tryckas på etiketten" i bilagorna 3, 4, 6 och 7, som skall förekomma på behållare och förpackning tillsammans med eventuell information om försiktighetsåtgärder för kosmetiska produkter som används i yrkesmässig verksamhet, särskilt av frisörer. Om detta är ogörligt av praktiska skäl, skall denna information finnas på en bipacksedel, bifogad etikett, tejp eller kort och konsumenten skall hänvisas till denna information genom att antingen en förkortad upplysning eller den symbol som anges i bilaga 8 skall förekomma på behållaren och förpackningen."
g) En förteckning över beståndsdelar i fallande ordning efter vikt då de tillsätts produkten. Denna förteckning skall föregås av ordet "innehåll". Om detta är ogörligt av praktiska skäl, skall uppgift om beståndsdelarna finnas på en bipacksedel, bifogad etikett, tejp eller kort och konsumenten skall hänvisas till denna information genom att antingen en förkortad upplysning eller den symbol som anges i bilaga 8 skall förekomma på behållaren och förpackningen."
- Kompletterande tekniskt material som används vid framställningen men som inte förekommer i slutprodukten.
I fråga om kosmetiska produkter som används i estetiskt syfte och som förekommer i flera nyanser får samtliga färgämnen som används i hela färgskalan nämnas i förteckningen, om uttrycket "kan innehålla" läggs till.
8. Följande två stycken skall läggas till sist i artikel 6.1:
9. Följande skall läggas till sist i artikel 6.3:
"2. De kan dock kräva att de uppgifter som anges i artikel 6.1 b-6.1 d och 6.1 f skall avfattas åtminstone på deras nationella eller officiella språk. De får även kräva att de uppgifter som anges i artikel 6.1 g skall avfattas på ett språk som konsumenterna kan förstå utan svårighet. Kommissionen skall därför i enlighet med förfarandet i artikel 10 fastställa en gemensam nomenklatur för beståndsdelar."
Varje medlemsstat skall utse en behörig myndighet och sända uppgifter om detta till kommissionen, som skall offentliggöra denna information i Europeiska gemenskapernas officiella tidning."
1. Tillverkaren eller dennes representant eller den person för vars räkning en kosmetisk produkt tillverkas eller den som är ansvarig för att en importerad kosmetisk produkt släpps ut på gemenskapsmarknaden skall i förebyggande syfte hålla följande information omedelbart tillgänglig för de behöriga myndigheterna i den medlemsstat det gäller på den adress som anges i märkningen enligt artikel 6.1 a:
c) Tillverkningsmetoden, som skall överensstämma med god tillverkningssed enligt gemenskapslagstiftning eller, om tillämplig sådan saknas, enligt lagstiftningen i den berörda medlemsstaten. Den person som är ansvarig för tillverkningen eller för den första importen till gemenskapen skall ha sådana yrkesmässiga kvalifikationer eller sådan erfarenhet som krävs i lagstiftning och praxis i den medlemsstat där tillverkningen eller den första importen sker.
e) Namn på och adress till den eller de experter som ansvarar för den bedömning som avses i d. Sådana experter skall ha ett examensbevis enligt definitionen i artikel 1 i direktiv 89/48/EEG i farmaci, toxikologi, dermatologi, medicin eller liknande ämne.
2. Den bedömning av säkerheten för människors hälsa som avses i punkt 1 d skall utföras enligt den princip om god laboratoriesed som fastställs i rådets direktiv 87/18/EEG av den 18 december 1986 om harmonisering av lagar och andra författningar om tillämpningen av principerna för god laboratoriesed och kontrollen av tillämpningen vid prov med kemiska ämnen(*).
5. Medlemsstaterna skall utse de behöriga myndigheter som avses i punkterna 1 och 4 och sända uppgifter om dessa till kommissionen som skall offentliggöra denna information i Europeiska gemenskapernas officiella tidning.
14. Bilaga 8, som återges i bilagan till detta direktiv, skall läggas till.
2. Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att säkerställa att sådana produkter som avses i punkt 1 inte kan säljas eller avyttras till konsumenter efter den 31 december 1997.
När en medlemsstat antar sådana bestämmelser skall dessa innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
Vidare innehåller direktiv 93/40/EEG(8) bestämmelser för den fortsatta administrationen av godkännanden för försäljning, som medlemsstaterna har meddelat efter yttrande från Kommittén för veterinärmedicinska läkemedel enligt direktiv 87/22/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att följa detta direktiv med verkan från och med den 1 januari 1995. De skall genast underrätta kommissionen om detta.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av kommissionens förslag(1),
med beaktande av följande: I rådets direktiv 74/577/EEG(4) fastställs bestämmelser om bedövning av djur före slakt.
Det är därför nödvändigt att fastställa gemensamma miniminormer för skydd av djur vid tidpunkten för slakt eller avlivning för att säkerställa en rationell utveckling av produktionen och för att underlätta genomförandet av den inre marknaden för djur och animalieprodukter.
Bestämmelserna bör även säkerställa ett tillfredsställande skydd vid tidpunkten för slakt eller avlivning av djur som inte omfattas av konventionen.
Direktiv 74/577/EEG bör upphöra att gälla.
- tekniska eller vetenskapliga experiment i samband med förfarandena i punkt 1, vilka utförs under tillsyn av en behörig myndighet,
4. Fasthållning: Varje metod som tillämpas för att begränsa djurets rörelseförmåga i syfte att underlätta bedövning eller avlivning.
7. Slakt: Avlivning av djur genom avblödning.
Artikel 3
Artikel 4
1. Hovdjur, idisslare, svin, kaniner och fjäderfä som förs till slakterier för att slaktas skall
c) bedövas före slakt eller avlivas omedelbart i enlighet med bilaga C,
3. Medlemsstaternas behöriga myndigheter kan under iakttagande av fördragets allmänna bestämmelser vad gäller anläggningar som omfattas av undantag enligt artikel 4 och artikel 13 i direktiv 64/433/EEG, artikel 4 i direktiv 91/498/EEG och artikel 7 och artikel 18 i direktiv 71/118/EEG, avstå från att tillämpa punkt 1 a vad gäller kreatur, och från punkt 1 a samt metoderna för bedövning och slakt i bilaga C vad gäller fjäderfä, kaniner, svin, får och getter, under förutsättning att kraven som fastställs i artikel 3 uppfylls.
2. Lämplig reservutrustning och reservinstrument skall finnas på slaktplatsen att användas i nödsituationer. De skall underhållas och besiktigas regelbundet.
Den behöriga myndigheten skall säkerställa att personer som arbetar med slaktning har nödvändig yrkesskicklighet och yrkesmässigt kunnande.
KAPITEL III Slakt och avlivning utanför slakterier
2. Medlemsstaterna kan emellertid bevilja undantag från punkt 1 beträffande fjäderfä, kaniner, svin, får och getter som slaktas eller avlivas utanför slakterier av sin ägare för dennes personliga bruk, under förutsättning att artikel 3 efterlevs och att svin, får och getter först blir bedövade.
2. Djur som uppföds för pälsens skull skall avlivas i enlighet med bilaga F.
Artikel 9 och artikel 10 skall inte tillämpas beträffande djur som i en nödsituation måste avlivas omedelbart.
KAPITEL IV Slutbestämmelser
2. a) Bilagorna till detta direktiv skall ändras av rådet på förslag från kommissionen i enlighet med förfarandet i punkt 1, i synnerhet för att anpassa dem till den tekniska och vetenskapliga utvecklingen.
- andra gaser än de som avses i bilaga C eller kombinationer av dessa som används vid avlivning,
c) Trots vad som sägs i a, och senast den 31 december 1995, skall kommissionen i enlighet med förfarandet i artikel 16 lämna in en rapport till Ständiga veterinärkommittén, som utarbetats på grundval av ett yttrande från Vetenskapliga veterinärmedicinska kommittén, tillsammans med relevanta förslag för fastställande av
d) I avvaktan på att b och c skall genomföras skall nationella bestämmelser på området fortsätta att gälla under iakttagande av fördragets allmänna bestämmelser.
Kommissionen skall underrätta medlemsstaterna om resultaten av kontrollerna.
4. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 16.
För att kött skall få importeras från tredje land skall det hälsointyg som åtföljer köttet kompletteras med ett intyg som visar att ovanstående krav har uppfyllts.
2. Kommissionens representant skall förelägga kommittén ett utkast till de åtgärder som skall vidtas. Kommittén skall avge ett yttrande om utkastet inom den tid som dess ordförande fastställt beroende på hur brådskande ärendet är. Yttrandet skall avges av den majoritet som fastställs i artikel 148.2 i fördraget beträffande beslut som rådet skall anta på kommissionens förslag. Medlemsstaternas representanters röster skall vägas på det sätt som anges i samma artikel. Ordföranden skall inte delta i omröstningen.
Om rådet inte har fattat beslut före utgången av en period på tre månader från den dag då saken förelades dem, skall de föreslagna åtgärderna antas av kommissionen utom då rådet har uttalat sig mot de aktuella åtgärderna med enkel majoritet.
Artikel 18
2. Från och med den dag som fastställs i punkt 1 får medlemsstaterna, under iakttagande av fördragets allmänna bestämmelser, inom sina områden upprätthålla eller tillämpa mer restriktiva bestämmelser än de som omfattas av detta direktiv. De skall underrätta kommissionen om alla sådana åtgärder.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av följande: Det är nödvändigt att anta tillämpningsföreskrifter för förordning (EEG) nr 3911/92, som bl.a. föreskriver inrättandet av en exportlicensordning för vissa kategorier av kulturföremål som anges i bilagan till den förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 3
3. Formulären skall tryckas och fyllas i på ett av gemenskapens officiella språk, bestämt av de behöriga myndigheterna i den utfärdande medlemsstaten. De behöriga myndigheterna i den medlemsstat där formuläret uppvisas får begära att det översätts till det officiella språket eller ett av de officiella språken i den medlemsstaten. I så fall skall översättningskostnaderna bäras av innehavaren av licensen.
- för att vidta nödvändiga åtgärder för att undvika att formulären förfalskas. De sätt för identifiering som antas av medlemsstaterna för detta ändamål skall anmälas till kommissionen för att vidarebefordras till de behöriga myndigheterna i de andra medlemsstaterna.
Artikel 4
3. När en sändning innehåller ett antal kulturföremål är det de behöriga myndigheterna som skall bestämma om en eller flera exportlicenser bör utfärdas för sändningen i fråga.
- ett exemplar märkt nr 1 skall utgöra ansökan,
Artikel 6
- dokumentation som innehåller alla relevanta upplysningar om kulturföremålen och deras rättsliga status vid tidpunkten för ingivande av ansökan, i förekommande fall med hjälp av stödjande handlingar (fakturor, expertvärderingar etc),
5. För att exportlicens skall beviljas skall de vederbörligen ifyllda formulären läggas fram för de behöriga myndigheter som utsetts av medlemsstaterna enligt artikel 2.2 i grundförordningen. När myndigheten har beviljat exportlicens skall exemplar 1 behållas av den myndigheten och de återstående exemplaren återsändas till innehavaren av exportlicensen eller till dennes representant.
- Det exemplar som är avsett för innehavaren av licensen.
2. Efter att ha fyllt i fält 19 B skall det tullkontor som är behörigt att ta emot exportdeklarationen återsända det exemplar som är avsett för innehavaren av licensen till deklaranten eller dennes representant.
1. Exportlicensens giltighetstid får inte överstiga tolv månader räknat från utfärdandedagen.
Artikel 10
Denna förordning träder i kraft den 1 april 1993.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Enligt rådets förordning (EEG) nr 845/72 av den 24 april 1972 om särskilda åtgärder för att främja silkesodling(2), senast ändrad genom förordning (EEG) nr 2059/92(3), beviljas stöd för de lådor med silkesfjärilsägg som ger upphov till en lyckad maskodling. Den tidpunkt när det ekonomiska målet har uppnåtts kan därför normalt anses vara den 1 augusti varje regleringsår. Detta datum kan därför användas som den avgörande händelsen för den jordbruksomräkningskurs som skall tillämpas på stöd för odling av silkesmask.
Enligt artikel 11.1 i förordning (EEG) nr 1068/93 skall den jordbruksomräkningskurs som gäller i början av regleringsåret tillämpas på hektarstödet för lin och hampa. I artikel 10.3 i samma förordning fastställs att den avgörande faktorn för stöd för privat lagring av lin- och hampfibrer skall vara den dag när kontraktet för varje enskilt parti börjar gälla. Förordningarna (EEG) nr 876/75 och (EEG) nr 1426/86 kan därför upphävas.
Artikel 2
Förordning (EEG) nr 876/75 och förordning (EEG) nr 1426/86 skall upphöra att gälla.
KOMMISSIONENS FÖRORDNING (EEG) nr 2040/93 av den 27 juli 1993 om fastställande av storleken på produktionsstöd för matpotatis på Madeira och storleken på produktionsstöd för sättpotatis och endiver på Azorerna, som fastställts i ecu av rådet och reducerats till följd av centralkursjusteringar
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas avseende den gemen-samma jordbrukspolitiken(1), särskilt artikel 9.1 i denna, och
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för utsäde.
Det stöd som avses i artiklarna 16 och 27 i förordning (EEG) nr 1600/92, och som har sänkts i enlighet med artikel 2 i förordning (EEG) nr 3824/92, fastställs till 494 ecu per hektar.
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag, och
Leveranser av bortsorterade ägg bör begränsas till sådana livs-medelsindustriföretag som godkänts i enlighet med rådets direktiv 89/437/EEG av den 20 juni 1989 om hygien-och hälsoproblem som påverkar tillverkningen och utsläppandet på marknaden av äggprodukter(3), för att säkerställa att sådana ägg hanteras korrekt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Artikel 4.1 a skall ersättas med följande:
4. Artikel 7 a skall ersättas med följande:
"a) Namnet eller firmabeteckningen och adressen till det företag som har förpackat äggen eller låtit förpacka dem; namn, firmanamn eller varumärke som används av det företaget och som kan vara ett varumärke som används gemensamt av ett antal företag, får anges om det inte innehåller någon kommentar eller symbol som är oförenlig med denna förordning i fråga om äggens kvalitet eller färskhet, typen av produktionssystem som används vid produktionen eller äggens ursprung."
7. Artikel 10.2 e skall ersättas med följande:
"2. När det gäller lösviktsförsäljning av ägg skall kontrollnumret på den förpackningsanläggning som klassificerade äggen anges eller, i fråga om importerade ägg, det tredje land där äggen har sitt ursprung liksom datum för minsta hållbarhetstid, åtföljt av lämpliga förvaringsinstruktioner."
Artikel 3
RÅDETS FÖRORDNING (EEG) nr 2847/93 av den 12 oktober 1993 om införande av ett kontrollsystem för den gemensamma fiskeripolitiken
med beaktande av kommissionens förslag(),
För att nå detta mål måste ett sådant system innehålla föreskrifter för kontroll av att åtgärderna för bevarande och förvaltning av fiskeresurserna, strukturåtgärderna och åtgärderna avseende en gemensam marknadsorganisation genomförs; det måste också innehålla vissa bestämmelser om sanktioner ifall åtgärderna inte genomförs omfattande hela fiskerisektorn, från producenten till konsumenten.
Erfarenheten från tillämpningen av rådets förordning (EEG) nr 2241/87 av den 23 juli 1987 om vissa åtgärder för kontroll av fisket() visar att det är nödvändigt att skärpa kontrollen av tillämpningen av föreskrifterna för bevarande av fiskeresurserna.
För att kunna övervaka alla fångster och landningar måste medlemsstaterna kontrollera den verksamhet som gemenskapens fiskefartyg bedriver i alla marina farvatten, samt all annan verksamhet som är förknippad med denna och har på så vis möjlighet att granska tillämpningen av bestämmelserna för den gemensamma fiskeripolitiken.
Genom att medlemsstaterna i samarbete med kommissionen genomför pilotprojekt som kan tillämpas på vissa kategorier av fartyg, kan rådet före den 1 januari 1996 avgöra om det finns anledning att införa ett övervakningssystem via satellit eller något annat system.
Det är viktigt att vid landningen närmare klargöra och bekräfta uppgifterna i loggböckerna; de personer som har hand om landningen och avsättningen av fångsterna måste därför anmäla vilka mängder som landats, lastats om, bjudits ut till försäljning eller köpts.
Begränsningar av fångsterna måste förvaltas såväl på medlemsstats- som gemenskapsnivå. Medlemsstaterna bör registrera landningarna och anmäla dem till kommissionen på elektronisk väg. Undantag från denna skyldighet måste därför kunna göras för små mängder som landas, emedan en elektronisk överföring i sådana fall skulle innebära en oproportionerligt stor administrativ och ekonomisk belastning för medlemsstaternas myndigheter.
För att hantera insamlingen och behandlingen av uppgifterna behöver databaser upprättas som särskilt gör det möjligt att samköra data. Kommissionen och dess inspektörer bör därför ha tillgång till dessa databaser på elektronisk väg för att kunna granska dem.
Det är nödvändigt att gottgöra den skada som en medlemsstat lidit som inte har förbrukat sin kvot, tilldelning eller andel av ett bestånd eller grupp av ett bestånd när fisket stoppas till följd av att en TAC är förbrukad. Av denna anledning bör ett kompensationssystem införas.
Ett av huvudsyftena med den gemensamma fiskeripolitiken är att anpassa fångstkapaciteten till de tillgängliga resurserna. Enligt artikel 11 i förordning (EEG) nr 3760/92 är det rådets uppgift att lägga fast mål och strategier för en omläggning av fiskeansträngningen. Det är också nödvändigt att se till att åtgärderna rörande den gemensamma marknadsorganisationen respekteras, särskilt av de personer som berörs av dem. Det är därför av avgörande betydelse att varje medlemsstat, utöver de finansiella kontroller som redan finns föreskrivna i gemenskapsbestämmelserna, gör tekniska kontroller för att se till att de av rådet fastställda bestämmelserna följs.
De åtgärder som vidtas till följd av överträdelserna kan variera från ett land till ett annat, vilket får fiskarna att känna sig orättvist behandlade. Frånvaron av avskräckande straffpåföljder i några medlemsstater minskar kontrollernas effektivitet. Följaktligen bör medlemsstaterna vidta nödvändiga icke diskriminerande åtgärder för att förebygga och beivra oegentligheter, särskilt genom att införa ett straffsystem som effektivt berövar lagöverträdarna det ekonomiska utbytet av överträdelserna.
För vissa åtgärder som avses i denna förordning är det lämpligt att fastställa tillämpningsföreskrifter.
Förordning (EEG) nr 2241/87 bör upphävas, med undantag av artikel 5 som fortfarande gäller fram till dess att de listor som avses i artikel 6.2 i denna förordning antagits.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- åtgärderna avseende den gemensamma organisationen av marknaden,
Artikel 2
Medlemsstaterna skall anmäla till kommissionen vilka åtgärder som vidtagits för att säkerställa att dessa förfaranden följs.
Artikel 3
Medlemsstaterna får samtidigt genomföra pilotprojekt för att utvärdera användningen av automatiska anordningar för positionsregistrering.
1. Varje medlemsstat skall själv och för egen räkning genomföra den i artikel 2 angivna inspektionen och övervakningen med hjälp av ett inspektionssystem som medlemsstaten själv fastlägger.
Artikel 5
b) det förfarande som inspektörer och befälhavare på fiskefartyg skall följa när en inspektör vill göra ett besök ombord,
e) märkning och identifiering av fiskefartygen och deras fiskeredskap,
h) det system som skall tillämpas med avseende på de fiskefartyg som för ett tredje lands flagg för att ge upplysning om deras rörelser och vilka fiskeprodukter de har ombord.
2. De arter som i enlighet med punkt 1 skall antecknas i loggboken är de arter som omfattas av TAC:er eller kvoter samt övriga arter som finns på de listor som rådet antar med kvalificerad majoritet på förslag av kommissionen.
5. Rådet kan på kommissionens förslag med kvalificerad majoritet besluta om andra undantag än det som avses i punkt 4.
7. Befälhavarna på gemenskapens fiskefartyg skall registrera de uppgifter som avses i punkterna 1 och 3, antingen i maskinläsbar form eller på papper.
1. Den befälhavare på ett fiskefartyg inom gemenskapen som önskar använda landningsställen vilka är belägna i en annan medlemsstat än flaggmedlemsstaten skall minst två timmar i förväg till de behöriga myndigheterna i denna medlemsstat anmäla
2. Den befälhavare enligt punkt 1 som underlåter att göra anmälan kan bli utsatt för lämpliga sanktioner av de behöriga myndigheterna.
1. Befälhavarna på sådana fiskefartyg inom gemenskapen som har en största längd av minst 10 m, eller deras ställföreträdare, skall efter varje resa inom 48 timmar efter landningen lämna in en deklaration till de behöriga myndigheterna i den medlemsstat där landningen äger rum. Befälhavaren är ansvarig för deklarationens riktighet, som minst skall innehålla uppgift om de landade mängderna av varje art som avses i artikel 6.2 och i vilket område de fångats.
Varje medlemsstat skall därför utarbeta en provtagningsplan och sända den till kommissionen. Resultaten av de kontroller som görs skall regelbundet meddelas kommissionen.
1. De auktionsinrättningar eller andra av medlemsstaterna bemyndigade organ som ansvarar för den första saluföringen av de fiskeprodukter som landas i en medlemsstat skall vid första försäljningstillfället lämna in en avräkningsnota, för vars riktighet dessa organ skall ansvara, till de behöriga myndigheterna i den medlemsstat på vars territorium den första saluföringen sker. Detta ansvar omfattar bara den information som avses i punkt 3.
- Individuell storlek eller vikt för varje art, samt kvalitet, produktform och färskhet.
- Såväl säljarens som köparens namn.
- Distriktsbeteckning och namn på det fiskefartyg som landat ifrågavarande produkter.
5. Avräkningsnotorna som avses i punkt 1 skall inom 48 timmar efter försäljningen översändas till medlemsstaternas behöriga myndigheter eller andra bemyndigade organ, antingen på elektronisk väg eller på papper.
Dessa undantag får bara beviljas om medlemsstaten ifråga har infört ett godtagbart kontrollsystem.
Artikel 10
c) Befälhavaren på ett fiskefartyg som för ett tredje lands flagg eller är registrerat i ett tredje land skall minst 72 timmar i förväg anmäla till de behöriga myndigheterna i den medlemsstat vars landningsplatser han önskar utnyttja vid vilken tid han avser att anlöpa landningshamnen.
2. Kommissionen får enligt förfarandet i artikel 36, under en begränsad tid som kan förlängas, undanta vissa kategorier av fiskefartyg från ett tredje land från deras förpliktelse enligt punkt 1 c, eller fastställa en annan anmälningsfrist, där hänsyn tas till bland annat avstånden mellan fiskebankarna, landningsplatserna och hamnarna i vilka fartygen ifråga är registrerade eller förtecknade.
1. Utan att det påverkar tillämpningen av artiklarna 7, 8 och 9, skall befälhavaren på ett gemenskapsfartyg som
vid omlastningen eller landningen underrätta den medlemsstat vars flagg hans fartyg för eller i vilket fartyget är registrerat om gällande arter och mängder och datumet för omlastningen eller landningen samt fångstplatsen med hänvisning till det minsta område för vilket en TAC eller kvot fastställts.
När en omlastning eller en rad omlastningar ägt rum skall mottagarfartygets befälhavare inom 24 timmar lämna in dessa uppgifter till ovannämnda behöriga myndigheter.
3. Medlemsstaterna skall vidta nödvändiga åtgärder för att kontrollera riktigheten av de uppgifter som erhållits enligt punkterna 1 och 2 och i förekommande fall överlämna dessa uppgifter och resultaten av granskningen till den eller de medlemsstater där mottagarfartyget och det fartyg varifrån omlastning sker är registrerade, eller vars flagg de för.
Om omlastningen eller landningen beräknas ske mer än 15 dagar efter fångsten skall de upplysningar som krävs enligt artiklarna 8 och 11 senast 15 dagar efter fångsten överlämnas till de behöriga myndigheterna i den medlemsstat där fartyget är registrerat eller vars flagg det för.
2. Detta dokument skall innehålla uppgifter om
c) fiskmängderna (i kg beredd vikt) för varje transporterad art, namnet på avsändaren och platsen och datumet för lastningen.
a) Dokumentet enligt punkt 1 ersätts med en kopia av en av de deklarationer som avses i artiklarna 8 eller 10 i fråga om de transporterade mängderna.
6. Varje medlemsstat skall göra stickprovskontroller på sitt territorium för att undersöka om förpliktelserna enligt denna artikel uppfylls.
1. Medlemsstaterna skall se till att alla landningar som äger rum i en medlemsstat enligt artiklarna 8, 9 och 10 registreras. De kan därför kräva att den första saluföringen sker genom offentlig auktion.
4. De medlemsstater som omfattas av undantaget i punkt 3 skall utarbeta en provtagningsplan för att bedöma storleken på de fångster som landats i de olika berörda hamnarna. Denna plan skall ha godkänts av kommissionen innan något undantag får göras. Medlemsstaten skall regelbundet sända resultaten av dessa bedömningar till kommissionen.
En sådan anmälan till kommissionen skall innehålla uppgift om fångstplatsen enligt artiklarna 6 och 8 samt om de berörda fiskefartygens nationalitet.
2. Kommissionen skall hålla de upplysningar som den tagit emot enligt denna artikel tillgängliga för medlemsstaterna genom dataöverföring.
Artikel 16
2. På kommissionens anmodan skall den medlemsstat där landningen äger rum, fångsten för första gången bjuds ut till försäljning eller där omlastningen sker sända in dessa upplysningar till kommissionen, samtidigt som den sänder dem till den medlemsstat där fartyget är registrerat.
2. Kontrollåtgärderna skall säkerställa att ägarna eller befälhavarna uppfyller följande förpliktelser:
- Flaggmedlemsstaten skall närmare underrättas om alla omlastningar av fisk till fiskefartyg från tredje land och om landningar som sker direkt i tredje land.
1. Varje medlemsstat skall före utgången av den första månaden i varje kvartal på elektronisk väg anmäla till kommissionen vilka mängder som tagits i de farvatten som anges i artikel 17 och som landats under föregående kvartal, samt lämna kommissionen alla de upplysningar som erhållits i enlighet med artikel 17.2.
3. Före den 1 oktober varje år skall kommissionen se till att medlemsstaterna får tillgång till den information som den erhållit enligt denna artikel.
2. För att underlätta denna granskning skall varje medlemsstat upprätta en elektronisk databas, där sådana data som avses i punkt 1 registreras.
4. En medlemsstat som beviljats sådana undantag skall under en tid av tre år föra ett icke elektroniskt register över de uppgifter som avses i punkt 1 och upprätta en provtagningsplan, som skall godkännas av kommissionen, så att en kontroll av uppgifternas riktighet skall kunna göras på platsen. Kommissionen skall på eget initiativ kunna företa granskningar på platsen för att kunna utvärdera provtagningsplanens effektivitet.
Artikel 20
a) Nätredskapen, vikterna och liknande utrustning skall lösgöras från trålborden, sveplinorna, trålvarpen och repen.
Varje ändring av en tidigare använd maskstorlek, liksom av fångstsammansättningen ombord vid tidpunkten för denna ändring skall därför skrivas in i loggboken och landningsdeklarationen. I speciella fall skall närmare bestämmelser om hur en stuvningsplan över bearbetade produkter för varje art skall utarbetas och hållas uppdaterad antas i enlighet med det förfarande som fastställs i artikel 36, med angivande av produkternas placering under däck.
b) speciella regler skall gälla för användningen av nät med olika maskstorlek vid speciella typer av fiske.
2. Varje medlemsstat skall fastställa ett datum när fångsterna ur ett kvoterat bestånd eller en kvoterad grupp av bestånd, som tagits av sådana fiskefartyg som för dess flagg eller är registrerade i den staten skall anses ha förbrukat den kvot som den tilldelats för detta bestånd eller denna grupp av bestånd. Från detta datum skall den tills vidare förbjuda nämnda fartyg att fiska ur detta bestånd eller denna grupp av bestånd och att bevara ombord, omlasta och landa fisk som fångats efter detta datum, och fastställa ett datum fram till vilket det är tillåtet att lasta om och landa fångster eller lämna in de senaste fångstdeklarationerna. Denna åtgärd skall omgående anmälas till kommissionen, som sedan skall informera de övriga medlemsstaterna om den.
Gemenskapens fiskefartyg skall upphöra med att fiska en art ur ett bestånd eller en grupp av bestånd som omfattas av en kvot eller TAC den dag när den kvot som tilldelats denna stat för beståndet eller gruppen av bestånd ifråga anses vara förbrukad, eller den dag när TAC:en för de arter som utgör detta bestånd eller denna grupp av bestånd anses vara förbrukad; dessa fartyg skall också upphöra med att bevara ombord, lasta om, landa eller låta lasta om eller landa fångster ur de bestånd eller grupper av bestånd som tagits efter denna dag.
Tillämpningsföreskrifter för denna punkt skall fastställas i enlighet med det förfarande som anges i artikel 36, särskilt beträffande bestämningen av ifrågavarande mängder.
Flaggmedlemsstaten skall meddela kommissionen och de övriga medlemsstaterna namnet och distriktsbeckningen på det fartyg som underkastats sådan ytterligare kontroll.
2. Rådet skall på kommissionens förslag med kvalificerad majoritet anta avdragsbestämmelser i enlighet med de mål och förvaltningsstrategier som anges i artikel 8 i förordning (EEG) nr 3760/92, och skall då i första hand ta hänsyn till följande parametrar:
- De berörda beståndens biologiska tillstånd.
Artikel 25
b) Anpassning av fiskekapaciteten genom temporärt eller definitivt stopp.
e) Utveckling av vattenbruket och kustområdena.
1. Tillämpningsföreskrifter för artikel 25 kan antas i enlighet med det förfarande som anges i artikel 36, särskilt med avseende på kontrollen av
c) fiskefartygens stillaliggandeperiod,
Artikel 27
- den landningsdeklaration som avses i artikel 8,
3. De åtgärder som avses i artikel 19.3, 19.4 och 19.5 skall tillämpas.
1. För att säkerställa att de tekniska aspekterna av de föreskrifter om åtgärder som fastställs i förordning (EEG) nr 3759/92 av den 17 december 1992 om den gemensamma organisationen av marknaden för fiske- och vattenbruksprodukter() följs skall varje medlemsstat på sitt territorium organisera regelbundna kontroller av alla dem som berörs av tillämpningen av dessa åtgärder.
b) prisreglering, särskilt vid
Medlemsstaterna skall göra jämförelser mellan dokumenten avseende den första saluföringen av de mängder som anges i artikel 9 och de landade mängder som dokumenten anger, särskilt med avseende på deras vikt.
4. Denna artikel skall inte inverka på de nationella bestämmelserna om sekretess vid rättsligt förfarande.
Inför besök på platsen skall kommissionen utfärda skriftliga instruktioner åt sina inspektörer med angivande av deras befogenhet och ändamålet med deras uppdrag.
Om kommissionen eller dess ombud stöter på svårigheter under genomförandet av sina uppdrag, skall medlemsstaterna ställa medel till kommissionens förfogande så att den kan slutföra sin uppgift, och de skall ge inspektörerna möjlighet att utvärdera kontrollerna ifråga.
Vid inspektioner till havs eller från luften är fartygets eller flygplanets befälhavare ensam ansvarig för inspektionen med hänsyn till dennes myndigheters skyldighet att tillämpa denna förordning. De av kommissionens inspektörer som deltar i inspektionen skall följa de regler och den praxis som befälhavaren fastställer.
Efter denna kontroll skall kommissionen sända en utvärderingsrapport om programmet till den berörda medlemsstaten och eventuellt rekommendera den att vidta åtgärder för att förbättra genomförandet av kontrollerna.
Om de nationella bestämmelserna föreskriver sekretess under förundersökningen får denna information inte lämnas ut utan tillstånd från den behöriga juridiska instansen.
2. Om kommissionen finner att oegentligheter begåtts vid tillämpningen av denna förordning eller att de existerande kontrollmetoderna och kontrollbestämmelserna inte är effektiva, skall den meddela den eller de berörda medlemsstaterna, som då skall sätta igång en administrativ undersökning, i vilken tjänstemän från kommissionen kan delta.
3. När kommissionens inspektörer deltar i en undersökning skall denna alltid ledas av medlemsstatens tjänstemän. Kommissionens tjänstemän får inte på eget initiativ använda sig av de inspektionsbefogenheter som tilldelats de nationella inspektörerna. Men de skall ha tillgång till samma lokaler och handlingar som dessa inspektörer.
Artikel 31
3. Påföljderna av det rättegångsförfarande som avses i punkt 2 kan beroende på brottets allvar omfatta
- beslag av fartyget,
4. Bestämmelserna i denna artikel får inte hindra landnings- eller omlastningsmedlemsstaten från att överlåta den rättsliga uppföljningen av en överträdelse på de behöriga myndigheterna i registreringsmedlemsstaten, om denna samtycker till det, förutsatt att en sådan överlåtelse skapar bättre förutsättningar för att uppnå det resultat som avses i punkt 2. Landnings- eller omlastningsmedlemsstaten skall anmäla varje sådan överlåtelse till kommissionen.
2. Om landnings- eller omlastningsmedlemsstaten inte är densamma som flaggmedlemsstaten, och de behöriga myndigheterna inte i enlighet med sin nationella lagstiftning vidtar lämpliga åtgärder, inbegripet förvaltnings- eller straffrättsliga åtgärder mot de ansvariga fysiska eller juridiska personerna, eller inte överlåter den rättsliga uppföljningen i enlighet med artikel 31.4, får den mängd fisk som olovligen landats eller lastats om skrivas av från den medlemsstatens kvot.
Artikel 33
3. Flagg- eller registreringsmedlemsstaten skall omgående anmäla till kommissionen vilka åtgärder som vidtagits i enlighet med punkt 2, samt det berörda fartygets namn och distriktsbeteckning.
De skall varje år anmäla alla ändringar av böternas minimi- och maximibelopp för varje typ av överträdelse, samt alla andra slag av tillämpliga påföljder.
Artikel 35
När förfarandet i denna artikel skall tillämpas, skall ordföranden hänskjuta ärendet till Förvaltningskommittén för fiske och vattenbruk som inrättats genom förordning (EEG) nr 3760/92, nedan kallad "kommittén", antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat.
Rådet får fatta ett annat beslut med kvalificerad majoritet inom den tid som anges i föregående stycke.
2. Namnen på de fysiska eller juridiska personerna skall bara meddelas kommissionen eller en annan medlemsstat i de fall det uttryckligen anges i denna förordning, eller om det är nödvändigt för att förebygga eller beivra överträdelser eller granska uppenbara överträdelser.
4. De uppgifter som lämnas eller tas emot i en eller annan form med stöd av denna förordning omfattas av tystnadsplikt och skall åtnjuta samma skydd som liknande uppgifter åtnjuter, såväl genom den nationella lagstiftningen i de medlemsstater som tar emot uppgifterna som genom motsvarande bestämmelser som är tillämpliga på gemenskapens institutioner.
Denna artikel påverkar inte de skyldigheter som följer av internationella konventioner om ömsesidigt bistånd i straffrättsliga frågor.
9. Uppgifterna i denna förordning skall bevaras på ett sådant sätt att de berörda personerna bara kan identifieras under den tid som behövs för ändamålet ifråga.
Denna förordning skall gälla utan att det påverkar tillämpningen av eventuella nationella kontrollåtgärder som sträcker sig utanför minimikraven, under förutsättning att de är förenliga med gemenskapsrätten och den gemensamma fiskeripolitiken.
1. Förordning (EEG) nr 2241/87 skall upphöra att gälla den 1 januari 1994 med undantag för artikel 5, som skall fortsätta att gälla till dess förordningarna om utarbetande av de förteckningar som avses i artikel 6.2 i denna förordning har trätt i kraft.
Denna förordning träder i kraft den 1 januari 1994.
KOMMISSIONENS FÖRORDNING (EEG) nr 3063/93 av den 5 november 1993 om tillämpningsföreskrifter för rådets förordning (EEG) nr 2019/93 angående stödordningen för produktion av kvalitetshonung
med beaktande av rådets förordning (EEG) nr 2019/93 av den 19 juli 1993 om införandet av särskilda bestämmelser för de mindre Egeiska öarna rörande vissa jordbruksprodukter(1) särskilt artikel 12.4 i denna,
För att uppmuntra honungsproducenter som är medlemmar av organisationer, som överensstämmer med definitionen i rådets förordning (EEG) nr 1360/78 av den 19 juni 1978 om producentgrupper och sammanslutningar av dessa(3), senast ändrad genom förordning (EEG) nr 746/93(4) att förbättra sina saluföringssystem för att tillmötesgå marknadens krav och att främja kvalitetsprodukter, är beviljande av stöd avhängigt att producenterna genomför årliga initiativprog-ram, som godkänns av de myndigheter som Grekland har utsett. För att uppnå målen bör programmet vara inriktat dels på genetiska förbättringar, omställning av bikupor, mekanisering och löpande utbildning för biodlare i ny produktionsteknik, dels på marknadsundersökningar, forskning om nya förpacknings-metoder och säljfrämjande åtgärder.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommitttén för ägg.
Stödet till produktion av den kvalitetshonung som är specifik för de mindre Egeiska öarna och som innehåller en stor andel timjanhonung, betalas ut till grupper av honungsproducenter som är erkända enligt förordning (EEG) nr 1360/78, och som genomför initiativprogram för att förbättra villkoren för saluföring och marknadsföring av kvalitetshonung.
1. Initiativprogrammet skall ha följande mål:
- Främjande av försäljningen av kvalitetshonung genom marknadsundersökningar, utveckling av nya förpackningsmetoder, samt anordnande av och deltagande i varumässor och andra säljfrämjande åtgärder.
1. Stödansökan skall lämnas in till den behöriga myndigheten under den period som dessa fastställer, dock senast den 30 september varje år, när det gäller produktionen för följande år. Vid för sen inlämning sänks stödet med 20 %, utom i fall av force majeure. Om ansökan inlämnas mer än 20 dagar efter den ansökningsperiod som fastställts av den behöriga myndigheten, skall inget stöd betalas ut.
- Sammanslutningens eller biodlarens namn och adress.
3. När det totala antalet bikupor för vilka det ansöks om stöd överstiger det högsta tillåtna antalet bikupor enligt artikel 12.3 i förordning (EEG) nr 2019/93, skall den behöriga myndigheten fastställa en schablonmässig koefficient för sänkning av alla stödbelopp.
För år 1993 får emellertid stödet betalas ut senast den 28 februari 1994.
- Antal producentsammanslutningar och antal individuella biodlare som inkommit med stödansökningar.
- De initiativprogram som blivit godkända.
Artikel 6
Artikel 7
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande (),
Det är nödvändigt att utvidga tillämpningen av förordning (EEG) nr 2299/89 och klargöra dess bestämmelser, och dessa åtgärder bör vidtas på gemenskapsnivå för att säkerställa att förordningens syften uppnås i alla medlemsstater.
Icke-regelbunden lufttrafik är av stor betydelse i gemenskapens territorium.
Det är önskvärt att likadana produkter behandlas på samma sätt och att säkerställa en rättvis konkurrens mellan de båda typerna av lufttransportprodukter samt en opartisk spridning av information till konsumenten.
Det bör klargöras att förordning (EEG) nr 2299/89 bör tillämpas på de datoriserade bokningssystem som erbjuds till eller används av alla slutkonsumenter, antingen de är enskilda personer eller företag.
Om moderföretag vägrar att ge samma information om tidtabeller, biljettpriser och platstillgång till andra system än deras eget och vägrar ta emot bokningar från dessa system kan det allvarligt snedvrida konkurrensen mellan datoriserade bokningssystem.
Ett moderföretag kan i konkurrensen mellan lufttrafikföretag få orättvisa fördelar av att det kontrollerar sitt datoriserade bokningssystem. Därför är det nödvändigt med en fullständigt lika behandling av moderföretag respektive deltagande lufttrafikföretag i den utsträckning som ett moderföretag använder de tjänster i dess eget system som omfattas av denna förordning.
Fakturorna bör innehålla tillräckligt med information för att deltagande lufttrafikföretag och abonnenter skall kunna kontrollera sina kostnader. För att underlätta en sådan kontroll bör sådan information göras tillgänglig på magnetiska medier.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Denna förordning skall gälla för datoriserade bokningssystem i den utsträckning som de omfattar lufttransportprodukter som erbjuds eller används inom gemenskapens territorium, oavsett
P den geografiska belägenheten av de flygplatser mellan vilka lufttransporten äger rum.
a) separat lufttransportprodukt: lufttrafik för befordran av passagerare mellan två flygplatser, inklusive bitjänster och ytterligare förmåner som erbjuds till försäljning och/eller säljs som en integrerad del av lufttransporttjänsten.
d) regelbunden lufttrafik: en serie flygningar, där varje flygning uppfyller följande kriterier:
1. enligt en utgiven tidtabell, eller
f) datoriserat bokningssystem: ett datoriserat system som innehåller information om bland annat lufttrafikföretags
P biljettpriser, och
P att reservera platser eller
g) distributionstjänster: tjänster som en systemleverantör ställer till en abonnents eller konsuments förfogande för att förmedla information om lufttrafikföretags tidtabeller, platstillgång, biljettpriser och tjänster i samband med flygbefordran samt för att reservera platser och/eller utställa biljetter och för att tillhandahålla andra tjänster i samband härmed.
j) effektiv kontroll: ett förhållande som bygger på rättigheter, avtal eller andra grunder, som antingen var för sig eller tillsammans och med hänsyn till faktiska omständigheter och berörda rättsregler, ger en möjlighet att direkt eller indirekt utöva ett avgörande inflytande över ett företag, i synnerhet genom
k) deltagande lufttrafikföretag: ett lufttrafikföretag som har ett avtal med en systemleverantör om förmedling av sina lufttransportprodukter genom ett datoriserat bokningssystem. I den utsträckning som ett moderföretag använder tjänsterna i sitt eget datoriserade bokningssystem, som omfattas av denna förordning, betraktas det som ett deltagande lufttrafikföretag.
n) primär textbild: en textbild som ger omfattande och opartisk information om flygförbindelser mellan två orter inom en angiven tidsperiod.
Artikel 3
b) En systemleverantör får inte ställa som villkor för att få delta i leverantörens datoriserade bokningssystem att ett deltagande lufttrafikföretag inte samtidigt deltar i ett annat system.
4. Om en systemleverantör avser att förbättra de distributionstjänster han erbjuder eller den utrustning som används i samband med att dessa tjänster erbjuds, skall han erbjuda samtliga deltagande lufttrafikföretag, inklusive moderföretag, information om och möjlighet att få del av dessa förbättringar med samma skyndsamhet, på samma villkor och under samma förutsättningar med förbehåll för de tekniska begränsningar som ligger utanför systemleverantörens kontroll, och på ett sådant sätt att det inte är någon skillnad i tidsförloppet för genomförandet av de nya förbättringarna mellan moderföretag och deltagande lufttrafikföretag."
1. a) Ett moderföretag får inte diskriminera ett konkurrerande datoriserat bokningssystem genom att vägra att ge det senare, på begäran och med samma skyndsamhet, samma information om tidtabeller, biljettpriser och platstillgång avseende dess egna flygförbindelser, som det ger sitt eget datoriserade bokningssystem, eller att vägra distribuera sina lufttransportprodukter genom ett annat datoriserat bokningssystem, eller att vägra acceptera eller med samma skyndsamhet bekräfta en bokning som görs från ett konkurrerande datoriserat bokningssystem avseende dess egna lufttransportprodukter som det distribuerar genom sitt eget datoriserade bokningssystem. Moderföretaget skall bara vara förpliktat att acceptera och bekräfta de bokningar som överensstämmer med dess biljettpriser och villkor.
2. Skyldigheten enligt denna artikel skall inte gälla till förmån för ett konkurrerande datoriserat bokningssystem när, det enligt förfarandena i artikel 6.5 eller 7.3 och 7.4 har konstaterats att det datoriserade bokningssystemet bryter mot artikel 4a eller att en systemleverantör inte kan ge tillräckliga garantier för att skyldigheterna enligt artikel 6 om moderföretags obehöriga tillgång till information uppfylls."
2. En systemleverantör får inte reservera någon specifik dataladdnings- eller databehandlingsmetod eller någon annan distributionstjänst för ett eller flera av sina moderföretag.
1. b) En systemleverantör får inte avsiktligt eller av oaktsamhet visa oriktig eller vilseledande information i sitt datoriserade bokningssystem.
1. c) Vid presentation på en primär textbild får vid sammanställning och val av flygningar mellan två givna orter ingen diskriminering göras mellan flygplatser som betjänar samma ort.
3. När en systemleverantör lämnar information om biljettpriser skall textbilden vara opartisk och icke-diskriminerande och minst innehålla biljettpriserna för alla deltagande lufttrafikföretags flygningar som visas i den primära textbilden. Källan för sådan information skall vara godtagbar för de berörda deltagande lufttrafikföretagen och systemleverantörerna.
Artikel 6
b) Varje upplysning om avsättning, bokningar och försäljning skall ske på grundval av följande:
iii) Att alla förfrågningar om sådana uppgifter skall behandlas med samma omsorg och skyndsamhet, med förbehåll för den överföringsmetod som det enskilda lufttrafikföretaget väljer.
4. Systemleverantören skall inom tre månader efter denna förordnings ikraftträdande på begäran ställa till förfogande för alla deltagande lufttrafikföretag en utförlig beskrivning av de tekniska och administrativa åtgärder som han vidtagit för att uppfylla bestämmelserna i denna artikel.
"1. Förpliktelserna för en systemleverantör enligt artikel 3 och 4 P6 gäller inte mot ett moderföretag i ett tredje land, i den mån det företagets datoriserade bokningssystem utanför gemenskapens territorium inte erbjuder EG-lufttrafikföretag en behandling som är likvärdig med den som tillämpas enligt denna förordning och enligt kommissionens förordning (EEG) nr 83/91 ().
"5. b) Om rådet, på begäran av en medlemsstat, inte inom två månader efter kommissionens beslut beslutar annorlunda, skall kommissionens beslut träda i kraft."
3. Ett lufttrafikföretags villkor för att godkänna en resebyrå som sin agent med rätt att sälja och utställa biljetter för företagets lufttransportprodukter skall inte påverka tillämpningen av punkterna 1 och 2."
I sådana fall skall en systemleverantör bara ha rätt att få tillbaka de direkta kostnaderna för uppsägningen av avtalet.
a) att en primär textbild tillhandahålls för varje enskild transaktion enligt artikel 5, utom när en konsument begär information om endast ett lufttrafikföretag, eller när en konsument begär information om endast kombinerade lufttransportprodukter,
10. I artikel 10 skall punkterna 1 och 2 ersättas med följande:
P Typ av bokning i det datoriserade bokningssystemet.
P Identifieringskod för IATA/ARC agentur.
P Bokningsdatum (transaktionsdatum).
P Statuskod (bokningsstatus).
Fakturainformationen skall erbjudas på magnetiska medier.
11. Artikel 21 skall ersättas med följande:
12. Följande artikel skall införas:
2. Systemleverantören skall informera deltagande lufttrafikföretag och kommissionen om kontrollantens identitet minst tre månader innan utnämningen bekräftas och minst tre månader före varje årlig återutnämning. Om något av de deltagande lufttrafikföretagen inom en månad efter detta meddelande ifrågasätter kontrollantens förmåga att genomföra sina uppgifter enligt denna artikel, skall kommissionen inom ytterligare två månader och efter samråd med kontrollanten, systemleverantören och varje annan part som hävdar ett legitimt intresse besluta om kontrollanten skall ersättas."
1. Denna förordning inskränker inte tillämpningen av nationell lagstiftning om säkerhet, allmän ordning eller dataskydd.
"Artikel 23
15. Bilagan skall ersättas med bilagan till denna förordning.
2. De nya artiklarna 3.1 och 5.2 b i förordning (EEG) nr 2299/89 skall inte tillämpas förrän sex månader efter den dag som anges i punkt 1. Kommissionen får bevilja ytterligare 12 månaders uppskov till de datoriserade bokningssystem som av objektiva skäl inte kan uppfylla bestämmelserna i artiklarna 3.1 och 5.2 b.
av den 14 december 1993
RÅDETS BESLUT av den 20 december 1994 om ingående av tilläggsprotokollet till interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Rumänien, å andra sidan, och till Europaavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan (94/48/EG)
med beaktande av Europeiska rådets slutsatser från mötet i Köpenhamn den 21 och 22 juni 1993,
Detta tilläggsprotokoll bör godkännas.
Tilläggsprotokollet till interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Rumänien, å andra sidan, och till Europaavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan, godkänns på Europeiska gemenskapens vägnar.
Rådets ordförande bemyndigas att utse den person som skall ha befogenhet att underteckna tilläggsprotokollet på Europeiska gemenskapens vägnar.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Enligt artikel 24 i beslut 90/424/EEG införs möjligheten att vidta en gemenskapsfinansierad åtgärd för att utrota och övervaka de sjukdomar som finns angivna i förteckningen i bilagan till detta beslut.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Följande strecksatser skall läggas till under Grupp 1 i förteckningen i bilagan till beslut 90/424/EEG:
- Anaplasmos, som överförs av smittbärande insekter i de franska utomeuropeiska departementen".
KOMMISSIONENS BESLUT av den 8 februari 1994 om ändring av rådets direktiv 89/556/EEG om djurhälsovillkor för handel inom gemenskapen med och import från tredje land av embryon från tamdjur av nötkreatur (Text av betydelse för EES) (94/113/EG)
med beaktande av rådets direktiv 89/556/EEG av den 25 september 1989 om djurhälsovillkor för handel inom gemenskapen med och import från tredje land av embryon från tamdjur av nötkreatur(1), senast ändrat genom direktiv 93/52/EEG(2), särskilt artikel 16 i detta, och med beaktande av följande:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
Det är i första hand medlemsstaterna som har ansvaret för riktade åtgärder för bekämpning av bedrägeribrott. Detta kräver ett nära samarbete mellan medlemsstaterna och kommissionen.
Kommissionen bör därför kunna rådfråga en kommitté bestående av företrädare för medlemsstaterna, vilken kan rådfrågas om alla frågor som rör förebyggande verksamhet, samarbete mellan medlemsstaterna och kommissionen, bekämpning av bedrägeribrott samt alla andra frågor med anknytning till det rättsliga skyddet för gemenskapens finansiella intressen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Kommittén skall ha en företrädare för kommissionen som ordförande.
3. De synpunkter som lagts fram av företrädarna för medlemsstaterna skall föras till protokollet.
med beaktande av Fördraget om Europeiska unionen, särskilt artiklarna J 3 och J 11 i detta,
med beaktande av artikel C i Fördraget om Europeiska unionen.
a) I syfte att verka för att en heltäckande fred i Mellanöstern sluts på grundval av FN:s säkerhetsråds resolutioner skall Europeiska unionen
- bidra till utformningen av de framtida förbindelserna mellan regionens parter i arbetsgruppen för vapenkontroll och regional säkerhet.
- bevara sin ledande roll i arbetsgruppen för regional ekonomisk utveckling (REDWG) och utveckla sitt deltagande i andra multinationella grupper,
- fortsätta att driva frågan om de förtroendeskapande åtgärder som den har förelagt parterna,
Artikel 2
- lämnande av stöd enligt befintliga riktlinjer till de andra parterna i de bilateral förhandlingarna, allteftersom dessa gör betydande framsteg mot fred.
a) Europeiska unionen lämna bistånd,
Artikel 4
Artikel 5
Europeiska unionen bekräftar att den är villig att fatta ytterligare praktiska beslut inom ramen för denna gemensamma åtgärd allteftersom fredsprocessen utvecklas.
Artikel 8
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Den behöriga myndigheten i medlemsstaterna får, med användning av icke-diskriminerande veterinära stickprovskontroller på bestämmelseorterna för djur och produkter, kontrollera att de krav som fastställs i artikel 3 i direktiv 90/425/EEG är uppfyllda. Myndigheten får samtidigt utföra provtagning i enlighet med artikel 5.1 a.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av följande: Rätten till rättsligt skydd för kretsmönster i halvledarprodukter i gemenskapen gäller för personer som har rätt till skydd i enlighet med artikel 3.1-3.5 i direktiv 87/54/EEG.
Detta skydd har tidigare, baserat på ömsesidighet, beviljats personer från vissa länder och territorier utanför gemenskapen, i vissa fall permanent, genom beslut 90/510/EEG(2), i andra interimistiskt, genom beslut 93/16/EEG(3).
Detta avtal och avtalet om inrättandet av Världshandelsorganisationen kommer att träda i kraft den 1 januari 1995 eller snarast möjligt efter den dagen. De industrialiserade länder som är parter i avtalet om inrättandet av Världshandelsorganisationen kommer att ha en frist av ett år efter det avtalets ikraftträdande för att genomföra bestämmelserna i avtalet om handelsrelaterade aspekter på immateriella rättigheter.
Artikel 1
b) Bolag eller andra juridiska personer från Canada som bedriver verklig och stadigvarande industriell eller affärsmässig verksamhet i Canada skall behandlas som om de bedrev verklig och stadigvarande industriell eller affärsmässig verksamhet inom en medlemsstats territorium.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av följande: En expertgrupp från kommissionen har gjort ett inspektionsbesök i Turkiet för att undersöka under vilka förhållanden levande tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar produceras och släpps ut på marknaden.
De behöriga turkiska myndigheterna har åtagit sig att regelbundet och snabbt till kommissionen överlämna uppgifter om förekomsten av plankton som innehåller toxiner i upptagningsområdena.
I enlighet med artikel 9.3 c i direktiv 91/492/EEG bör en förteckning upprättas över de anläggningar från vilka import av tvåskaliga blötdjur, tagghudingar, manteldjur och marina snäckor och sniglar är tillåten. Anläggningar får tas upp i förteckningen endast om de är officiellt godkända av de behöriga myndigheterna i Turkiet. Det åligger de behöriga turkiska myndigheterna att se till att bestämmelserna i artikel 9.3 c i direktiv 91/492/EEG följs.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
- Avsändande land: TURKIET.
- Förpackningsdatum med angivande av minst dag och månad.
2. Intygen skall innehålla namn, tjänsteställning och underskrift av den veterinär som representerar Ministry of Agriculture and Rural Affairs och dettas officiella stämpel i en annan färg än den som använts för övriga noteringar.
KOMMISSIONENS BESLUT av den 16 december 1994 om särskilda villkor för godkännandet av de förpackningsanläggningar som avses i rådets direktiv 77/99/EEG och om bestämmelser om saluhållandet av produkter därifrån (94/837/EG)
De hygienvillkor som skall gälla för sådan verksamhet bör fastställas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Förpackningsanläggningar som tar bort innerförpackningen och förser produkterna med ny innerförpackning skall uppfylla gällande villkor enligt bilaga A, kapitlen I och II till direktiv 77/99/EEG och de relevanta villkoren enligt bilaga B, kapitel I punkterna 1 a, 1 b, 1 d, 1 e och 1 f samt 2 a, 2 c, 2 i och 2 j till ovannämnda direktiv.
Produkter från de förpackningsanläggningar som avses i artikel 1.2 skall märkas med ett kontrollmärke i enlighet med de bestämmelser som fastställs i bilaga B, kapitel VI till direktiv 77/99/EEG. Den behöriga myndigheten skall tilldela förpackningsanläggningarna ett kontrollmärke.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av rådets direktiv 90/539/EEG av den 15 oktober 1990 om djurhälsoproblem för handeln inom gemenskapen med och import av fjäderfä och kläckningsägg från tredje land(2), ändrat genom del 1 kapitel 2 avsnitt A punkt 4. b och 4. c i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt artikel 9a, 9b och 10b i detta,
med beaktande av rådets direktiv 92/118/EEG av den 17 december 1992 om djurhälso- och hygienkrav för handel inom gemenskapen med produkter som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A. I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG, samt för import till gemenskapen av sådana produkter(5), ändrat genom del 1 kapitel 4 punkt 4. c i bilaga 1 V E till akten om anslutningsvillkoren för Norge, Österrike, Finland och Sverige och om anpassningarna i de fördrag som ligger till grund för Europeiska unionen, särskilt kapitel 2 första strecksatsen i bilaga 2 till denna, och med beaktande av följande:
Mot bakgrund av detta bör endast ett kommissionsbeslut antas om godkännande av det operativa programmet.
Artikel 1
Det finska programmets åtgärder avseende avelsfjäderfä och dagsgamla kycklingar som skall ingå i flockar av avelshöns eller flockar av produktionsfjäderfä godkänns.
Artikel 4
Det finska programmets åtgärder avseende nötkött och svinkött godkänns.
Artikel 7
Finland skall på dagen för ikraftträdandet av anslutningsfördraget sätta i kraft de lagar och andra författningar som är nödvändiga för att vidta de åtgärder som avses i artiklarna 1, 2, 3, 4, 5, 6 och 7.
Artikel 10
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(2), och
Förpliktelsen att uppfylla en procentsats på 5 % per sektor och per tullkontor gör det svårare att koncentrera personella resurser på export med hög risk.
Med tanke på nödvändigheten av att bestämmelserna om kontroll av exportbidrag tillämpas effektivt överallt i gemenskapen och mot bakgrund av de ekonomiska riskerna för gemenskapens tillgångar, måste regler antas på gemenskapsnivå.
Förordning (EEG) nr 386/90 ändras på följande sätt:
- per produktsektor.
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
Beträffande produkterna nr 3, 5, 6 och 7 i bifogade tabell har Tullkodexkommitténs sektion för tulltaxe- och statistiknomenklatur inte avgivit något yttrande inom den tid som dess ordförande bestämt.
Artikel 1
Om inte annat följer av de åtgärder som gäller i gemenskapen beträffande system med dubbelkontroll och med övervakning i för- och efterhand av import av textilprodukter till gemenskapen, får de bindande klassificeringsbesked som getts ut av medlemsstaternas tullmyndigheter rörande klassificeringen av varor i Kombinerade nomenklaturen och som inte överensstämmer med denna förordning, fortsatt åberopas av mottagaren enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en tid av 60 dagar.
KOMMISSIONENS FÖRORDNING (EG) nr 2701/94 av den 7 november 1994 om ändring av bilagorna 1, 2, 3 och 4 till rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung (Text av betydelse för EES)
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa maximalt tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), senast ändrad genom kommissionens förordning (EG) nr 1430/94(2), särskilt artikel 6-8 i denna, och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: Kommissionens förordning (EEG) nr 2273/93(2), ändrad genom förordning (EG) nr 2202/94(3), som gäller från och med den 1 januari 1995, skall ändras så att den överensstämmer med bestämmelserna i anslutningsakten.
Artikel 1
Denna förordning träder i kraft om och när Anslutningsfördraget för Norge, Österrike, Finland och Sverige träder i kraft.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
En grupp sakkunniga från kommissionen har företagit en resa till Marocko för att försäkra sig om villkoren för produktion, lagerhållning och sändning av fiskeriprodukter avsedda för gemenskapen.
De villkor som gäller det intyg som avses i artikel 11.4 a i direktiv 91/493/EEG omfattar fastställandet av en förlaga till ett intyg, valet av det eller de språk som intyget skall vara avfattat på samt firmatecknarens tjänsteställning.
DEMA har lämnat en officiell försäkran att de bestämmelser som anges i kapitel V i bilagan till direktiv 91/493/EEG och de krav som är likvärdiga med dem som fastställs i det direktivet för godkännande av anläggningar är uppfyllda.
1. Det intyg som avses i artikel 2.1 bör vara upprättat på minst ett av de officiella språken i den medlemsstat där kontrollen utförs.
Detta beslut tillämpas från och med den 1 mars 1995.
KOMMISSIONENS FÖRORDNING (EG) nr 1368/95 av den 16 juni 1995 om ändring av förordning (EEG) nr 2921/90 om beviljande av stöd för framställningen av kasein och kaseinater av skummjölk
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter (1), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94 (2), särskilt artikel 11.3 i denna, och
Förordning (EEG) nr 2921/90 ändras på följande sätt:
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Gränsvärden för högsta tillåtna restmängder bör endast fastställas sedan prövningar gjorts av Kommittén för veterinärmedicinska läkemedel av all relevant information om den berörda substansens restmängder vad beträffar säkerheten för konsumenten av livsmedel med animaliskt ursprung samt restmängdernas inverkan på industriell förädling av livsmedel:
Vad gäller veterinärmedicinska läkemedel avsedda för värpfåglar, mjölkdjur och honungsbin, måste gränsvärden för högsta tillåtna restmängder även för ägg, mjölk och honung fastställas.
För att möjliggöra komplettering av vetenskapliga studier danofloxacin och erytromycin bör bilaga III föras till förordning (EEG) nr 2377/90.
Denna förordning bör träda i kraft efter en period på 60 dagar, för att möjliggöra för medlemsländerna att föra de justeringar av tillstånden som kan komma att bli nödvändiga, samt för att få ut de berörda veterinärmedicinska läkemedlen på marknaden, vilket beviljats i överensstämmelse med rådets direktiv 81/851/EEG (3), senast ändrat genom direktiv 93/40/EEG (4), vilket tar hänsyn till denna förordnings bestämmelser.
Artikel 1
Denna förordning träder i kraft den sextionde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för humanläkemedel och yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
Inom ramen för de beslut som rör tillstånden för utsläppande på marknaden av läkemedel fastställs i denna förordning vissa närmare föreskrifter för hur Ständiga kommittén för humanläkemedel och Ständiga kommittén för veterinärmedicinska läkemedel (nedan kallade "kommittén") skall genomföra det förfarande som föreskrivs i artikel 73 i förordning (EEG) nr 2309/93, i artikel 37b i rådets direktiv 75/319/EEG (2) eller i artikel 42k i rådets direktiv 81/851/EEG (3).
Utom i undantagsfall, då det förslag till beslut som utarbetats av kommissionen inte är förenligt med yttrandet från Europeiska läkemedelsmyndigheten, skall ett skriftligt förfarande enligt bestämmelserna i artikel 3 tillämpas.
Om en medlemsstat inom tidsfristen på trettio dagar inkommer med en skriftlig begäran, vederbörligen motiverad, om att förslaget till beslut skall behandlas vid ett sammanträde med kommittén skall emellertid det skriftliga förfarandet avslutas, och ordföranden skall snarast möjligt sammankalla kommittén.
Ett nytt förfarande skall öppnas inom trettio dagar efter det att kommissionen har mottagit myndighetens svar.
Artikel 6
Artikel 7
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av kommissionens förslag,
Införandet av enhetliga visumhandlingar är ett viktigt steg mot harmoniseringen av viseringspolitiken. Artikel 7a i fördraget fastställer att den inre marknaden skall omfatta ett område utan inre gränser, där fri rörlighet för personer säkerställs i enlighet med bestämmelserna i fördraget. Åtgärden i fråga skall även ses som sammanhängande med de åtgärder som skall antas för tillämpningen av avdelning VI i Fördraget om Europeiska unionen.
För att undvika att uppgifterna i fråga sprids till flera personer än nödvändigt är det också viktigt att endast ett organ i varje medlemsstat utses för tryckningen av den enhetliga visumhandlingen, dock utan hinder av att kunna ersättas av ett annat organ om så behövs. Av säkerhetsskäl skall varje medlemsstat underrätta kommissionen och de övriga medlemsstaterna om det behöriga organets namn.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
1. De specifikationer som avses i artikel 2 är hemliga och skall inte offentliggöras. De meddelas enbart till de organ som utses av medlemsstaterna för tryckning och till personer som vederbörligen auktoriserats av en medlemsstat eller av kommissionen.
1. Utan att det påverkar tillämpningen av mer långtgående bestämmelser om skydd av uppgifter har de personer som beviljats ett visum rätt att kontrollera de personuppgifter som finns på visumhandlingen och i förekommande fall att få dessa rättade eller borttagna.
I denna förordning avses med "visumhandling" ett tillstånd eller beslut av en medlemsstat, som krävs för inresa på dess territorium för
Artikel 6
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över detta förslag inom den tidsfrist som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall anta sitt yttrande med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Vid omröstning inom kommittén skall medlemsstaternas företrädares röster vägas enligt samma artikel. Ordföranden skall inte delta i omröstningen.
Om rådet inte har fattat något beslut inom två månader, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas, såvida inte rådet med enkel majoritet har uttalat sig emot förslaget.
Artikel 8
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande (2),
Det har visat sig att bestämmelserna om märkning av jordbruksprodukter och livsmedel som innehåller en ingrediens med jordbruksursprung, producerad av odlare eller uppfödare som genomför omläggning av produktionen till ekologiskt jordbruk, som upphör att gälla den 1 juli 1995, bör förlängas för att denna produktion trots sina merkostnader, genom en lämplig märkning av produkterna, skall kunna göras lönande för producenterna.
Det har också framkommit att den upplysning som anges i bilaga V bör förbli frivillig men att den, för att förhindra missbruk, också bör begränsas till försäljning av färdigförpackade livsmedel eller till direktförsäljning från producent eller beredare till slutkonsumenter med villkor att produktens sammansättning kan identifieras.
Det har framkommit att vissa av de produkter som användes i enlighet med vedertagna regler för ekologisk odling inom gemenskapen, innan förordning (EEG) nr 2092/91 antogs, inte har inkluderats i bilaga II till nämnda förordning. Användningen av dessa produkter bör tillåtas i den utsträckning som den också är tillåten i det konventionella jordbruket.
1. I artikel 1.2 ersätts datumet "den 1 juli 1992" med datumet "den 30 juni 1995."
3. Artikel 4.3 ersätts med följande text:
"6. `ingredienser`: ämnen (inbegripet tillsatsämnen) som används vid beredningen av de produkter som avses i artikel 1.1 b såsom de definieras i artikel 6.4 i direktiv 78/112/EEG om tillnärmning av medlemsstaternas lagstiftning om märkning, presentation och reklam i fråga om livsmedel."
10. `ingrediensförteckning`: en sådan ingrediensförteckning som avses i artikel 6 i direktiv 79/112/EEG."
"d) för produkter som beretts efter den 1 januari 1997, skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som producenten är underställd. Valet av om namn eller kodnummer skall användas vid märkning åligger medlemsstaten som skall meddela sitt beslut till kommissionen."
"3. Vid märkning av och reklam för en produkt som åsyftas i artikel 1.1 b får beskrivningen av den saluförda varan endast innehålla uppgifter som hänvisar till ekologisk produktion om följande villkor är uppfyllda:
c) produkten innehåller enbart ämnen som finns förtecknade i bilaga VI punkt a i deras egenskap av ingredienser som inte är av jordbruksursprung,
f) produkten har beretts eller importerats av en leverantör som är underkastad den kontroll som anges i artiklarna 8 och 9,
10. Artikel 5.4 ersätts med följande text:
"5. Produkter som är föremål för märkning och reklam i enlighet med styckena 1 och 3 kan vara försedda med uppgifter som hänvisar till omställningen till ekologiskt jordbruk under förutsättning att:
c) uppgifterna inte vilseleder konsumenterna beträffande skillnader i förhållande till produkter som uppfyller alla krav i styckena 1 eller 3. Efter den 1 januari 1996 skall nämnda uppgifter bestå av orden `producerad under omställning till ekologiskt jordbruk` och presenteras i en färg, ett format och i en typstil som inte får vara mer framträdande än beskrivningen av den saluförda varan. Orden `ekologiskt jordbruk` får inte vara mer framträdande än orden `produkt under omställning till`,
12. Följande punkt skall införas efter artikel 5.5:
b) produktens alla andra ingredienser av jordbruksursprung omfattas av bilaga VI punkt C eller har godkänts provisoriskt av en medlemsstat i enlighet med vidtagna genomförandeåtgärder, i förekommande fall i enlighet med punkt 7,
e) produkten eller dess ingredienser av jordbruksursprung som anges i punkt a har inte behandlats med andra ämnen än de som finns i bilaga VI punkt B,
h) för produkter som beretts efter den 1 januari 1997, skall märkningen inkludera namn på och/eller kodnummer för den myndighet eller det kontrollorgan som den leverantör som utfört den sista beredningsåtgärden är underställd. Valet av om namn eller kodnummer skall användas åligger medlemsstaten som skall meddela sitt beslut till kommissionen."
a) minst 50 % av produktens ingredienser av jordbruksursprung uppfyller kraven i punkt 3 a,
- förekommer uteslutande i ingrediensförteckningen i enlighet med direktiv 79/112/EEG, senast ändrat genom direktiv 89/395/EEG,
e) uppgifterna i ingrediensförteckningen presenteras i samma färg, format och typstil."
15. Artikel 5.9 ersätts med följande text och punkterna 10 och 11 läggs till:
11. Kommissionen skall före den 1 juli 1999 göra en förnyad granskning av bestämmelserna i denna artikel och artikel 10 och presentera lämpliga förslag för deras eventuella ändring."
1. Ekologisk produktion innebär vid framställning av de produkter som anges i artikel 1.1 a med undantag för utsäde och vegetativt förökningsmaterial följande
c) endast utsäde och vegetativt förökningsmaterial som har producerats med den ekologiska produktionsmetod som anges i stycke 2 får användas.
b) förfarandet i artikel 14 kan användas för att fatta beslut om:
- införande av procedurregler och kriterier rörande det i a angivna undantaget och information om detta till berörda yrkesorganisationer, andra medlemsstater samt kommissionen.
"Artikel 6a
3. Trots vad som sägs i punkt 2, får plantor som inte erhållits i överensstämmelse med den ekologiska produktionsmetoden användas under en övergångsperiod fram till den 31 december 1997 förutsatt att följande villkor är uppfyllda:
c) plantorna härstammar från en producent som har accepterat ett kontrollsystem som är likvärdigt med det system som avses i artikel 9 och som har accepterat att tillämpa förbehållet i punkt b. Denna bestämmelse träder i kraft den 1 januari 1996,
f) utan att detta påverkar någon inskränkning som följer av det i punkt 4 angivna förfarandet skall alla godkännanden som lämnats i enlighet med denna punkt återkallas när bristsituationen avhjälpts och de skall löpa ut senast den 31 december 1997.
- benämning för berörd sort och art,
- övriga upplysningar som begärts av kommissionen eller medlemsstaterna.
18. I artikel 7 skall följande stycke läggas till efter punkt 1:
20. I artikel 9.5 b ersätts ordet "avvikelser" med orden "avvikelser och/eller överträdelser".
23. I artikel 9 införs följande punkt efter punkt 6:
"11. Utan att det påverkar tillämpningen av punkterna 5 och 6 skall de behöriga kontrollorganen från och med den 1 januari 1998 uppfylla kraven i EN 45011 av den 26 juni 1989."
a) överensstämmer med artikel 5.1 eller 5.3,
d) i märkningen är försedda med tillverkarens, beredarens eller säljarens namn på och/eller firma samt namn på eller kodnummer för kontrollmyndigheten eller kontrollorganet och övriga uppgifter som krävs i enlighet med reglerna för märkning av livsmedel som gäller i enlighet med gemenskapens lagstiftning."
"Allmänna åtgärder för verkställighet
2. Medlemsstaterna skall vidta nödvändiga åtgärder för att undvika bedräglig användning av de uppgifter som anges i artikel 2 och/eller bilaga V."
30. I artikel 11.6 a ersätts den sista meningen med följande text:
"7. Kommissionen får på begäran av en medlemsstat i enlighet med det i artikel 14 angivna förfarandet godkänna ett tredje lands kontrollorgan, som den berörda medlemsstaten på förhand har utvärderat, och föra upp den på den förteckning som anges i punkt 1 a. Kommissionen skall underrätta det tredje landet om detta."
33. I artikel 13 ersätts sista strecksatsen med följande strecksats:
Denna förordning träder i kraft den sjunde dagen efter dess offentliggörande i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapens officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Förordning (EEG) nr 2137/93 skall upphöra att gälla.
KOMMISSIONENS FÖRORDNING (EG) nr 2916/95 av den 18 december 1995 om ändring av vissa förordningar om den gemensamma organisationen av marknaderna för fjäderfäkött och ägg och om det gemensamma handelssystemet för äggalbumin och mjölkalbumin
med beaktande av rådets förordning (EEG) nr 234/79 av den 5 februari 1979 om förfarandet vid anpassning av Gemensamma tulltaxans nomenklatur för jordbruksprodukter (1), ändrad genom förordning (EEG) nr 3209/89 (2), särskilt artikel 2.1 i denna,
med beaktande av rådets förordning (EEG) nr 2783/75 av den 29 oktober 1975 om det gemensamma handelssystemet för äggalbumin och mjölkalbumin (6), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige och genom förordning (EG) nr 3290/94, särskilt artiklarna 2.2, 3.4 och 4.4 i denna,
med beaktande av rådets förordning (EG) nr 3492/93 av den 13 december 1993 om vissa förfaranden för tillämpningen av Europaavtalet om upprättandet av en associering mellan Europeiska gemenskaperna och deras medlemsstater å ena sidan och Polen, å den andra sidan (11), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EEG) nr 1601/92 av den 15 juni 1992 om särskilda åtgärder för Kanarieöarna rörande vissa jordbruksprodukter (14), senast ändrad genom kommissionens förordning (EG) nr 2537/95 (15), särskilt artikel 3.4 i denna,
med beaktande av rådets förordning (EG) nr 3642/93 av den 20 december 1993 om vissa förfaranden vid tillämpning av interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Rumänien, å andra sidan (19), senast ändrad genom förordning (EG) nr 3379/94, särskilt artikel 1 i denna,
med beaktande av rådets förordning (EG) nr 1277/95 av den 29 maj 1995 om vissa förfaranden för tillämpningen av avtalet om frihandel och vissa handelsrelaterade frågor mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Litauen, å andra sidan (22), särskilt artikel 1 i denna, och med beaktande av följande:
1. KN-nummer 0207 31 skall ersättas med KN-nummer 0207 34. KN-nummer 0207 39 90 och 0207 50 skall ersättas med numren 0207 13 91, 0207 14 91, 0207 26 91, 0207 27 91, 0207 35 91, 0207 36 81, 0207 36 85 och 0207 36 89. Nummer 1602 32 skall införas efter nummer 1602 31
2. KN-nummer 0105 12 skall införas före KN-nummer 0105 19
- i artiklarna 1 och 3.1 b i kommissionens förordning (EEG) nr 903/90 (26).
- kommissionens förordning (EG) nr 1431/94 (29),
- kommissionens förordning (EG) nr 1484/95 (32),
"Artikel 1 Om inte annat föreskrivs i denna förordning skall Gemensamma tulltaxans tullsatser tillämpas för följande produkter:
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av kommissionens förslag (1),
med beaktande av följande: Gemenskapen är allvarligt oroad över fartygsolyckor där människoliv går till spillo.
Människors säkerhet till sjöss kan förbättras avsevärt om ISM-koden tillämpas strikt och tvingande.
En strikt och tvingande tillämpning av ISM-koden är nödvändig för att säkerställa att säkerhetsorganisationssystem inrättas och bibehålls på vederbörligt sätt på både företags- och fartygsnivå av företag som bedriver havsgående trafik med ro-ro-passagerarfartyg.
Fartygssäkerheten är flaggstaternas huvudansvar, och medlemsstaterna kan säkerställa att adekvata bestämmelser om säkerhetsorganisation följs av de fartyg som för deras flagg och de företag som bedriver trafik med dessa. Det enda sättet att garantera säkerheten på alla ro-ro-passagerarfartyg, oberoende av flagg, som bedriver eller önskar bedriva reguljär trafik från medlemsstaternas hamnar är att medlemsstaterna, som villkor för att bedriva reguljär trafik från deras hamnar, kräver att säkerhetsbestämmelserna verkligen följs.
Medlemsstaterna kan komma att anse det nödvändigt att delegera eller att förlita sig på specialiserade organ för att uppfylla sina förpliktelser enligt denna förordning. Det lämpliga sättet att säkerställa en enhetlig och tillräcklig kontrollnivå är att kräva att dessa organ endast får vara sådana som uppfyller kraven i rådets direktiv 94/57/EG av den 22 november 1994 om gemensamma regler och standarder för organisationer som utför inspektioner och utövar tillsyn av fartyg och för sjöfartsadministrationernas verksamhet i förbindelse därmed (5).
Ett snabbt införande av dessa säkerhetsregler medför särskilda tekniska och administrativa problem för Grekland på grund av det mycket stora antal företag som är etablerade i Grekland och bedriver färjetrafik under grekisk flagg och uteslutande mellan grekiska hamnar. Ett undantag under begränsad tid för att hantera denna situation bör därför beviljas under beaktande även av att reguljär passagerar- och färjetrafik mellan grekiska hamnar fram till och med den 1 januari 2004 undantagits från tillämpningen av rådets förordning (EEG) nr 3577/92 av den 7 december 1992 om tillämpning av principen om frihet att tillhandahålla tjänster på sjötransportområdet inom medlemsstaterna (cabotage) (6).
Syftet med denna förordning är att öka säkerheten vid ledning och drift av ro-ro-passagerarfartyg samt att förhindra förorening som orsakas av sådana fartyg i reguljär trafik till eller från hamnar i medlemsstater inom Europeiska gemenskapen, genom att säkerställa att företag som bedriver trafik med ro-ro-passagerarfartyg följer bestämmelserna i ISM-koden genom
Artikel 2
b) reguljär trafik: en serie av resor med ett ro-ro-passagerarfartyg som upprätthåller trafik mellan två eller flera platser, antingen
c) företag: ro-ro-passagerarfartygets ägare eller någon annan organisation eller person, t.ex. redaren eller den som hyr fartyget utan besättning, som har övertagit fartygsägarens ansvar för ro-ro-passagerarfartygets drift.
f) administration: regeringen i den stat vars flagg ro-ro-passagerarfartyget har rätt att föra,
i) skyddade vatten: områden där sannolikheten per år för att det bildas vågor med en signifikant våghöjd över 1,5 m är mindre än 10 % och inom vilka ett ro-ro-passagerarfartyg aldrig befinner sig på större avstånd än 6 nautiska mil från en plats där fartyg kan söka skydd och där nödställda kan ta sig iland.
Artikel 4
Artikel 5
För tillämpningen av punkt 13.2 i ISM-koden får en medlemsstat endast utfärda dokument om godkänd säkerhetsorganisation för ett företag som har sin huvudsakliga verksamhetsort på dess eget territorium. Före ett sådant utfärdande skall medlemsstaterna samråda med administrationen i de stater vars flagg ifrågavarande företags ro-ro-passagerarfartyg har rätt att föra, om denna administration inte är den utfärdande medlemsstatens.
5. För tillämpningen av denna förordning och särskilt artikel 6 skall varje medlemsstat godkänna ett dokument om godkänd säkerhetsorganisation eller ett certifikat om godkänd säkerhetsorganisation som utfärdats av administrationen i någon annan medlemsstat eller av en erkänd organisation som handlar på dess vägnar.
Artikel 6
Om en medlemsstat anser att ett företag, trots att det har ett dokument om godkänd säkerhetsorganisation, inte kan bedriva reguljär trafik med ett ro-ro-passagerarfartyg till eller från dess hamnar på grund av risk för allvarlig fara för säkerheten för liv eller egendom eller för miljön får rätten att bedriva denna trafik dras in tills faran har undanröjts.
För att kunna beakta ISM-kodens allmänna begrepp skall kommissionen tre år efter denna förordnings ikraftträdande se över genomförandet av förordningen och föreslå lämpliga åtgärder.
a) Definitionen av ISM-koden i artikel 2.
Artikel 10
3. a) Kommissionen skall själv anta förslaget om det är förenligt med kommitténs yttrande.
Artikel 11
RÅDETS BESLUT av den 25 juni 1996 om förbättring av gemenskapens jordbruksstatistik (96/411/EG)
med beaktande av kommissionens förslag (1),
I ramprogrammet 1993 1997 som avses i beslut 93/464/EEG fastställs bland annat behovet av att bättre utnyttja de resurser som ägnas åt jordbruksstatistik genom genomförandet av resultaten av den "övervakningsverksamhet" som utfördes under det föregående statistiska programmet, som avses i rådets resolution av den 19 juni 1989 om genomförandet av en plan för prioriterade åtgärder för statistik: Europeiska gemenskapernas statistiska program (1989 1992) (4).
Anpassningar på det nationella planet måste samordnas på gemenskapsnivå för att säkerställa att
c) olika medlemsstaters metodologiska undersökningar om effektiva sätt att möta de nya informationsbehoven är lämpliga.
Denna samordning uppnås bäst genom att fastställa en formell struktur som gör det möjligt att gemensamt studera tekniska begränsningar och preferenser samt att fatta beslut som tar hänsyn både till gemenskapsintressen och nationella intressen.
Nödvändiga åtgärder bör vidtas för en eventuell förlängning av detta beslut inom ramen för nästa ramprogram för prioriterade åtgärder för statistik avseende åren efter 1997.
Artikel 1
Artikel 2
a) fastställa en gemensam plan för samordning av arbetet och en allmän ram för nödvändiga metodologiska beskrivningar,
Artikel 3
Artikel 4
2. Varje årlig teknisk handlingsplan skall innehålla en detaljerad verksamhetsplan för det kommande året och en preliminär tidsplan för de två följande åren. Vid utarbetandet av denna tidsplan skall hänsyn tas till följande:
c) Nödvändiga och tillgängliga resurser för alla planerade åtgärder.
Medlemsstaterna skall senast den 31 mars varje år (år n) överlämna
c) information om viktiga, större åtgärder som planeras för eller avses genomföras under de två följande åren (åren n + 2 och n + 3) och som är av betydelse för syftet med detta beslut.
Artikel 6
2. Kommissionen skall varje år i samband med den tekniska handlingsplanen och i enlighet med förfarandet i artikel 10 fastställa beloppet för gemenskapsbidraget till varje medlemsstat.
Flexibilitet
Anpassning till nya omständigheter
Ständiga kommittén för jordbruksstatistik
b) De åtgärder som medlemsstaterna föreslår för det kommande året och utsikterna för de följande två åren.
e) Eventuella ändringar i bilagorna I och II.
Kommissionen skall vidta de åtgärder som är nödvändiga för tillämpningen av detta beslut. Den skall biträdas av Ständiga kommittén för jordbruksstatistik, nedan kallad "kommittén".
Om de föreslagna åtgärderna inte är förenliga med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall besluta med kvalificerad majoritet.
Rapport
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
En anmälan om utsläppande på marknaden av en sådan produkt har inlämnats till den behöriga myndigheten i en medlemsstat (Nederländerna).
Efter att ha granskat de handlingar som inlämnats enligt direktiv 90/220/EEG och beaktat all den information som överlämnats av medlemsstaterna har kommissionen kommit fram till följande slutsatser:
- Det föreligger inga säkerhetsskäl för att på etiketten ange att produkten erhållits genom genetisk förändring.
Artiklarna 11.6 och 16.1 i direktivet ger ytterligare skydd om ny kunskap om risker förknippade med produkten blir tillgänglig.
Artikel 1
i) Barnase-genen från Bacillus amyloliquefaciens (ribonukleas) med promotorn PTA29 från Nicotiana tabaccum och terminatorn från nopalinsyntasgenen från Agrobacterium tumefaciens.
2. Medgivandet avser utsäde av alla hybrider mellan denna produkt och icke genetiskt modifierad cikoria.
- skall användas för odlingsverksamhet.
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Föreskrifterna i den mauretanska lagstiftningen i fråga om inspektion om hygienkontroll av fiskeriprodukter kan betraktas som likvärdiga med dem som fastställs genom direktiv 91/493/EEG.
Det är lämpligt att i enlighet med artikel 11.4 b i direktiv 91/493/EEG anbringa ett märke med uppgifter om det tredje landets namn och ursprungsanläggningens eller frysfartygets godkännandenummer på förpackningen för fiskeriprodukterna.
De åtgärder om föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
2. I intyget skall finnas namn och tjänstebeteckning på representanten för "Ministère des Pêches et de l'Économie Maritime - Centre National de Recherches Océanographiques et des Pêches - Département Valorisation et Inspection Sanitaire (MPEM - CNROP - DVIS)", dennes namnteckning samt den officiella stämpeln för MPEM - CNROP - DVIS; allt detta skall vara i en annan färg än övriga uppgifter i intyget.
KOMMISSIONENS BESLUT av den 14 oktober 1996 om särskilda importvillkor för fiskeri- och vattenbruksprodukter med ursprung i Elfenbenskusten (Text av betydelse för EES) (96/609/EG)
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktion och utsläppande på marknaden av fiskeriprodukter (1), senast ändrat genom direktiv 95/71/EG (2), särskilt artikel 11 i detta, och med beaktande av följande:
"Ministère de l'agriculture et des ressources animales - Direction générale des ressources animales (MARA-DGRA)" kan på ett effektivt sätt granska tillämpningen av den gällande lagstiftningen.
I enlighet med artikel 11.4 c i direktiv 91/493/EEG är det viktigt att fastställa en förteckning över godkända anläggningar. Denna förteckning bör fastställas på grundval av ett meddelande från Ministère de l'agriculture et des ressources animales - Direction générale des ressources animales (MARA-DGRA) till kommissionen. Det åligger alltså MARA-DGRA att försäkra sig om att de åtgärder som föreskrivs i detta syfte i artikel 11.4 i direktiv 91/493/EEG efterlevs.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 4
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande (2),
2. I rådets direktiv 88/299/EEG (6) fastställs villkor för undantag från förbudet att handla med vissa djurkategorier som anges i artikel 7 i direktiv 88/146/EEG, samt kött från dessa.
5. Resultaten från den undersökning som genomfördes av kommissionen 1990 till 1992 i medlemsstaterna visar på stor tillgång av â-agonister i animalieproduktionen vilket gynnar illegal användning.
8. Det är dessutom nödvändigt att garantera alla konsumenter samma villkor vid anskaffande av kött och livsmedel från kött, samt att erbjuda dem en produkt som motsvarar deras förväntningar. Med tanke på konsumenternas mottaglighet kan möjligheterna att få avsättning för produkterna i fråga härigenom enbart öka.
11. Levande djur som behandlas på detta sätt i terapeutiskt eller zootekniskt syfte och kött från dessa djur kan i princip inte bli föremål för handel med tanke på den inverkan det skulle ha på en effektiv kontroll av systemet. Undantag från detta förbud kan emellertid göras under vissa villkor beträffande handel inom gemenskapen och import från tredje land av djur avsedda för avel samt av uttjänta avelsdjur.
14. Direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG bör upphävas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Dessutom avses med
c) zooteknisk behandling:
d) illegal behandling: användning av icke godkända ämnen eller produkter eller användning av enligt gemenskapslagstiftningen godkända ämnen eller produkter för andra ändamål eller på andra villkor än vad som föreskrivs i gemenskapslagstiftningen eller - i förekommande fall - i de olika nationella lagstiftningarna.
a) Tillförsel av ämnen med tyreostatisk, östrogen, androgen eller gestagen verkan, samt â-agonister till ett husdjur eller vattenbruksdjur, oavsett på vilket sätt det sker.
d) Avyttring av kött från djur som avses i b.
Trots artikel 2 och 3, får medlemsstaterna tillåta följande:
- slag av godkända produkter,
Detta register skall på begäran ställas till behörig myndighets förfogande.
ii) â-agonister i form av injektion för att motverka livmoderkontraktioner hos kor i samband med kalvning.
Utan att det påverkar tillämpningen av första stycket i punkt 2 ii är emellertid terapeutisk behandling förbjuden för produktionsdjur, inklusive uttjänta avelsdjur.
Medlemsstaterna kan emellertid tillåta att synkronisering av östrus samt förberedelser av donatorer och recipienter för implantation av embryon inte utförs av veterinär utan endast på dennes ansvar.
Behandling i zootekniskt syfte är emellertid förbjuden på produktionsdjur, inklusive under gödningsperiod för uttjänta avelsdjur.
2. Följande kan emellertid inte tillåtas enligt punkt 1:
ii) Produkter där karenstiden är längre än 15 dygn efter behandling.
- med okända användningsvillkor,
Artikel 7
2. Kött eller produkter från djur som tillförts ämnen med östrogen, androgen eller gestagen verkan eller â-agonister kan enligt reglerna om undantag från detta direktiv avyttras för konsumtion endast om djuren i fråga har behandlats med veterinärmedicinska läkemedel som uppfyller kraven i artikel 6, och under förutsättning att den föreskrivna karenstiden har iakttagits innan djuren slaktas.
1) Att innehav av ämnen som avses i artikel 2 och artikel 3 a begränsas till personer som har tillstånd enligt nationell lagstiftning i enlighet med artikel 1 i direktiv 90/676/EEG (15), vid import, tillverkning, lagring, distribution, försäljning eller användning.
b) om djur behandlas illegalt,
3) Att sökande efter
a) visar på förekomst av ämnen eller produkter där användning eller innehav är förbjudet eller förekomsten av restsubstanser från ämnen vars tillförsel inneburit illegal behandling, skall dessa ämnen eller produkter beslagtas medan djur som eventuellt behandlats, eller deras kött, placeras under officiell kontroll till dess att nödvändiga påföljder genomförts,
Utan att det påverkar tillämpningen av direktiv 81/851/EEG skall företag som köper eller tillverkar ämnen med tyreostatisk, östrogen, androgen eller gestagen verkan eller â-agonister och de företag som har något slag av tillstånd för att utöva handel med nämnda substanser, samt de företag som köper eller producerar farmaceutiska produkter och veterinärmedicinska läkemedel utifrån dessa ämnen, upprätta ett register i kronologisk ordning över tillverkade eller införskaffade produkter och dem som överlåtits eller används för tillverkning av läkemedelspreparat och veterinärmedicinska läkemedel och till vem dessa har överlåtits eller sålts.
När resultaten av de kontroller som utförts i en medlemsstat visar att kraven i detta direktiv inte iakttagits i djurens eller produkternas ursprungsland, skall den behöriga myndigheten i den medlemsstaten tillämpa reglerna i rådets direktiv 89/608/EEG av den 21 november 1989 beträffande ömsesidigt stöd mellan medlemsstaternas administrativa myndigheter, samt samarbetet mellan dessa och kommissionen, i syfte att garantera att lagstiftningen på det veterinära och zootekniska området tillämpas korrekt (17).
2. Medlemsstaterna skall dessutom säkerställa att import från tredje land som förekommer på en av de listor som avses i punkt 1 förbjuds
ii) som tillförts de ämnen eller produkter som avses i artikel 3 a, utom om tillförseln sker enligt bestämmelser och krav i artikel 4, 5 och 7 i detta direktiv och om den karenstid som tillåts i de internationella rekommendationerna iakttagits,
4. Kontroller beträffande import från tredje land skall utföras enligt föreskrifterna i artikel 4.2 c i rådets direktiv 91/496/EEG av den 15 juli 1991 om fastställande av regler för hur veterinärkontroller skall organiseras för djur som importeras till gemenskapen från tredje land (18) och som enligt artikel 8.2 i rådets direktiv 90/675/EEG av den 10 december 1990 om principerna för organisering av veterinärkontroller av produkter som förs in i gemenskapen (19) från tredje land.
Artikel 13
Artikel 14
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
KOMMISSIONENS DIREKTIV 96/28/EG av den 10 maj 1996 om anpassning till teknisk utveckling av rådets direktiv 76/116/EEG om tillnärmning av medlemsstaternas lagstiftning om gödselmedel (Text av betydelse för EES)
med beaktande av rådets direktiv 76/116/EEG av den 18 december 1975 om tillnärmning av medlemsstaternas lagstiftning om gödselmedel (1), senast ändrat genom direktiv 89/530/EEG (2), särskilt artikel 9.1 i detta, och
För att nya gödselmedel skall kunna dra fördel av den "EEG-märkning" som avses i bilaga II i direktiv 76/116/EEG måste de läggas till bilaga I till det direktivet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Det gödselmedel som anges i bilaga I till detta direktiv skall läggas till del A punkt 1 "Kvävegödselmedel".
Artikel 3
Artikel 4
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande (1),
Erfarenheten visar att det har förekommit fall av bedräglig verksamhet på grund av den strukturella obalansen mellan de mervärdeskattesatser som medlemsstaterna tillämpar för jordbruksprodukter från blomster- och trädgårdsodling. Eftersom den strukturella obalansen direkt kan hänföras till tillämpningen av artikel 12.3 d bör detta ändras.
Artikel 1
2. Följande punkt skall införas i artikel 28.2:
Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
2. I sin resolution av den 15 januari 1985 om förbättring av energibesparingsprogrammen i medlemsstaterna (4) uppmanade rådet medlemsstaterna att fortsätta och i förekommande fall öka sina ansträngningar att främja en mer rationell användning av energi genom att utveckla en samordnad politik i fråga om energibesparingsåtgärder.
5. Det är nödvändigt att utgå från en hög skyddsnivå när det gäller förslagen om tillnärmning av bestämmelser i medlemsstaternas lagar och andra författningar rörande hälsa, säkerhet, miljöskydd och konsumentskydd. Detta direktiv garanterar en hög skyddsnivå för miljön och konsumenterna samtidigt som det syftar till en betydande förbättring av kylskåps och frysars energieffektivitet.
8. Rådets beslut 89/364/EEG av den 5 juni 1989 om ett åtgärdsprogram för gemenskapen för förbättrad effektivitet i elutnyttjandet (5) har den dubbla målsättningen att uppmuntra konsumenterna att välja apparater och utrustning som är mest energieffektiva samt att förbättra apparaternas och utrustningens energieffektivitet.
11. De åtgärder för en förbättrad energieffektivitet som genomförts på de senaste modellerna av kylskåp och frysar som finns på marknaden ökar inte påtagligt deras tillverkningskostnader och kan uppvägas inom några få år, eller till och med ännu snabbare, av de elektricitetsbesparingar de innebär. Denna beräkning tar inte hänsyn till den ytterligare fördel det innebär att externa kostnader i samband med elproduktionen försvinner, såsom exempelvis koldioxidutsläpp (CO2) och andra föroreningar.
14. Detta direktiv som syftar till att avlägsna tekniska hinder för en förbättrad energieffektivitet hos kylskåp och frysar för hushållsbruk skall följa den "nya metoden" som fastställs i rådets resolution av den 7 maj 1985 om en ny metod för teknisk harmonisering och standardisering (9) i vilken det uttryckligen bestäms att rättslig harmonisering begränsas till att genom direktiv anta de grundläggande krav vilka skall uppfyllas av varor som släpps ut på marknaden.
17. Med hänsyn till den internationella handeln bör internationell standard användas. Elförbrukningen för kylskåp och frysar definieras av Europeiska standardiseringsorganisationens standard EN 153 från juli 1995, på grundval av en internationell standard.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 3
3. a) Om kyl- och frysapparater omfattas av andra direktiv i vilka andra frågor behandlas och i vilka EG-märkning också föreskrivs innebär denna märkning att sådana kyl- och frysapparater skall förutsättas överensstämma även med bestämmelserna i dessa direktiv om det inte finns bevis om motsatsen.
De förfaranden som skall tillämpas för bedömning av överensstämmelse och de skyldigheter som rör EG-märkning av kyl- och frysapparater anges i bilaga II.
2. Det är förbjudet att på kyl- och frysapparaterna anbringa märkningar som skulle kunna vilseleda tredje man i fråga om EG-märkningens betydelse och grafiska utformning. Annan märkning får anbringas på apparaterna, emballaget, bruksanvisningen eller andra handlingar endast om EG-märkningen förblir synlig och läsbar.
2. Om överträdelsen fortgår skall medlemsstaten i enlighet med artikel 7 vidta alla nödvändiga åtgärder för att begränsa eller förbjuda att varan i fråga släpps ut på marknaden eller säkerställa att den tas ur försäljning.
2. Medlemsstaten skall utan dröjsmål underrätta kommissionen om och ange skälen för en sådan åtgärd. Kommissionen skall underrätta de övriga medlemsstaterna om detta.
Artikel 9
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 10
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100 a i detta,
Bestämmelserna i detta direktiv är förenliga med yttrandet från Kommittén för anpassning till tekniska framsteg, som upprättades i direktiv 74/150/EEG.
Bilaga I och II som är bilagor till rådets direktiv 76/432/EEG (3) ändras i enlighet med bilagan till detta direktiv.
- vägra att bevilja EG-typgodkännande eller ett sådant dokument som avses i artikel 10.1 sista strecksatsen i direktiv 74/150/EEG eller nationellt typgodkännande för en traktortyp, eller
- får vägra att bevilja nationellt typgodkännande
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 1 oktober 1997. De skall genast underrätta kommissionen om detta.
Artikel 4
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 100a i detta,
i enlighet med det i artikel 189b i fördraget angivna fördraget (3), och
De metoder som används vid officiella provningar i medlemsstaterna för att bestämma fibersammansättningen för textilvaror bör vara enhetliga både vad beträffar förbehandlingen av provet och den kvantitativa analysen.
I fråga om binära blandningar för vilka det inte finns någon enhetlig analysmetod på gemenskapsnivå, får det laboratorium som ansvarar för provningen bestämma sammansättningen av sådana blandningar. De får därvid använda någon vedertagen metod och ange resultatet i analysrapporten samt hur tillförlitlig den använda metoden är, i den mån detta är känt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Artikel 3
Det laboratorium som ansvarar för provningen av binära blandningar för vilka det inte finns någon enhetlig analysmetod på gemenskapsnivå skall bestämma sammansättningen av sådana blandningar genom att använda en vedertagen metod och ange resultatet i analysrapporten och hur tillförlitlig den använda metoden är, i den mån detta är känt.
2. Kommittén skall själv fastställa sin arbetsordning.
1. När det förfarande skall tillämpas som anges i denna artikel skall ärendet hänskjutas till kommittén av ordföranden, antingen på hans eget initiativ eller på begäran av en företrädare för en medlemsstat.
b) Om förslaget inte är förenligt med kommitténs yttrande, eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas.
Artikel 7
Direktiven som nämns i bilaga III del A upphävs utan att detta påverkar medlemsstaternas skyldigheter vad gäller de tidsfrister för överförande som anges i bilaga III del B.
Detta direktiv riktar sig till medlemsstaterna.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande (2), och
Olikheterna i nationell lagstiftning i fråga om sätten att kommersiellt bedriva transport på inre vattenvägar gynnar inte den inre marknadens funktion inom denna sektor, och därför bör på gemenskapsnivå gemensamma bestämmelser införas för hela marknaden för transport på inre vattenvägar, i enlighet med rådets resolution av den 24 oktober 1994 om strukturella förbättringar av transport på inre vattenvägar (4).
Med hänsyn till subsidiaritetsprincipen är det både nödvändigt och tillräckligt att på gemenskapsnivå fastställa en enhetlig tidsplan för successiv liberalisering av marknaden, samtidigt som ansvaret för genomförandet av liberaliseringen överlåts på medlemsstaterna.
Artikel 1
b) transportör: den som äger eller bedriver transport med ett eller flera fartyg på inre vattenvägar,
Artikel 2
Med undantag från artikel 2 får medlemsstaterna under en övergångsperiod fram till den 1 januari 2000 upprätthålla ett system med obligatoriska minimitaxor och system med befraktning i turordning under förutsättning
Artikel 4
b) Transporter som inte kan utföras effektivt av dessa system, bland annat
Artikel 5
- föreskriva att enstaka eller upprepade transporter, som erbjudits två gånger efter varandra inom systemet med befraktning i turordning utan att ha funnit någon användare, skall tas ur detta system och förhandlas fritt.
- Tidsavtal, inbegripet hyresavtal, enligt vilket transportören ställer ett eller flera fartyg med besättning till en kunds exklusiva förfogande för en fastställd tid för att transportera de varor den senare anförtror honom mot betalning av ett fastställt dagsbelopp. Avtalet skall ingås fritt mellan parterna.
Artikel 7
3. En medlemsstats begäran om att lämpliga åtgärder skall vidtas skall åtföljas av alla uppgifter som krävs för en bedömning av den ekonomiska situationen inom sektorn i fråga, bland annat
- prognoser om utvecklingen av efterfrågan.
Artikel 8
Yttrandet skall protokollföras, och dessutom har varje medlemsstat rätt att begära att få sin uppfattning tagen till protokollet.
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 1 januari 1997 och skall genast underrätta kommissionen om detta.
Artikel 10
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från sektionen för tulltaxe- och statistiknomenklatur inom tullkodexkommittén.
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas inom den gemensamma jordbrukspolitiken (3), senast ändrad genom förordning (EG) nr 150/95 (4), särskilt artikel 6.2 i denna, och
Vad gäller stöd till privat lagring av skummjölkspulver föreskrivs det i artikel 5 i förordning (EEG) nr 1362/87 att kontraktsparten vid export av skummjölkspulver genom undantag från gällande bestämmelser kan sälja ut lager när en kontraktsperiod på 30 dagar har löpt ut. Denna undantagsbestämmelse används sällan och försvårar i onödan förvaltning av ordningen. Den bör därför upphävas.
Artikel 1
"a) har framställts av en produktionsenhet som förbundit sig att löpande föra de register som avses i artikel 2.1 b i förordning (EG) nr 322/96,".
Artikel 2
"1. Anbudsgivare får delta i anbudsförfaranden endast
3. I artikel 7.1 andra stycket skall punkt c ersättas med följande:
"Artikel 9
- Om proteinhalten i den fettfria torrsubstansen är minst 35,6 % skall uppköpspriset vara det pris som anges i anbudet.
Proteinhalten fastställs enligt den metod som anges i bilaga I till förordning (EG) nr 322/96."
I bilagan till förordning (EEG) nr 1756/93 skall punkt 1 i avdelning C.I i del C och punkt 3 i del D ersättas med följande:
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 235 i detta,
KOMMISSIONENS FÖRORDNING (EG) nr 779/96 av den 29 april 1996 om tillämpningsföreskrifter till rådets förordning (EEG) nr 1785/81 i fråga om informationslämnande inom sockersektorn
med beaktande av rådets förordning (EEG) nr 1785/81 av den 30 juni 1981 om den gemensamma organisationen av marknaden för socker (1), senast ändrad genom förordning (EG) nr 1101/95 (2), särskilt artikel 39 i denna, och
För att noggrant kunna följa utvecklingen av handeln med tredje land behövs en nära och regelbunden övervakning med hänsyn till de intressekonflikter som kan uppkomma beroende på å ena sidan gemenskapens åtaganden inom ramen för ovan nämnda jordbruksavtal och åtgärder som kan behöva vidtas i samband med detta, särskilt i fråga om tillämpningen av artikel 23.4a i förordning (EEG) nr 1785/81, och å andra sidan gemenskapens åtaganden inom ramen för Internationella sockeravtalet. Det finns anledning för kommissionen att från början ha tillgång till relevant regelbunden information, inte bara vad gäller import och export av sådana produkter som omfattas av fastställda avgifter eller bidrag där licens utfärdas i enlighet med kommissionens förordning (EG) nr 1464/95 av den 27 juni 1995 om särskilda tillämpningsföreskrifter för systemet med import- och exportlicenser för socker (11), ändrad genom förordning (EG) nr 2136/95 (12), och när det gäller att iaktta de mera allmänna bestämmelserna i kommissionens förordning (EEG) nr 3719/88 (13), senast ändrad genom kommissionens förordningar (EG) nr 2137/95 (14) och (EEG) nr 3665/87 (15), senast ändrad genom förordning (EG) nr 1384/95 (16), utan även om import och export av sådana produkter som exporterats utan bidrag, med eller utan utfärdad licens, särskilt enligt bestämmelserna om aktiv förädling. Även importen av förmånssocker bör kunna följas för att ge möjlighet till effektiv tillämpning av bestämmelserna i kommissionens förordning (EEG) nr 2782/76 av den 17 november 1976 om fastställande av tillämpningsföreskrifter för import av förmånssocker (17), senast ändrad genom förordning (EEG) nr 1714/88 (18).
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för socker.
Vad gäller interventionsåtgärder som vidtagits i enlighet med artiklarna 9.1 och 11.1 i förordning (EEG) nr 1785/81 skall varje medlemsstat varje vecka, med avseende på närmast föregående vecka, till kommissionen anmäla
c) de kvantiteter vitsocker och råsocker, angivna i icke omräknad vikt, som sålts av interventionsorganet.
Artikel 3
2. På begäran av kommissionen, med avseende på en bestämd period, anmäla de kvantiteter vitsocker och råsocker som har denaturerats och ange vilken av de metoder som anges i bilagan till förordning (EEG) nr 100/72, som har använts.
1. Senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, anmäla de kvantiteter vitsocker, råsocker och sirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans för vilka:
2. Senast vid utgången av september månad varje år, med avseende på närmast föregående regleringsår, anmäla de kvantiteter vitsocker, råsocker och sirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans, fördelade på de produkter som räknas upp i bilagan till förordning (EEG) nr 1010/86, för vilka
3. Senast vid utgången av september månad varje år, med avseende på närmast föregående regleringsår, anmäla de kvantiteter basprodukter som avses i punkt 2 ovan vilka använts för framställning av sådana mellanprodukter som räknas upp i bilagan till förordning (EEG) nr 1729/78.
1. Varje vecka, med avseende på närmast föregående vecka:
- råsocker angivet i icke omräknad vikt KN-nr 1701 11 90 och 1701 12 90,
- inulinsirap uttryckt som torrsubstans, socker/isoglukos ekvivalent, KN-nr ex 1702 60 90,
d) med angivande av exportbidrag fastställda i enlighet med artikel 17.5 andra stycket a i förordning (EEG) nr 1785/81 de kvantiteter vitsocker, råsocker och sackarossirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans, för vilka exportlicens har utfärdats för att exportera i form av produkter enligt artikel 1.1 b i rådets förordning (EEG) nr 426/86 (29).
a) de kvantiteter - med angivande av exportbidrag för varje kvantitet - socker och sirap uttryckt som vitsocker, som avses i artikel 2 i förordning (EG) nr 1464/95, vilka exporterats i obearbetat skick utan exportlicens,
d) med angivande av exportbidrag fastställda i enlighet med artikel 17.5 andra stycket a i förordning (EEG) nr 1785/81 de kvantiteter vitsocker, råsocker och sackarossirap uttryckt som vitsocker, samt de kvantiteter isoglukos uttryckt som torrsubstans, som exporterats i form av produkter enligt bilaga I i rådets förordning (EEG) nr 804/68 (30), samt produkter enligt bilagan till kommissionens förordning (EG) nr 1222/94 (31),
Artikel 6
2. För varje kvartal, senast vid utgången av den tredje kalendermånaden efter det kvartal anmälan avser, de kvantiteter socker, uttryckt som vitsocker, som
Artikel 7
2. För varje kvartal, senast vid utgången av den andra kalendermånaden efter det kvartal anmälan avser, var för sig de kvantiteter socker som införts från tredje land och utförts i form av ersättningsprodukter inom ramen för förfarandet för aktiv förädling enligt definition i artikel 116 i förordning (EEG) nr 2913/92 (32).
1. Att senast vid utgången av varje kalendermånad, med avseende på närmast föregående kalendermånad, till kommissionen anmäla de kvantiteter socker, angivet i icke omräknad vikt, för vilka importlicenser har utfärdats i enlighet med förordning (EEG) nr 2782/76, med angivande av varje ursprungsland var för sig.
b) kopior av de dokument som avses i artikel 7.2 i förordning (EEG) nr 2782/76,
3. Att senast vid utgången av oktober månad varje år till kommissionen överlämna en förteckning över intyg och attester som utfärdats i enlighet med artiklarna 6 och 7 i förordning (EEG) nr 2782/76 och ange
c) den totala kvantiteten råsocker, angiven i ton i icke omräknad vikt, som är avsedd för direkt konsumtion,
Varje medlemsstat skall till kommissionen anmäla följande:
3. Före den 15 september varje år för vart och ett av de sockerproducerande, isoglukosproducerande och inulinsirapproducerande företagen på dess territorium, anmäla den slutliga produktionen under det närmast föregående regleringsåret av socker, isoglukos och inulinsirap, fastställd i enlighet med artikel 3.3 i förordning (EEG) nr 1443/82.
a) de kvantiteter socker, isoglukos och inulinsirap som avsatts på dess territorium för konsumtion,
Utan att det påverkar tillämpningen av artikel 2.1 andra stycket i förordningen (EEG) nr 2670/81 skall varje medlemsstat före den 15 mars varje år, med avseende på närmast föregående regleringsår, till kommissionen anmäla de kvantiteter C-socker, C-isoglukos och C-inulinsirap som enligt artikel 1.1 i förordning (EEG) nr 2670/81 anses vara avsatt på gemenskapens inre marknad.
1. Före den femtonde dagen varje månad, med avseende på den närmast föregående kalendermånaden, anmäla de totala kvantiteter B-socker och C-socker som i förekommande fall har förts över enligt artikel 27 i förordning (EEG) nr 1785/81.
- vad gäller produktionen av betsocker i Spanien skall datumet den 1 mars ersättas med den 15 april,
1. De godkännanden som avses i artikel 2.1 c och d i förordning (EEG) nr 1358/77 samt i förekommande fall godkännanden som har dragits tillbaka med stöd av artikel 1 i förordning (EEG) nr 1998/78.
b) de kvantiteter som har avsatts enligt artikel 12.1 i förordning (EEG) nr 1998/78.
1. Före den 1 september varje år, med avseende på närmast föregående regleringsår, och före den 1 januari varje år, med avseende på närmast föregående produktionsår, uppgifter rörande försörjningsbalanserna för socker, isoglukos och inulinsirap för ifrågavarande period enligt exemplet i bilaga II.
Varje medlemsstat skall för varje kalendermånad och senast vid utgången av den tredje påföljande kalendermånaden till kommissionen lämna de statistiska uppgifter som rör gemenskapens åtaganden inom ramen för Internationella sockeravtalet i enlighet med exemplen i bilagorna IV och V.
a) närmast föregående vecka: referensperioden från torsdag till onsdag,
Artikel 17
Artikel 18
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
I artikel 9 i förordning (EG) nr 2494/95 krävs att medlemsstaterna behandlar insamlade data/uppgifter så att HIKP kan tas fram som omfattar kategorierna COICOP (Classification of individual consumption by purpose) och där dessa kategorier behöver anpassas.
De åtgärder som denna förordning föreskriver överensstämmer med yttrandet från Statistiska programkommittén (SPC), inrättad genom rådets beslut 89/382/EEG, Euratom (2).
Artikel 1
Artikel 2
Artikel 3
Artikel 4
Artikel 5
Artikel 6
KOMMISSIONENS BESLUT av den 28 januari 1997 om fastställandet av ett identifieringssystem för förpackningsmaterial i enlighet med Europaparlamentets och rådets direktiv 94/62/EG om förpackningar och förpackningsavfall (Text av betydelse för EES) (97/129/EG)
med beaktande av Europaparlamentets och rådets direktiv 94/62/EG av den 20 december 1994 om förpackningar och förpackningsavfall (1), särskilt artikel 8.2 i detta, och
De åtgärder som avses i detta beslut är förenliga med yttrandet från den kommitté som inrättas genom artikel 21 i direktiv 94/62/EG.
Målet med detta beslut, vilket omfattar alla förpackningar enligt direktiv 94/62/EG, är att fastställa den numrering och de förkortningar som identifieringssystemet bygger på och ange vilket/vilka förpackningsmaterial som använts, samt specificera vilka material som bör omfattas av identifieringssystemet.
- De definitioner som anges i artikel 3 i direktiv 94/62/EG skall gälla om tillämpligt.
Numreringen och förkortningarna i identifieringssystemet skall vara de som anges i bilagorna.
Artikel 4
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av rådets direktiv 89/130/EEG, Euratom av den 13 februari 1989 om harmonisering av beräkningen av bruttonationalinkomst till marknadspris (1), och
Det är därför nödvändigt att uttolka reglerna för nuvarande upplaga av ENS i enlighet med dessa grundprinciper, så att det kan fastställas hur denna inkomst skall bokföras.
Artikel 1
Om det inte sker någon utdelning av inkomsten, skall denna behandlas som en inkomst utbetald av institutet för kollektiv investering till dess aktieägare, som dessa omedelbart återinvesterar i institutet för kollektiv investering. Detta innebär att inkomsten måste bokföras som kapital- och företagarinkomster på samma sätt som när det gäller utdelning av inkomst. Motsvarande summa kommer att bokföras på aktieägarnas finanskonto under posten aktier.
KOMMISSIONENS BESLUT av den 17 februari 1997 om förfarandet för bestyrkande av överensstämmelse av byggprodukter enligt artikel 20.2 i rådets direktiv 89/106/EEG beträffande konstruktionsvirke o.d. med tillbehör (Text av betydelse för EES) (97/176/EG)
med beaktande av rådets direktiv 89/106/EEG av den 21 december 1988 om tillnärmning av medlemsstaternas lagar och andra författningar om byggprodukter (1), ändrat genom direktiv 93/68/EEG (2), särskilt artikel 13.4 i detta, och med beaktande av följande:
De två förfarandena i artikel 13.3 beskrivs i detalj i bilaga III till direktiv 89/106/EEG. Det är därför nödvändigt att, i enlighet med bilaga III, klart specificera de metoder med vilka de två förfarandena skall genomföras för varje produkt eller produktgrupp, eftersom bilaga III anger att vissa system i första hand skall användas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Förfarandet för bestyrkande av överensstämmelse enligt bilaga III skall anges i uppdragen för harmoniserade standarder.
KOMMISSIONENS BESLUT av den 2 oktober 1997 om ändring av beslut 93/53/EEG om inrättande av en vetenskaplig kommitté för ursprungsbeteckningar, geografiska beteckningar och särartsskydd (Text av betydelse för EES) (97/656/EG)
med beaktande av följande: Det är lämpligt att närmare fastställa de villkor som skall gälla för medlemmarna i kommittén i deras tjänsteutövande.
Beslut 95/53/EEG ändras på följande sätt:
2. Artikel 6.2 skall ersättas med följande:
2. De får inte för yrkesmässiga syften använda de uppgifter som kommit till deras kännedom under och efter deras mandat som medlemmar i kommittén."
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
Kommissionens beslut 97/613/EG (2) av den 8 september 1997 om ett tillfälligt förbud mot import av pistaschmandlar och vissa produkter som är framställda från dessa, som har sitt ursprung i eller försänds från Iran gäller fram till den 15 december 1997 och bör upphävas.
Detta utgör en allvarlig fara för folkhälsan i gemenskapen och det är absolut nödvändigt att vidta skyddsåtgärder på gemenskapsnivå.
Pistaschmandlar och vissa produkter som är framställda av dessa skall ha producerats, sorterats, hanterats, bearbetats, förpackats och transporterats i överensstämmelse med god hygienisk sed. Det är nödvändigt att fastställa halten av aflatoxin B1 och den totala aflatoxinhalten i prover tagna från sändningen omedelbart innan den lämnar Iran.
Samråd har ägt rum med medlemsstaterna den 29 oktober 1997 och den 10 november 1997.
Detta beslut upphäver beslut 97/613/EG av den 8 september 1997 om ett tillfälligt förbud mot import av pistaschmandlar och vissa produkter som är framställda från dessa, som har sitt ursprung i eller försänds från Iran.
- pistaschmandlar som omfattas av KN-nummer 0802 50 00,
2. Pistaschmandlar och produkter som är framställda från dessa, och som har sitt ursprung i, eller sänds från Iran, skall endast införas i gemenskapen via en av de införselorter som anges i bilaga II.
5. De behöriga myndigheterna skall säkerställa att prover tas från varje sändning och att dessa analyseras för att fastställa halten av aflatoxin B1 och den totala aflatoxinhalten, och skall informera kommissionen om resultaten av dessa analyser.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Detta direktiv om benämningar på textilier föreskriver etiketter eller märkning eller angivelse av benämningarna på produktens textilfibrer för att säkerställa att konsumenternas intressen säkras genom rätt information.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1) Nummer 2 ändras på följande sätt:
2) Nummer 30 ändras på följande sätt:
4) Ett nytt nr 31 införs enligt följande:
- Texten i kolumnen "beteckning" skall vara "polyimid".
- En hänvisning till fotnoten har bifogats efter texten i kolumnen "beteckning". Fotnotens text skall vara följande:
Artikel 2
2) Ett nytt nr 31 införs enligt följande:
3) Ett nytt nr 32 införs enligt följande:
4) Ett nytt nr 33 införs enligt följande:
Artikel 3
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 57.2, 66 och 100a i detta,
i enlighet med det i artikel 189b i fördraget angivna förfarandet (3), och
3. De upphandlande myndigheter som omfattas av avtalet rättar sig efter direktiven 92/50/EEG, 93/36/EEG och 93/37/EEG, i dessas lydelse enligt det här direktivet, och tillämpar samma bestämmelser som gäller för tjänsteleverantörer, leverantörer och entreprenörer i tredje land som undertecknat avtalet, handlar i enlighet med avtalet.
6. När upphandlande myndigheter tilldelar ett kontrakt på sätt som avses med avtalet, måste möjligheterna att få tillgång till offentliga tjänste-, varu- samt bygg- och anläggningskontrakt som i enlighet med fördraget är tillgängliga för företag och produkter från medlemsstater, vara minst lika förmånliga som villkoren för tillgång till sådana offentliga upphandlingskontrakt inom Europeiska unionen som enligt bestämmelserna i avtalet tillämpas för företag och produkter med ursprung i tredje land som undertecknat avtalet.
9. Därför bör tillämpligheten av vissa av anpassningarna i direktiv 92/50/EEG utökas till att gälla alla tjänster som omfattas av detta direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"1. a) Det här direktivet gäller för
i) som tilldelas av de upphandlande myndigheter som anges i bilaga I till direktiv 93/36/EEG, förutsatt att det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 130 000 särskilda dragningsrätter (SDR) i ecu,
Den beräkningsmetod som avses i den här punkten skall på förslag av kommissionen ses över av Rådgivande kommittén för offentlig upphandling, i princip två år efter det att den tillämpats för första gången.
B) Punkt 8 utgår.
De upphandlande myndigheterna får emellertid besluta att viss information som rör tilldelningen av kontrakt och som nämns i första stycket inte skall lämnas ut om det bedöms att detta skulle hindra lagarnas tillämpning eller strida mot allmänintresset eller vara till skada för offentliga eller privata företags legitima kommersiella intressen eller för lojal konkurrens mellan tjänsteleverantörer.
"1. Denna artikel skall tillämpas på formgivningstävlingar som anordnas som led i ett förfarande för att tilldela ett kontrakt om tjänster med ett uppskattat värde, exklusive mervärdesskatt, på minst
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen ii för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i artikel 1 b, utom dem som nämns i bilaga I till direktiv 93/36/EEG.
- det tröskelvärde som avses i artikel 7.1 a andra strecksatsen i för de tjänster som avses i bilaga I A, utom tjänsterna i kategori 8 och telekommunikationstjänsterna i kategori 5, med CPC-referensnumren 7524, 7525 och 7526, som tilldelas av de upphandlande myndigheter som avses i bilaga I till direktiv 93/36/EEG, eller
"2. Tidsfristen för mottagande av anbud enligt punkt 1 får ersättas av en tidsfrist som är tillräckligt lång för att de berörda parterna skall ha möjlighet att lägga in giltiga anbud, och som i allmänhet inte understiger 36 dagar, men som aldrig är kortare än 22 dagar räknat från dagen för avsändande av meddelandet om upphandling, om de upphandlande myndigheterna har avsänt det preliminära förhandsmeddelande som avses i artikel 15.1, utformat enligt förlagan i bilaga III A (förhandsinformation), till Europeiska gemenskapernas officiella tidning minst 52 dagar och högst tolv månader före insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 15.2, och om det preliminära förhandsmeddelandet dessutom innehåller minst den information som föreskrivs i förlagan i bilaga III B (öppet förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
6. I artikel 23 blir den nu befintliga texten punkt 1 och följande punkt läggs till:
- att anbudets sekretess består i avvaktan på utvärderingen, och
7. Följande artikel förs in:
2. Den statistiska rapporten skall innehålla åtminstone följande:
- antal och värden för kontrakt som av varje upphandlande myndighet tilldelas över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, tjänstekategori i enlighet med den terminologi som anges i bilaga I och nationalitet för den tjänsteleverantör som tilldelas kontraktet samt, i fråga om förhandlade förfaranden, med uppdelning enligt artikel 11 under angivande av antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
d) Alla andra statistiska upplysningar som skall bestämmas i enlighet med förfarandet i artikel 40.3 och som begärs i enlighet med avtalet.
9. Bilaga III ersätts med den text som framgår av bilaga II till det här direktivet.
1. I artikel 5
i) de i artikel 1 b angivna upphandlande myndigheterna, inklusive kontrakt som tilldelas av de upphandlande myndigheterna inom försvarssektorn som anges i bilaga I i den mån det gäller varor som inte omfattas av bilaga II, om det uppskattade värdet, exklusive mervärdesskatt, uppgår till minst 200 000 särskilda dragningsrätter (SDR) i ecu,
c) Motvärdet i ecu och nationella valutor för de tröskelvärden som avses i a skall i princip revideras vartannat år med verkan från och med den 1 januari 1996. Beräkningen av detta motvärde skall grundas på det dagliga genomsnittsvärdet för dessa valutor uttryckt i ecu och för ecun uttryckt i SDR under de sista 24 månaderna fram till den sista augusti som föregår revisionen per den 1 januari.
B) läggs följande punkt till:
"1. De upphandlande myndigheterna skall inom 15 dagar efter det att en skriftlig begäran inkommit underrätta varje anbudssökande eller anbudsgivare vars ansökan eller anbud har förkastats om orsakerna till att hans ansökan eller anbud förkastats samt underrätta varje anbudsgivare som lämnat ett godtagbart anbud om utformningen av och de relativa fördelarna med det antagna anbudet samt namnet på den anbudsgivare som tilldelats kontraktet.
3. I artikel 10 skall följande punkt föras in:
"3 a. Tidsfristen för mottagande av anbud enligt punkt 3 får förkortas till 26 dagar, om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 9.1, utformat enligt förlagan i bilaga IV A (Förhandsinformation), till Europeiska gemenskapernas officiella tidning åtminstone 52 dagar och högst tolv månader före dagen för insändandet till Europeiska gemenskapernas officiella tidning av det meddelande om upphandling som avses i artikel 9.2, och om förhandsmeddelandet dessutom innehåller åtminstone den information som föreskrivs i förlagan i bilaga IV C (selektivt förfarande) eller, beroende på omständigheterna, i bilaga IV D (förhandlat förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
- att varje anbud innehåller de upplysningar som krävs för att utvärdera det,
- att öppnande av anbuden äger rum efter utgången av den tidsfrist som bestäms för avgivande av dessa."
3. Kommissionen skall på grundval av gjorda rättelser, ändringar eller tillägg uppdatera bilaga I i enlighet med det förfarande som anges i artikel 32.2 och skall se till att den offentliggörs i Europeiska gemenskapernas officiella tidning.
a) När det gäller de upphandlande myndigheter som avses i bilaga I
b) När det gäller övriga upphandlande myndigheter som omfattas av detta direktiv, antal och värden för kontrakt som tilldelas av varje kategori av upphandlande myndighet över tröskelvärdet, med uppdelning, så långt det är möjligt, efter förfarande, varukategori i enlighet med den terminologi som avses i artikel 9.1 och nationalitet för den varuleverantör som tilldelas kontraktet, fördelat enligt artikel 6 med uppgift om antal och värden för de kontrakt som tilldelas varje medlemsstat och tredje land.
3. Kommissionen skall enligt den förfarande som anges i artikel 32.2 bestämma arten av de statistiska upplysningar som krävs enligt det här direktivet."
Direktiv 93/37/EEG ändras på följande sätt:
"1. Det här direktivet gäller för
2. a) Motvärdet i ecu och nationella valutor för det tröskelvärde som fastställs i punkt 1 skall i princip revideras vartannat år med verkan från den 1 januari 1996. Beräkningen av detta motvärde skall grundas på den genomsnittliga dagskursen för ecun, uttryckt i SDR, och för dessa nationella valutor uttryckt i ecu under de sista 24 månaderna fram till den sista augusti som föregår revisionen per den 1 januari.
B) Följande punkt läggs till:
"1. De upphandlande myndigheterna skall inom 15 dagar efter det att en skriftlig begäran inkommit underrätta varje anbudssökande eller anbudsgivare vars ansökan eller anbud har förkastats om orsakerna till att hans ansökan eller anbud förkastats samt underrätta varje anbudsgivare som lämnat ett godtagbart anbud om utformningen av och de relativa fördelarna med det antagna anbudet samt namnet på den anbudsgivare som tilldelats kontraktet.
3. Artikel 12.2 ersätts med följande text:
"4. Tidsfristen för mottagande av anbud enligt punkt 3 får förkortas till 26 dagar, om de upphandlande myndigheterna har avsänt det förhandsmeddelande som avses i artikel 11.1, utformat enligt förlagan i bilaga IV A (Förhandsinformation), till Europeiska gemenskapernas officiella tidning minst 52 dagar och högst tolv månader före dagen för insändandet av det meddelande om upphandling som avses i artikel 11.2, och om förhandsmeddelandet dessutom innehåller minst den information som föreskrivs i förlagan i bilaga IV C (selektivt förfarande) eller, beroende på omständigheterna, i bilaga IV D (förhandlat förfarande), förutsatt att denna information fanns tillgänglig vid tidpunkten för meddelandets offentliggörande."
- att varje anbud innehåller de upplysningar som krävs för att utvärdera det,
- att öppnande av anbuden äger rum efter utgången av den tidsfrist som gäller för avgivande av dessa."
"1. För att möjliggöra bedömning av resultatet av tillämpningen av detta direktiv skall medlemsstaterna till kommissionen översända en statistisk rapport rörande de kontrakt för bygg- och anläggningsarbeten som under det föregående året tilldelats av de upphandlande myndigheterna senast den 31 oktober 1997 och därefter senast den 31 oktober varje år.
- det beräknade sammanlagda värdet för kontrakt som tilldelats av varje upphandlande myndighet under tröskelvärdet,
c) När det gäller de upphandlande myndigheter som anges i bilaga I till direktiv 93/36/EEG, antal och sammanlagt värde för kontrakt som tilldelats av varje upphandlande myndighet enligt undantagen från avtalet. När det gäller övriga upphandlande myndigheter som avses med detta direktiv, det sammanlagda värdet för kontrakt som tilldelats av varje kategori av upphandlande myndighet enligt undantagen från avtalet.
8. Bilaga IV ersätts med den text som framgår av bilaga IV till det här direktivet.
När en medlemsstat antar de bestämmelser som avses i första stycket skall de innehålla en hänvisning till det här direktivet eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Detta direktiv riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
I artikel 12 föreskrivs att tillverkare eller importörer av vissa ämnen som kan utgöra en allvarlig risk för människor eller miljön, kan åläggas att lämna de uppgifter som de har tillgång till.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Relevant information om exponering av människor eller miljön för ett ämne omfattar utsläpp av ämnet eller exponering av människor eller delar av miljön för ämnet under olika stadier av ämnets livscykel i enlighet med artikel 3.3 och bilaga 1 A till förordning (EG) nr 1488/94, där
- ett ämnes livscykel omfattar tillverkning, transport, lagring, blandning till en beredning eller annan bearbetning, användning och bortskaffade eller återvinning.
RÅDETS FÖRORDNING (EG) nr 552/97 av den 24 mars 1997 om tillfälligt upphävande av allmänna tullförmåner för Unionen Myanmar
med beaktande av rådets förordning (EG) nr 3281/94 av den 19 december 1994 om tillämpning av ett fyraårigt system med allmänna tullförmåner (1995-1998) för vissa industriprodukter med ursprung i utvecklingsländerna (1), särskilt artikel 12.3 i denna,
med beaktande av Europaparlamentets yttrande (4),
Enligt artikel 9 i förordning (EG) nr 3281/94 och artikel 9 i förordning (EG) nr 1256/96 kan förmånerna i fråga helt eller delvis tillfälligt upphävas under omständigheter som inbegriper utövande av någon form av tvångsarbete såsom det definieras i Genèvekonventionerna av den 25 september 1926 och den 7 september 1956 och i Internationella arbetsorganisationens (ILO) konventioner nr 29 och 105.
Kommissionen har i samråd med kommittén för förvaltningen av allmänna tullförmåner undersökt klagomålet av den 7 juni 1995 och de fakta som de klagande framlagt har bedömts vara tillräckliga för att inleda en undersökning. Kommissionen fattade beslut om detta i ett tillkännagivande av den 16 januari 1996 (6).
Kommissionen har, i syfte att komplettera de uppgifter som den har inhämtat i samband med undersökningen, uppmanat myndigheterna i Myanmar att samarbeta genom att tillåta en undersökningsdelegation inresa i landet. Myndigheterna i Myanmar har inte efterkommit denna uppmaning och eftersom villkoren i artikel 11.5 i förordning (EG) nr 3281/94 följaktligen är uppfyllda kan slutsatserna grundas på tillgängliga uppgifter.
En rapport om undersökningens slutsatser har överlämnats till kommittén för förvaltningen av allmänna tullförmåner enligt artikel 12.1 i förordning (EG) nr 3281/94.
Varor som redan avsänts till Europeiska gemenskapen bör undantas från detta upphävande av förmåner under förutsättning att de avsänts före den dag när denna förordning träder i kraft.
De allmänna tullförmåner enligt förordning (EG) nr 3281/94 och förordning (EG) nr 1256/96 är härmed tillfälligt upphävda för Unionen Myanmar.
Artikel 3
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I avdelning IV i förordning (EG) nr 2200/96 fastställs interventionsordningen för de produkter som avses i artikel 1.2 i denna. Tillämpningsföreskrifter till dessa bestämmelser bör därför fastställas.
För att tillämpa de begränsningar som föreskrivs i artiklarna 23 och 24 i förordning (EG) nr 2200/96 är det lämpligt att definiera den "saluförda kvantiteten" av en produkt som saluförs en producentorganisation med hänsyn till den faktiska produktion som producentorganisationen i fråga är upphov till, produktionen från andra producentorganisationer liksom produktionen från producenter som inte är anslutna till någon producentorganisation.
För att undvika oriktigheter vid tillämpningen av ordningen och garantera öppenhet och insyn bör producentorganisationerna i förväg meddela varje återtagande till kontrollmyndigheterna. Om ett sådant meddelande inte har lämnats får produkten avsättas först efter tillstånd från medlemsstaten. Dessutom måste ett kommunikationssystem inrättas, både för producentorganisationerna och för medlemsstaterna.
Bestämmelserna i kommissionens förordning (EEG) nr 3587/86 (3), senast ändrad genom förordning (EG) nr 1363/95 (4), (EEG) nr 827/90 (5), senast ändrad genom förordning (EG) nr 771/95 (6), (EEG) nr 2103/90 (7), ändrad genom förordning (EG) nr 1363/95, (EEG) nr 2276/92 (8), senast ändrad genom förordning (EG) nr 1363/95 och (EG) nr 113/97 (9), som har blivit föråldrade eller som skall ersättas av bestämmelserna i denna förordning, bör upphöra att gälla.
Artikel 1
1. Med produkter som "återtagits från marknaden" eller produkter som "inte saluförts" avses enligt denna förordning sådana produkter som inte sålts genom en producentorganisation, i enlighet med den interventionsordning som avses i förordning (EG) nr 2200/96.
1. För varje produkt skall den av en producentorganisation "saluförda kvantitet" som nämns i artikel 23.3 i förordning (EG) nr 2200/96 vara summan av
c) den produktion som framställts av medlemmar i andra producentorganisationer och som saluförts genom den berörda producentorganisationen i enlighet med artikel 11.1 c 3 andra och tredje strecksatsen i förordning (EG) nr 2200/96.
Artikel 4
Artikel 5
b) den produktion som medlemmarna i andra producentorganisationer salufört genom den berörda producentorganisationen i enlighet med artikel 11.1 c 3 andra och tredje strecksatsen i förordning (EG) nr 2200/96,
Artikel 6
1. De representativa marknader som avses i artikel 28.1 i förordning (EG) nr 2200/96 skall motsvaras av dem som anges i bilaga II till denna förordning.
1. Producentorganisationerna eller deras sammanslutningar skall minst 24 timmar i förväg underrätta de behöriga nationella myndigheterna om varje återtagande samt tillhandahålla en detaljerad förteckning över de produkter som avses för intervention, den kvantitet som beräknas för varje produkt.
b) Vid början av varje regleringsår uppgifterna om de uppodlade arealerna för varje produkt och eventuellt för varje sort.
2. Vid slutet av varje regleringsår skall medlemsstaterna för varje berörd produkt meddela kommissionen de uppgifter som anges i bilaga IV. Dessa uppgifter skall meddelas
3. Om medlemsstaterna inte lämnar in de uppgifter som avses i punkt 2 och om de meddelade uppgifterna med hänsyn till de objektiva fakta som kommissionen förfogar över verkar oriktiga, kan kommissionen i avvaktan på att ovan nämnda uppgifter läggs fram tillfälligt upphöra med den utbetalning av förskotten på de beräknade utgifter som avses i artikel 5.2 a i rådets förordning (EEG) nr 729/70 (10).
1. De produkter som återtagits från marknaden under ett visst regleringsår får ställas till förfogande för välgörenhetsorganisationer som godkänts av medlemsstaterna på deras begäran för gratis utdelning i enlighet med bestämmelserna i artikel 30.1 a första och tredje strecksatsen i förordning (EG) nr 2200/96.
b) föra särskilda räkenskaper över den aktuella verksamheten,
a) Välgörenhetsorganisationer som har tillstånd att genomföra utdelning på medlemsstatens territorium av produkter som har återtagits från marknaden.
De av medlemsstaterna utvalda institutioner som avses i artikel 30.1 a andra strecksatsen i förordning (EG) nr 2200/96 måste uppfylla villkoren i artikel 11.2 i denna förordning.
Vid slutet av varje regleringsår skall medlemsstaterna till kommissionen vidarebefordra de uppgifter om gratis utdelning som avses i bilaga VI.
2. För avsända produkter utgår inget exportbidrag. På tulldokumentet för export, transiteringshandlingen samt det kontrolldokument T 5 som eventuellt utfärdats skall uppgiften "utan bidrag" anges.
Om gratis utdelning sker utanför gemenskapen skall schablonbeloppen som avses i bilaga V täcka avståndet mellan platsen för återtagandet och den plats där sändningen lämnar gemenskapen.
- namnet på de mottagande organisationerna,
- vilka transportmedel som använts.
2. Enligt punkt 1 skall producentorganisationerna vid regleringsårets början ingå avtal med de välgörenhetsorganisationer som godkänts i enlighet med artikel 11.2 och 11.3 samt underrätta de behöriga nationella myndigheterna om dessa avtal så snart de ingåtts. Dessa myndigheter får fastställa en frist för slutandet av sådana avtal.
- den för varje produkt sannolika utdelningskvantiteten,
- den överenskomna överlåtelseplatsen,
5. Medlemsstaterna skall senast en månad efter det att avtalen slutits meddela kommissionen de uppgifter som avses i punkt 4.
- kvantiteten berörda produkter,
Artikel 17
De skall dessutom förvissa sig om att de produkter som inte saluförts överensstämmer med gällande normer, om sådana normer har fastställts med tillämpning av artikel 2.2 i förordning (EG) nr 2200/96.
Kontrollerna skall genomföras för varje producentorganisation minst en gång per regleringsår och den skall för varje produkt omfatta minst 10 % av betalningsansökningarna.
a) att verksamheten i fråga utförs på ett korrekt sätt,
2. Kontrollen enligt punkt 1 består av dokumentkontroller och fysiska kontroller, vilka skall avse berörda producentorganisationer och välgörenhetsorganisationer. Kontrollerna får bestå av stickprovskontroller som genomförs varje regleringsår och de skall avse minst 10 % av de utdelade kvantiteterna.
Artikel 19
b) de produkter som inte saluförts inte har avsatts i enlighet med artikel 30 i förordning (EG) nr 2200/96,
3. I händelse av uppsåtlig falskdeklaration eller av grov vårdslöshet skall den berörda producentorganisationen inte erhålla gemenskapskompensation för återtagande under det regleringsår för vilket oegentligheten konstaterats.
2. Godkännandet av den välgörenhetsorganisation som avses i artikel 11.2 dras in. Indragningen skall verkställas omedelbart, den skall gälla under minst ett regleringsår samt förlängas med hänsyn till hur allvarlig oegentligheten är.
Den avsändare som har fått transportkostnaderna täckta som avses i artikel 15 skall återbetala den dubbla summan av de belopp som erhållits för transportkostnader, ökad med en ränta beräknad på grundval av den tid som förflutit mellan utbetalningen och mottagarens återbetalning.
Artikel 21
Artikel 23
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Gemenskapens normer för frukt och grönsaker är utspridda på en rad gemenskapsbestämmelser. Det är nödvändigt att harmonisera vissa av dessa bestämmelser för att uppnå en enhetlig tillämpning av dessa normer och av kontrollen av deras överensstämmelse.
En kategori III har fastställts i de förordningar i vilka normer för purjolök, aubergine, zucchini, tomater, lök, endiver, körsbär, jordgubbar, brysselkål, bordsdruvor, trädgårdssallad, endivsallad, gurkor, citrusfrukter, äpplen och päron har fastställts. Denna kategori III tillämpades enbart i undantagsfall och har förlorat sin betydelse för färsk frukt och färska grönsaker. De internationella normerna innehåller ingen sådan kategori och för enkelhetens skull bör den tas bort i gemenskapens normer.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"Packare och/eller avsändare. Namn och adress eller officiellt utfärdat eller godkänt märke. Om en kod (ett märke) används skall "packare och/eller avsändare (eller motsvarande förkortning)" anges vid denna kod (detta märke)."
"Ursprungsland och eventuellt produktionsområde eller nationell, regional eller lokal benämning."
Artikel 2
KOMMISSIONENS FÖRORDNING (EG) nr 1054/97 av den 11 juni 1997 om klassificeringen av vissa varor i Kombinerade nomenklaturen
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 866/97 (2), särskilt artikel 9 i denna, och med beaktande av följande:
Med tillämpning av dessa allmänna regler måste de varor som beskrivs i första kolumnen i tabellen i bilagan till den här förordningen hänföras till de nummer i Kombinerade nomenklaturen som anges i andra kolumnen med stöd av den motivering som anges i tredje kolumnen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Nederländerna har begärt att kommissionen skall anpassa den årliga maximala fiskeansträngningsnivå som beviljats den nederländska flottan för vissa kvoter som de har tilldelats i enlighet med rådets förordning (EG) nr 390/97 av den 20 december 1996 om fastställande, för vissa fiskbestånd och grupper av fiskbestånd, av totala tillåtna fångstmängder under 1997 och av vissa villkor för fångsten (3), senast ändrad genom förordning (EG) nr 711/97 (4).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I kommissionens förordning (EG) nr 716/96 (3), senast ändrad genom förordning (EG) nr 2423/96 (4), föreskrivs undantagsåtgärder till stöd för nötköttsmarknaden i Förenade kungariket, särskilt genom att utbetalning till producenten av 0,9 ecu per kg levande vikt tillåts för djur som slaktas enligt den plan som föreskrivs i förordningen. Med hänsyn till prisutvecklingen i Förenade kungariket bör detta belopp justeras för kor samtidigt som en högsta tillåten vikt föreskrivs för djur som slaktas enligt planen. Denna högsta tillåtna vikt bör fastställas med hänsyn till den genomsnittliga vikten för kor. Följaktligen bör även gemenskapens bidrag, uttryckt i ecu per djur, justeras.
Artikel 1
- 0,9 ecu per kg levande vikt när det gäller alla andra djur.
- 2, när det gäller kor, och
Ett förskott på 80 % av det medfinansierade beloppet skall i enlighet med artikel 1.2 betalas ut efter det att de uppköpta djuren slaktats.
Om denna förbindelse inte görs skall det pris som skall betalas enligt punkt 1 för djuret i fråga nedsättas till ett belopp motsvarande det belopp som tillämpas för säsongsutjämningsbidraget. Om en premieansökan lämnas in för djuret i fråga, skall den berörda producenten tvingas betala tillbaka ett belopp motsvarande det belopp som tillämpas för säsongsutjämningsbidraget av det pris han erhållit för djuret i fråga. I båda dessa fall skall den andel medfinansiering från gemenskapen som avses i punkt 3 nedsättas med ett belopp motsvarande det belopp som skall tillämpas för säsongsutjämningsbidraget.
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 130 w i detta,
Verkningarna av en ekonomi som baseras på framställning av narkotika - eller som gör stora förtjänster på detta - på strukturen hos ett samhälle under utveckling, äventyrar en harmonisk integration av landet i världsekonomin.
Det är lämpligt att ge de utvecklingsländer som begär det ett institutionellt stöd för att de skall kunna bekämpa narkotikan mer effektivt.
Den fjärde AVS-EG-konventionen och de avtal om samarbete, association eller partnerskap som har ingåtts mellan gemenskapen och utvecklingsländerna innehåller klausuler om samarbete i kampen mot narkotikamissbruk och illegal handel med narkotika, kontroll av handeln med prekursorer, kemiska produkter och psykotropa ämnen samt utbyte av relevant information, inklusive åtgärder när det gäller penningtvätt. Det finns också ett samband mellan kampen mot narkotika och narkotikamissbruk och målen för samarbetet mellan gemenskapen och utvecklingsländerna.
En effektiv kamp mot narkotika måste också omfatta åtgärder mot penningtvätt som härrör från narkotikahandel, såsom antagandet av en lämplig rättslig ram och lämpliga mekanismer i berörda länder.
Ett finansiellt referensbelopp, i betydelsen enligt punkt 2 i förklaringen från Europaparlamentet, rådet och kommissionen av den 6 mars 1995 (3) har införts i den här förordningen för perioden 1998-2000 utan att detta påverkar den budgetansvariga myndighetens befogenheter enligt fördraget.
Inom ramen för sin politik för utvecklingssamarbete och med beaktande av de skadliga verkningarna på utvecklingsinsatserna som framställning, saluförande och konsumtion av narkotika har, skall gemenskapen genomföra samverkansåtgärder inom området narkotika och narkotikamissbruk i utvecklingsländerna, varvid företräde skall ges åt dem som har visat politisk vilja på högsta nivå att lösa sina problem med narkotika. Förekomsten av en sådan vilja kan manifesteras bl.a. genom ratificering av konventionen från 1961, ändrad genom protokollet från 1972, konventionen från 1971 och konventionen från 1988. Utvecklingsländernas engagemang skall ta sig uttryck bl.a. i genomförandet av inhemsk lagstiftning mot penningtvätt som härrör från illegal handel med narkotika.
Artikel 3
Samarbete inom gemenskapen skall ha formen av en dialog som återspeglar de genuina kulturskillnader som påverkar synen på problem som är knutna till narkotikan; detta är avgörande för att se till att strategierna för narkotikakontroll blir socialt och politiskt möjliga att genomföra.
- Utveckling av den institutionella kapaciteten, särskilt för att:
- Minska efterfrågan främst genom analys av fenomenet på lokal nivå, inrättandet av kontrollmekanismer riktade mot handeln med och konsumtionen av narkotika liksom av psykotropa ämnen, behandling och återanpassning av narkotikamissbrukare, och även att minska riskerna. Dessa aktioner bör integreras i den politik som förs på hälso- och utbildningsområdet, utveckling och kamp mot fattigdom och ekonomisk och social utslagning.
Särskild uppmärksamhet skall ägnas åt att få lokalbefolkningen och målgrupper att delta när aktionerna beslutas, planeras och genomförs.
Samarbetsparter som är berättigade till finansiellt stöd enligt denna förordning skall vara regionala och internationella organisationer, särskilt UNDCP, lokala och i medlemsstaterna förankrade icke-statliga organisationer, nationella, regionala och lokala styrande organ och myndigheter, organisationer förankrade i lokalsamhället, institut samt offentliga och privata aktörer.
2. Gemenskapens finansiering kan, beroende på behoven för varje åtgärd, täcka såväl investeringskostnader, med undantag av fastighetsköp, som driftskostnader i utländsk eller inhemsk valuta. Med undantag av utbildningsprogrammen skall dock driftskostnaderna normalt täckas endast under inledningsfasen, för att sedan gradvis minska.
5. Möjligheter till samfinansiering med andra bidragsgivare, i synnerhet medlemsstaterna, kan undersökas.
a) inrätta ett system för systematiskt utbyte och analys av information om finansierade åtgärder samt de åtgärder som gemenskapen och medlemsstaterna har för avsikt att finansiera,
Artikel 7
Det finansiella referensbeloppet för att genomföra detta program är 30 miljoner ecu för perioden 1998-2000.
1. Kommissionen skall ansvara för bedömning, godkännande och förvaltning av de åtgärder som omfattas av denna förordning enligt gällande budgetförfaranden och andra gällande förfaranden, särskilt de som föreskrivs i budgetförordningen för Europeiska gemenskapernas allmänna budget.
- Kulturella och sociala aspekter samt genus- och miljöaspekter.
3. Beslut om finansiering som överskrider 2 miljoner ecu för enskilda åtgärder enligt denna förordning samt alla förändringar som ger en ökning på mer än 20 % av den summa som ursprungligen godkänts för en sådan åtgärd, skall fattas enligt det förfarande som föreskrivs i artikel 10.
5. I alla överenskommelser eller kontrakt om finansiering som ingås enligt denna förordning, skall föreskrivas särskilt att kommissionen och revisionsrätten kan utföra kontroller på plats i enlighet med de sedvanliga villkor som kommissionen fastställer inom ramen för gällande bestämmelser, särskilt bestämmelserna i budgetförordningen för Europeiska gemenskapernas allmänna budget.
8. Leveranser skall härröra från medlemsstaterna, mottagarlandet eller andra utvecklingsländer. I vederbörligen styrkta undantagsfall kan leveranser härröra från andra länder.
- klart definierade och övervakade mål samt genomförandeindikatorer för samtliga projekt.
2. Kommissionens företrädare skall förelägga kommittén ett utkast till de åtgärder som skall vidtas. Kommittén skall yttra sig över utkastet inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Den skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Medlemsstaternas röster skall vägas enligt bestämmelserna i samma artikel. Ordföranden får inte rösta.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
1. Efter varje budgetår skall kommissionen överlämna en årsrapport till Europaparlamentet och rådet med en sammanfattning av de åtgärder som finansierats under budgetåret samt en utvärdering av hur denna förordning genomförts under denna period.
3. Kommissionen skall, senast en månad efter det att den fattat sitt beslut, informera medlemsstaterna om godkända åtgärder och projekt med uppgift om kostnad, art, mottagarland och parter.
KOMMISSIONENS BESLUT av den 25 februari 1998 om ett frågeformulär för medlemsstaternas rapporter om genomförande av rådets direktiv 94/67/EG om förbränning av farligt avfall (genomförande av rådets direktiv 91/692/EEG) (Text av betydelse för EES) (98/184/EG)
med beaktande av rådets direktiv 91/692/EEG av den 23 december 1991 om att standardisera och rationalisera rapporterna om genomförandet av vissa direktiv om miljön (1), särskilt artiklarna 5 och 6 i detta,
Rapporten skall utarbetas på grundval av frågeformulär eller mallar som kommissionen fastställer i enlighet med förfarandet i artikel 6 i direktiv 91/692/EG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
För detta ändamål bör beslut 94/411/EG ändras genom att dess bilaga II ersätts.
Artikel 1
Detta beslut riktar sig till medlemsstaterna.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113, tillsammans med artikel 228.2 första meningen och 228.3 första stycket, samt artikel 228.4 i detta,
Vissa genomförandeuppgifter har anförtrotts den gemensamma kommitté som inrättas genom avtalet, särskilt befogenheten att ändra vissa aspekter av de sektoriella bilagorna till detta.
Artikel 1
Artikel 2
1. Gemenskapen skall i den gemensamma kommitté som föreskrivs i artikel XI i avtalet och i de gemensamma sektoriella grupper som föreskrivs i artikel XII i avtalet och som inrättas genom de sektoriella bilagorna företrädas av kommissionen, som skall biträdas av den särskilda kommitté som utsetts av rådet. Kommissionen skall efter samråd med denna särskilda kommitté verkställa de utseenden, det informationsutbyte och de framställningar om kontroller som avses i artiklarna IX, X, XI.3 c och e, XII b och XIII i avtalet och i motsvarande bestämmelser i de sektoriella bilagorna.
RÅDETS DIREKTIV 98/29/EG av den 7 maj 1998 om harmonisering av huvudbestämmelserna för kreditförsäkringar för medellånga och långa exportaffärer
med beaktande av kommissionens förslag, och
(3) Skillnaderna mellan medlemsstaternas nu existerande statsstödda system för kreditförsäkringar för medellånga och långa exportaffärer med avseende på de huvudsakliga beståndsdelarna i försäkringsskyddet, premiebestämmelserna och täckningspolitiken kan leda till att konkurrensen mellan företag inom gemenskapen snedvrids.
(6) Regeringars (eller särskilda av regeringar kontrollerade institutioners) tillhandahållande av exportkreditgarantisystem eller exportkreditförsäkringssystem till premier som är otillräckliga för att täcka systemens långsiktiga kostnader och förluster betraktas som förbjudna exportsubventioner i det avtal om subventioner och utjämningsåtgärder som ingicks inom ramen för de multilaterala handelsförhandlingarna i Uruguayrundan (1986-1994) (1) (se artikel 3.1 a och bilaga I j till avtalet).
(9) Både harmonisering och samarbete är huvudsakliga och avgörande faktorer för gemenskapsexportens konkurrenskraft på marknader utanför gemenskapen.
(12) Den 15 maj 1991 gav den nämnda arbetsgruppen mandat till experter från var och en av de dåvarande medlemsstaterna vilka, under namnet Expertgruppen för den inre marknaden 1992, den 27 mars 1992, den 11 juni 1993 och den 9 februari 1994 lade fram rapporter, som innehöll ett antal förslag.
(15) Denna begynnande harmonisering av exportkreditförsäkringarna bör ses som ett steg i riktning mot samstämmighet mellan medlemsstaternas olika system.
Tillämpningsområde
Artikel 2
Artikel 3
Artikel 4
Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Den skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Kommittén skall fatta sitt beslut med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Medlemsstaternas röster skall vägas enligt bestämmelserna i samma artikel. Ordföranden får inte rösta.
- Får rådet fatta ett annat beslut med kvalificerad majoritet inom den tid som anges i första strecksatsen.
Kommissionen skall senast den 31 december 2001 förelägga rådet en rapport om de erfarenheter som gjorts och den samstämmighet som uppnåtts vid tillämpning av bestämmelserna i detta direktiv.
De förfaranden som föreskrivs i detta direktiv kompletterar dem som inrättas genom beslut 73/391/EEG (6).
Direktiv 70/509/EEG och direktiv 70/510/EEG upphävs.
Artikel 9
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande (2),
(2) Arbetstagarnas sociala skydd säkerställs genom lagstadgade system för social trygghet som supplerar kompletterande system för social trygghet.
(5) Ingen pension eller förmån bör omfattas både av bestämmelserna i detta direktiv och av förordningarna (EEG) nr 1408/71 och (EEG) nr 574/72 och därför kan ett kompletterande pensionssystem, som ligger inom dessa förordningars räckvidd därför att en medlemsstat har avgett en förklaring av denna innebörd enligt artikel 1 j i förordning (EEG) nr 1408/71, inte omfattas av bestämmelserna i detta direktiv.
(8) Den fria rörligheten för personer, som är en av de grundläggande rättigheterna i fördraget, är inte begränsad till anställda utan omfattar också egenföretagare.
(11) Medlemsstaterna bör vidta de åtgärder som behövs för att se till att förmåner enligt kompletterande pensionssystem betalas ut till försäkringstagare och före detta försäkringstagare samt till andra personer som är berättigade enligt sådana system i alla medlemsstater, eftersom alla restriktioner för betalningar och kapitalrörelser är förbjudna enligt artikel 73 b i fördraget.
(14) De arbetstagare som utövar sin rätt till fri rörlighet bör på ett adekvat sätt informeras av arbetsgivare, förvaltare eller andra som har ansvar för förvaltningen av de kompletterande pensionssystemen, särskilt vad gäller de val och de alternativ som erbjuds dem.
(17) I enlighet med subsidiaritets- och proportionalitetsprinciperna i artikel 3 b i fördraget kan målen för detta direktiv inte i tillräcklig utsträckning uppnås av medlemsstaterna utan de kan uppnås bättre på gemenskapsnivå. Detta direktiv går inte utöver vad som är nödvändigt för att uppnå dessa mål.
SYFTE OCH RÄCKVIDD
Artikel 2
DEFINITIONER
a) kompletterande pension: ålderspension och, om det föreskrivs i bestämmelserna för ett i enlighet med nationell lagstiftning och praxis inrättat kompletterande pensionssystem, invaliditets- och efterlevandeförmåner som är avsedda att komplettera eller ersätta de förmåner som de lagstadgade systemen för social trygghet föreskriver för samma försäkringsfall,
d) intjänade pensionsrättigheter: alla rättigheter till förmåner som erhålls efter uppfyllande av de krav som ställs enligt reglerna för ett kompletterande pensionssystem och, i förekommande fall, enligt nationell lagstiftning,
KAPITEL III
Likabehandling i fråga om bevarande av pensionsrättigheter
Gränsöverskridande betalningar
Avgifter till kompletterande pensionssystem från eller för utsända arbetstagare
Artikel 7
KAPITEL IV
Medlemsstaterna kan föreskriva att bestämmelserna i artikel 6 skall tillämpas endast på utsändningar som påbörjas 25 juli 2001.
Artikel 10
De skall underrätta kommissionen om vilka nationella myndigheter som skall kontaktas vad avser tillämpningen av detta direktiv.
Rapporten skall behandla direktivets tillämpning och skall vid behov innehålla förslag till ändringar som kan behöva göras.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande (2),
Produktionen av potatis och tomater intar en viktig plats inom gemenskapens jordbruk. Potatis- och tomatskörden hotas ständigt av skadegörare.
En av skadegörarna på potatis och tomat är Ralstonia solanacearum (Smith) Yabuuchi m.fl., den sjukdomsalstrande organism som orsakar mörk ringröta hos potatis och bakteriologisk vissnesjuka hos potatis och tomat. Sjukdomar som orsakats av denna sjukdomsalstrande organism har brutit ut i några delar av gemenskapen, och det existerar fortfarande några begränsade smittkällor.
Åtgärderna måste beakta att systematiska officiella undersökningar är nödvändiga för att lokalisera den sjukdomsalstrande organismen. Sådana undersökningar bör omfatta besiktningar och där så är lämpligt stickprovskontroller och test, eftersom sjukdomen under vissa miljömässiga omständigheter kan förbli latent och obemärkt både i potatisens förökningsmaterial och i lagrade potatisknölar. Spridningen av den sjukdomsalstrande organismen inom förökningsmaterialet är inte den viktigaste faktorn, men eftersom den sjukdomsalstrande organismen kan spridas med ytvatten och genom vissa besläktade vilda växter av familjen Solanaceae, utgör bevattning av potatis- och tomatgrödor med angripet vatten en smittorisk för sådana grödor. Den sjukdomsalstrande organismen kan också övervintra i självsådda (övervintrade) potatis- och tomatplantor, och dessa kan utgöra en smittkälla då de för över smittan från en odlingssäsong till nästa. Den sjukdomsalstrande organismen sprids också genom att potatisplantor angrips vid kontakt med smittad potatis och vid kontakt med utrustning för sättning, upptagning och hantering eller med transport- och lagringsbehållare som har angripits av skadegöraren vid tidigare kontakt med smittad potatis.
För att närmare kunna besluta om dessa allmänna åtgärder, liksom om de strängare eller ytterligare åtgärder som medlemsstaterna vidtar för att förhindra att den sjukdomsalstrande organismen förs in till deras territorium, är det önskvärt att medlemsstaterna samarbetar nära med kommissionen inom Ständiga kommittén för växtskydd (nedan kallad kommittén).
Detta direktiv rör de åtgärder som i medlemsstaterna skall vidtas mot Ralstonia solanacearum (Smith) Yabuuchi m.fl., tidigare känd som Pseudomonas solanacearum (Smith) Smith (nedan kallad skadegöraren) för att, såvitt avser skadegörarens värdväxter, vilka förtecknas i del 1 i bilaga I, (nedan kallade det förtecknade växtmaterialet),
c) om det konstateras förekomst av den, förhindra dess spridning och bekämpa den i syfte att utrota den.
2. De officiella undersökningar som anges i punkt 1 skall genomföras
c) när så är lämpligt på annat material i enlighet med lämpliga metoder.
4. Följande bestämmelse skall antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
- De lämpliga metoderna för de undersökningar som avses i punkt 2 första stycket under c.
Medlemsstaterna skall säkerställa att misstänkt förekomst eller bekräftad närvaro av skadegöraren på deras territorium rapporteras till deras egna ansvariga officiella organ.
2. I avvaktan på bekräftelse eller vederläggande av misstänkt förekomst enligt punkt 1, i varje enskilt fall av misstänkt förekomst där antingen
b) vidta åtgärder för att spåra den misstänkta förekomstens ursprung,
4. Följande bestämmelse får antas i enlighet med förfarandet i artikel 16a i direktiv 77/93/EEG:
1. Om ett officiellt eller officiellt övervakat laboratorietest som, med avseende på det förtecknade växtmaterialet, använder den lämpliga metod som anges i bilaga II, eller i andra fall, någon annan officiellt godkänd metod, bekräftar skadegörarens förekomst i ett stickprov som tagits på grund av detta direktiv, skall de ansvariga officiella organen i en medlemsstat, med beaktande av sunda vetenskapliga principer, skadegörarens biologiska egenskaper och de särskilda systemen för produktion, marknadsföring och bearbetning av skadegörarens värdväxt i den medlemsstaten,
ii) Förklara följande angripet: Det förtecknade växtmaterialet, sändningen och/eller partiet som stickprovet togs från, maskinerna, fordonet, fartyget, lagret, eller delar av dessa, och alla andra föremål, inklusive förpackningsmaterialet som har varit i kontakt med det förtecknade växtmaterial från vilket stickprovet togs. I förekommande fall även förklara följande som angripet: Det eller de fält, den eller de enheter för skyddad växtproduktion och den eller de produktionsplatser där det förtecknade växtmaterialet har skördats och från vilka stickprovet tagits. I fråga om de stickprov som tagits under växtsäsongen förklara följande för angripet: Det eller de fält, den eller de produktionsplatser, och i förekommande fall den eller de enheter för skyddad växtproduktion som stickprovet togs ifrån.
b) I fråga om grödor från värdväxter som inte nämns under a, då det har konstaterats att det finns en risk vid produktionen av det förtecknade växtmaterialet vidta följande åtgärder:
iii) Fastställa det troliga angreppet och avgränsa ett område i enlighet med punkterna a iii respektive a iv i förhållande till produktionen av det förtecknade växtmaterialet.
ii) Förklara det ytvatten som provet eller proven har tagits från för angripet i den utsträckning som det är lämpligt och på grundval av undersökningen enligt punkt i.
Medlemsstaterna skall samtidigt till kommissionen överlämna en tilläggsanmälan enligt 3 a i bilaga V. Innehållet i denna anmälan enligt detta stycke skall omedelbart överlämnas till kommitténs ledamöter.
1. Medlemsstaterna skall föreskriva att det förtecknade växtmaterial som förklarats för angripet enligt artikel 5.1 a ii inte får planteras och att det, under övervakning av och med godkännande av deras ansvariga officiella organ, skall underkastas någon av bestämmelserna i punkt 1 i bilaga VI, så att det kan fastställas att det inte finns någon identifierbar risk för att skadegöraren sprids.
4. Utan att det påverkar tillämpningen av de åtgärder som genomförs enligt punkterna 1 3 skall medlemsstaterna föreskriva att ett antal åtgärder skall genomföras enligt punkterna 4.1 och 4.2 i bilaga VI inom det område som avgränsas enligt artikel 5.1 a iv och 5.1 c iii. Uppgifter om dessa åtgärder skall varje år anmälas till de andra medlemsstaterna och till kommissionen. Innehållet i denna anmälan för överlämnas till kommittén.
De ovannämnda testerna skall utföras av en medlemsstat
ii) genom tester av allt ursprungligt klonurval av utsädespotatis eller tidigare generationer inklusive det ursprungliga klonurvalet i de fall då inget släktskap genom klon har påvisats och
- Tillämpningsföreskrifterna i punkt 1, andra stycket, punkt a.
Medlemsstaterna skall förbjuda innehav och hantering av skadegöraren.
Artikel 10
Artikel 12
2. Medlemsstaterna skall omedelbart till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv. Kommissionen skall underrätta de övriga medlemsstaterna om detta.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europaparlamentets yttrande (2),
(2) Råolja och petroleumprodukter som importeras spelar fortfarande en viktig roll i gemenskapens energiförsörjning. Varje svårighet, även om den är tillfällig, som leder till att leveranserna av dessa produkter begränsas, eller till att deras pris stiger avsevärt på de internationella marknaderna skulle kunna orsaka allvarliga störningar i gemenskapens ekonomiska verksamhet. Gemenskapen måste därför vara i stånd att upphäva eller åtminstone minska de skadeverkningar som skulle kunna uppstå i sådana fall. Det är nödvändigt att uppdatera direktiv 68/414/EEG så att det anpassas till den verklighet som råder på gemenskapens inre marknad och till utvecklingen på oljemarknaderna.
(5) Lagerhållningen av olja måste vara så organiserad att den inte förhindrar att den inre marknaden fungerar väl.
(8) Lagren måste stå till medlemsstaternas förfogande om det uppstår svårigheter med oljeförsörjningen. Medlemsstaterna bör ha befogenhet och möjlighet att kontrollera användningen av lagren så att de utan dröjsmål kan göras tillgängliga för de områden där behovet av oljeleveranser är störst.
(11) I syfte att organisera lagerhållningen får medlemsstaterna använda sig av ett system med ett lagerhållande organ eller en enhet som skall förvalta alla eller en del av de lager som utgör lagerhållningsskyldigheten. Eventuell överskjutande del bör hållas av raffinaderier och andra marknadsaktörer. Partnerskap mellan staten och branschen är nödvändigt för att lagerhållningssystemen skall fungera effektivt och säkert.
(14) Det finns ett behov av att anpassa och förenkla gemenskapens system för statistisk rapportering av oljelager.
(17) Det är lämpligt att bygga ut den administrativa tillsynen av lagren och att inrätta verkningsfulla system för kontroll och verifiering av lagren. Införandet av ett sådant kontrollsystem kräver ett sanktionssystem.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Medlemsstaterna skall anta de lagar och andra författningar som är lämpliga för att, om inte annat följer av bestämmelserna i artikel 7, inom gemenskapen, alltid hålla sina lager av petroleumprodukter på en nivå som för varje typ av petroleumprodukter, enligt förteckningen i artikel 2, motsvarar minst 90 dagars genomsnittlig, daglig inhemsk förbrukning under det föregående kalenderåret enligt artikel 4.
3. För att kunna uppfylla kraven i punkterna 1 och 2 får medlemsstaterna besluta att använda sig av ett lagerhållande organ eller en enhet med ansvar för att hålla alla lagren eller en del av dessa.
En medlemsstats lagerhållningsskyldighet skall baseras på det föregående kalenderårets inhemska förbrukning. Vid början av varje kalenderår skall medlemsstaterna göra en ny beräkning av sin lagerhållningsskyldighet senast den 31 mars varje år och säkerställa att de uppfyller sina nya skyldigheter så snart som möjligt och i vart fall senast den 31 juli varje år.
Obligatoriska lager enligt artikel 1 får hållas i form av råolja, halvfabrikat och färdiga produkter.
- på grundval av raffinaderiernas produktionsprogram i den berörda staten under innevarande år, eller
a) Punkt 1 skall ersättas med följande:
I dessa fall skall den medlemsstat på vars territorium lagren hålls inom ramen för ett sådant avtal inte hindra att dessa lager överförs till de andra medlemsstaterna, för vars räkning lagren hålls enligt avtalet. Den skall kontrollera dessa lager i enlighet med förfarandena som närmare anges i det avtalet men inte räkna in dem i sitt statistiska sammandrag. Den medlemsstat för vars räkning lagren hålls får räkna in dem i sitt statistiska sammandrag.
Avtalen skall uppfylla följande villkor:
- De skall närmare ange de förfaranden som skall användas för att kontrollera och identifiera de lager som föreskrivs, bland annat metoder för att utföra inspektioner och för samarbetet under dessa.
När lager, upprättade enligt sådana avtal, inte ägs av det företag, det organ/enhet som har skyldighet att hålla lager, utan hålls tillgängliga för företaget, organet/enheten av ett annat företag, organ/enhet, skall följande villkor uppfyllas:
- Uppgifter om var lagren är belägna och/eller om de företag som håller lagren tillgängliga för det företag, organ/enhet som har rätt till dem, liksom lagrade kvantiteter och produktkategorier eller uppgift om att det rör sig om lagrad råolja, skall anges.
"Följaktligen skall särskilt följande uteslutas från det statistiska sammandraget: inhemsk råolja som ännu inte utvunnits, mängder som skall användas till bunkring för havsgående fartyg, mängder i direkt transitering, frånsett de i punkt 2 angivna lagren, mängder i rörledningar, tankbilar och tankvagnar på järnväg, i lagertankar på detaljistmarknaden samt hos små förbrukare. De mängder som innehas av de väpnade styrkorna och de som innehas av oljebolag för deras räkning skall också uteslutas från det statistiska sammandraget." 8. Följande artikel skall införas:
9. Följande artikel skall införas:
Artikel 2
1. Medlemsstaterna skall före den 1 januari 2000 sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
På grund av Hellenska republikens särskilda situation garanteras den en ej förnybar extra period på tre år för att tillämpa detta direktivs skyldigheter vad gäller att låta mängder som används till bunkring av internationellt flyg ingå när det gäller att beräkna inhemsk förbrukning.
Artikel 6
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Gränsvärden bör fastställas först efter det att Kommittén för veterinärmedicinska läkemedel har granskat all relevant information beträffande säkerheten med restmängder av ämnet i fråga för den som konsumerar livsmedel med animaliskt ursprung samt restmängdernas påverkan på den industriella bearbetningen av livsmedel.
För veterinärmedicinska läkemedel som är avsedda för äggläggande fåglar, mjölkdjur eller honungsbin, måste gränsvärden även fastställas för ägg, mjölk eller honung.
För att möjliggöra komplettering av vetenskapliga studier, bör giltighetstiden för temporära MRL, tidigare definierad i bilaga III i förordning (EEG) nr 2377/90, förlängas för penetamat.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av följande: I förordning (EG) nr 3051/95 föreskrivs att företag och medlemsstater skall följa bestämmelserna i Internationella säkerhetsorganisationskoden, som antogs av Internationella sjöfartsorganisationen (IMO) genom församlingens resolution A.741 (18) av den 4 november 1993, för ro-ro-fartyg i trafik till eller från hamnar i medlemsstater inom gemenskapen.
Det är lämpligt att säkerställa att giltigheten för vissa dokument och certifikat som redan utfärdats inte påverkas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Det åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för humle.
Bilagan till denna förordning skall ersätta bilagan till förordning (EEG) nr 3077/78.
KOMMISSIONENS FÖRORDNING (EG) nr 726/98 av den 31 mars 1998 om ändring av förordning (EG) nr 2543/95 om tillämpningsföreskrifter för ordningen med exportlicenser inom olivoljesektorn
med beaktande av rådets förordning nr 136/66/EEG av den 22 september 1966 om den gemensamma organisationen av marknaden för oljor och fetter (1), senast ändrad genom förordning (EG) nr 1581/96 (2), särskilt artiklarna 2 och 3 i denna, och
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för oljor och fetter.
Förordning (EG) nr 2543/95 ändras på följande sätt:
1. Punkt 3 skall ersättas med följande:
b) 1 ecu per 100 kg netto i övriga fall."
3. Artikel 3 skall ändras på följande sätt:
2. Första stycket i punkt 2 skall ersättas med följande:
"Dessa åtgärder skall gälla exportlicenser med förutfastställelse av bidraget, och får variera mellan produktkoderna i nomenklaturen över exportbidrag för jordbruksprodukter."
5. Följande stycke skall läggas till:
1. I punkt 1 första stycket skall "torsdag" ersättas med "fredag".
3. I punkt 1 b skall "måndagen innan" ändras till "från och med föregående period fredag till och med torsdag, med separat angivelse för licenser med förutfastställelse av bidraget i förhållande till licenser utan förutfastställelse av bidraget".
5. I punkt 2 tredje strecksatsen skall "i förekommande fall" läggas till framför "tillämplig".
7. I punkt 3 skall följande läggas till:
Artikel 2
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av följande: I kommissionens förordning (EEG) nr 1722/93 av den 30 juni 1993 om tillämpningsföreskrifter för rådet förordningar (EEG) nr 1766/92 och (EEG) nr 1418/76 om produktionsbidrag inom spannmåls- respektive rissektorn (5), senast ändrad genom kommissionens förordning (EG) nr 1516/95 (6), föreskrivs att det vid beräkning av produktionsbidrag skall göras åtskillnad mellan stärkelse av majs, vete, potatis och ris, å ena sidan, och stärkelse av korn och havre, å andra sidan. I praktiken har visat sig att det inte längre är nödvändigt att fastställa ett särskilt belopp för stärkelse av korn och havre, och att det enhetliga bidragsbeloppet hädanefter kan tillämpas på all stärkelse utan risk för att otillbörlig kompensation ges.
I förordningen förskrivs för närvarande att medlemsstaterna varje månad till kommissionen skall överlämna de statistiska uppgifter som både omfattar de kvantiteter stärkelse som har fått produktionsbidrag och de produkter i vilka stärkelse har använts. Det har blivit uppenbart att detta informationslämnande sker onödigt ofta och att det vore lämpligt att ersätta det med kvartalsvisa meddelanden.
"Artikel 3
i) marknadspriset på majs i gemenskapen, giltigt i fem dagar före den dag det fastställs, med hänsyn tagen till priserna för vete, och
3. Det bidrag som skall utbetalas skall beräknas i enlighet med punkt 2 och multipliceras med koefficienten i bilaga II, vilken motsvarar KN-numret för den stärkelse som faktiskt används för att framställa de godkända produkterna.
"3. Bidragslicensen skall innefatta de upplysningar som anges i artikel 5.2, och dessutom bidragssatsen och den sista dag då licensen är giltig, som skall vara den sista dagen i den femte månaden efter den månad då licensen utfärdades.
Om någon av de kvantiteter stärkelse som anges i licensen bearbetas under det regleringsår för spannmål som följer på det år då ansökan inkom, skall dock det bidrag som skall utbetalas för den stärkelse som bearbetas under det nya regleringsåret justeras med skillnaden mellan det interventionspris som tillämpas under den månad då bidragslicensen utfärdas och det som tillämpas under bearbetningsmånaden, multiplicerad med koefficienten 1,60. Den omräkningskurs som skall användas för att uttrycka bidragsbeloppet i nationell valuta skall vara den som gäller den dag då stärkelsen bearbetas."
4) I artikel 10.4 skall följande stycke läggas till:
Inom tre månader från utgången av varje kvartal skall medlemsstaterna underrätta kommissionen om typen, kvantiteterna och ursprunget (majs, vete, potatis, korn, havre eller ris) av den stärkelse för vilken bidrag har utbetalats och om typen och kvantiteterna av de produkter till vilka stärkelsen har använts."
KOMMISSIONENS FÖRORDNING (EG) nr 1549/98 av den 17 juli 1998 om komplettering av bilagan till förordning (EG) nr 1107/96 beträffande registrering av geografiska beteckningar och ursprungsbeteckningar enligt förfarandet i artikel 17 i rådets förordning (EEG) nr 2081/92 (Text av betydelse för EES)
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska beteckningar och ursprungsbeteckningar för jordbruksprodukter och livsmedel (1), senast ändrad genom kommissionens förordning (EG) nr 1068/97 (2), särskilt artikel 17.2 i denna, och av följande skäl:
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för geografiska och ursprungsbeteckningar.
Bilagan till förordning (EG) nr 1107/96 skall kompletteras med beteckningarna i bilagan till denna förordning.
KOMMISSIONENS FÖRORDNING (EG) nr 1900/98 av den 4 september 1998 om ändring av bilaga I till rådets förordning (EEG) nr 2092/91 om ekologisk produktion av jordbruksprodukter och uppgifter därom på jordbruksprodukter och livsmedel
med beaktande av rådets förordning (EEG) nr 2092/91 av den 24 juni 1991 om ekologisk produktion av jordbruksprodukter och uppgifter därom på jordbruksprodukter och livsmedel (1), senast ändrad genom kommissionens förordning (EG) nr 1488/97 (2), särskilt artikel 13 första och andra strecksatsen i denna, och
Vissa komponenter, särskilt halm och gödsel, kan dock för tillfället inte erhållas i tillräckligt stora mängder från ekologisk produktion. Därför bör en lämplig övergångsperiod fastställas så att producenterna kan anpassa sig till de nya kraven.
Övergångsperiodens varaktighet kan komma att ses över om situationen på något sätt förändras när det gäller tillgången på halm och gödsel från ekologisk odling.
Artikel 1
1. Denna förordning träder i kraft den 1 december 1998.
- produkter som anges i punkt 5.2 i bilagan och som inte kommer från jordbruksföretag där en ekologisk produktionsmetod används, men som vid behov uppfyller de krav som anges i del A i bilaga II till förordning (EEG) nr 2092/91,
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
med beaktande av Fördraget om upprättandet av ett gemensamt råd och en gemensam kommission för Europeiska gemenskaperna,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
De regler för avrundning av penningbelopp som fastställs i rådets förordning (EG) nr 1103/97 av den 17 juni 1997 om vissa bestämmelser som har samband med införandet av euron (3) skall tillämpas.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EEG) nr 1898/87 av den 2 juli 1987 om skydd av beteckningar som används vid saluhållande av mjölk och mjölkprodukter (2), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 4.2 i denna, och
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandena från berörda förvaltningskommittéer.
"b) Den genomsnittliga fetthalten får inte avvika med mer än en procentenhet från den angivna halten. Fetthalten i de enskilda proven får avvika med endast två procentenheter från den angivna halten.
Artikel 2
med beaktande av protokoll nr 3 om stadgan för Europeiska centralbankssystemet och Europeiska centralbanken (nedan kallad stadgan), särskilt artikel 19.2 i denna,
med beaktande av kommissionens yttrande (3)
(2) Enligt artikel 19.2 i stadgan skall rådet bland annat fastställa basen för minimireserverna och den högsta tillåtna kvoten mellan dessa reserver och basen för dem.
(5) För att systemet med åläggande av minimireserver skall kunna vara ett effektivt verktyg för förvaltning av penningmarknaden och monetär styrning måste det ha en sådan struktur att ECB har förmåga och flexibilitet nog att tillämpa krav på reserver mot bakgrund av och med hänsyn tagen till förändringar i fråga om de ekonomiska och finansiella förhållandena i de deltagande medlemsstaterna. I detta avseende måste ECB vara flexibel nog att reagera för ny betalningsteknik, såsom utvecklingen av elektroniska pengar. För att begränsa möjligheterna att kringgå kraven på minimireserver får ECB tillämpa dem på skyldigheter som härrör från poster utanför balansräkningen, särskilt poster som - antingen enskilt eller i kombination med andra poster i eller utanför balansräkningen - är jämförbara med skyldigheter som är upptagna i balansräkningen.
(8) ECBS och ECB har anförtrotts uppgiften att förbereda de penningpolitiska instrumenten så att de kan ha trätt i kraft fullt ut när den tredje etappen av den ekonomiska och monetära unionen inleds (nedan kallad tredje etappen). Ett väsentligt inslag i dessa förberedelser är att innan den tredje etappen inleds ha antagit de ECB-förordningar enligt vilka instituten måste hålla minimireserver från och med den 1 januari 1999. Det är önskvärt att under 1998 underrätta marknadsaktörerna om de detaljerade bestämmelser som ECB kan anse sig behöva anta för att genomföra systemet med minimireserver. Det är därför nödvändigt att från och med dagen för den här förordningens ikraftträdande utrusta ECB med föreskrivande befogenheter.
2) nationell centralbank: en deltagande medlemsstats centralbank,
5) sanktioner: böter, viten, straffränta och räntelös insättning.
ECB kan på icke-diskriminerande grunder undanta institut från kraven på minimireserver enligt kriterier som fastställs av ECB.
1. I basen för de minimireserver som ECB enligt artikel 19.1 i stadgan kan ålägga institut att hålla skall, om inte annat följer av bestämmelserna i punkterna 2 och 3, ingå
iii) skyldigheter som ett institut helt eller delvis har gentemot andra institut enligt villkor som fastställs av ECB, och inte heller
3. ECB kan på icke-diskriminerande grunder tillåta att vissa typer av tillgångar undantas från kategorier av skyldigheter som ingår i basen för minimireserverna.
1. Reservkvoterna, som ECB får fastställa enligt artikel 19.1 i stadgan, får inte överstiga 10 % av någon relevant skyldighet som utgör en del av basen för minimireserverna, men kan vara 0 %.
Föreskrivande befogenheter
Rätt att inhämta och verifiera uppgifterna
3. Rätten att verifiera uppgifter skall inbegripa rätten att
c) ta kopior av eller göra utdrag ur sådana räkenskaper och register, och
4. ECB får delegera verkställandet av de rättigheter som avses i punkterna 1-3 till de nationella centralbankerna. I enlighet med första strecksatsen i artikel 34.1 i stadgan skall ECB ha befogenhet att i en förordning ytterligare precisera villkoren för utövande av kontrollrätten.
1. Om ett institut underlåter att hålla alla eller delar av de minimireserver som krävs enligt den här förordningen och de ECB-förordningar eller ECB-beslut som är knutna till denna förordning, får ECB förelägga institutet endera av följande sanktioner:
2. När en sanktion föreläggs enligt punkt 1 skall principerna och förfarandena i förordning (EG) nr 2532/98 tillämpas. Artikel 2.1 och 2.3 och artikel 3.1-3.4 i den förordningen skall dock inte vara tillämpliga, och de tidsfrister som avses i artikel 3.6-3.8 skall förkortas till femton dagar.
Slutbestämmelser
av den 16 december 1998
VERKSTÄLLANDE KOMMITTÉN HAR FATTAT DETTA BESLUT
Det ligger i alla Schengenstaters intresse att inom ramen för sin gemensamma politik avseende rörligheten för personer fastställa enhetliga regler för utfärdande av viseringar för att undvika eventuella negativa följder när det gäller inresor till territoriet och den inre säkerheten.
Detta formulär medger en stor flexibilitet när det gäller användningen och skall anpassas till den rättsliga situationen för varje avtalsslutande part eftersom Schengenstaterna för närvarande använder mycket olika formulär för olika typer av åtaganden.
- Utseendet och strukturen.
1. Följande punkt skall läggas till i kapitel V punkt 1.4 i de gemensamma konsulära anvisningarna: "I de fall då det enligt Schengenstaternas nationella lagstiftning föreligger krav på inbjudningar av privatpersoner eller affärsmän, åtagandeförklaringar eller bevis för att bostad finns skall dessa dokument framläggas i form av ett enhetligt formulär(1)."
4. De modelldokument som utarbetats av de avtalsslutande parterna skall bifogas de gemensamma konsulära anvisningarna som bilaga 15.
7. Dokumentet skall utarbetas på minst tre språk.
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
Kommissionen skall välja det av de två förfaranden, enligt artikel 13.3 i direktiv 89/106/EEG för bestyrkande av överensstämmelse av en produkt, som är "minst betungande och samtidigt förenligt med kraven på säkerhet". Detta innebär att det är nödvändigt att besluta om huruvida en tillverkningskontroll i fabriken under tillverkarens ansvar är ett nödvändigt och tillräckligt villkor för bestyrkande av överensstämmelse för en bestämd produkt eller produktgrupp, eller om det av orsaker som rör uppfyllandet av de kriterier som avses i artikel 13.4 krävs att ett godkänt certifieringsorgan deltar.
Det förfarande som avses i artikel 13.3 a motsvarar de system som anges i det första alternativet utan fortlöpande övervakning, samt i det andra och det tredje alternativet i punkt 2 ii i bilaga III och det förfarande som avses i artikel 13.3 b motsvarar de system som anges i punkt 2 i i bilaga III, samt i det första alternativet med fortlöpande övervakning i punkt 2 ii i bilaga III.
Artikel 1
För de produkter som anges i bilaga II skall överensstämmelsen bestyrkas genom ett förfarande där, förutom ett system för tillverkningskontroll i fabriken som genomförs av tillverkaren, även ett godkänt certifieringsorgan tar del i bedömningen och övervakningen av tillverkningskontrollen eller av själva produkten.
Artikel 4
av den 28 juni 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
2. Direktiv 91/682/EEG skall upphöra att gälla från och med den 1 juli 1999 och ersättas med direktiv 98/56/EG.
5. Detta system innehåller också uppgifter om upprätthållande av sorter och om skillnader i förhållande till de mest liknande sorterna.
8. De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga kommittén för förökningsmaterial av prydnadsväxter.
I detta direktiv fastställs ytterligare genomförandebestämmelser för de listor över sorter av prydnadsväxter och förökningsmaterial av prydnadsväxter som förs av leverantörer i enlighet med artikel 9.1 fjärde strecksatsen i direktiv 98/56/EG.
i) Sortens namn, i tillämpliga fall tillsammans med dess allmänt kända synonymer.
iv) Om möjligt, uppgifter om hur sorten skiljer sig från de sorter som mest liknar den.
Direktiv 93/78/EEG skall upphöra att gälla från och med det datum som avses i artikel 4 i detta direktiv.
2. När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Medlemsstaterna skall besluta om hur en sådan hänvisning skall göras.
EUROPAPARLAMENTETS OCH RÅDETS DIREKTIV 1999/92/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
1. I artikel 137 i fördraget föreskrivs att rådet genom direktiv får anta minimikrav för att, främst i fråga om arbetsmiljön främja förbättringar för att garantera en högre skyddsnivå för arbetstagares säkerhet och hälsa.
4. En förutsättning för att kunna säkerställa arbetstagarnas säkerhet och hälsa är att minimikraven för förbättring av säkerhet och hälsa för arbetstagare som kan utsättas för fara orsakad av explosiv atmosfär iakttas.
7. I Europaparlamentets och rådets direktiv 94/9/EG av den 23 mars 1994 om tillnärmning av medlemsstaternas lagstiftning om utrustning och säkerhetssystem avsedda för användning i explosionsfarliga omgivningar(5) fastställs att det på grundval av artikel 137 i fördraget skall utarbetas ett kompletterande direktiv som i synnerhet skall täcka explosionsfara till följd av användning av en viss utrustning eller till följd av typer av och metoder för installation av utrustning.
10. En bedömning av explosionsrisker kan krävas enligt annan gemenskapslagstiftning. För att undvika onödigt dubbelarbete bör arbetsgivaren, i enlighet med nationell praxis, ha möjlighet att slå ihop dokument, delar av dokument eller liknande rapporter som skall utarbetas i enlighet med annan lagstiftning till en enda säkerhetsrapport.
13. Förebyggande åtgärder måste vid behov kompletteras med andra åtgärder som genomförs när antändning har skett. Högsta möjliga skyddsnivå uppnås genom att förena förebyggande åtgärder med andra åtgärder som begränsar de skadliga effekterna för arbetstagarna av en explosion.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
2. Direktivet skall inte tillämpas på
c) framställning, hantering, användning, förvaring och transport av explosiva substanser eller instabila kemiska substanser.
3. Bestämmelserna i direktiv 89/391/EEG och de tillämpliga särdirektiven skall tillämpas fullt ut på det område som avses i punkt 1, utan att det påverkar tillämpningen av strängare och/eller mer specifika bestämmelser i det här direktivet.
I det här direktivet avses med explosiv atmosfär en blandning under atmosfäriska förhållanden av luft och brännbara ämnen i form av gas, ånga, dimma eller damm, i vilken förbränningen efter antändning sprider sig till hela den oförbrända blandningen.
Artikel 3
- förhindra att explosiv atmosfär bildas, eller, där verksamhetens art inte medger detta,
Dessa åtgärder skall vid behov kombineras och/eller kompletteras med åtgärder som förhindrar spridning av explosioner och de skall ses över regelbundet och, i alla händelser, när betydande ändringar genomförs.
1. När arbetsgivaren utför de skyldigheter som fastställs i artiklarna 6.3 och 9.1 i direktiv 89/391/EEG skall denne bedöma de särskilda risker som uppstår genom explosiv atmosfär och åtminstone ta hänsyn till
- installationerna, ämnen som används, processerna och möjlig växelverkan mellan dessa,
2. Områden som genom öppningar har eller kan få förbindelse med områden där explosiv atmosfär kan uppstå skall beaktas vid bedömningen av explosionsrisker.
För att säkerställa arbetstagarnas säkerhet och hälsa och i enlighet med de grundläggande principerna för riskbedömning och de principer som anges i artikel 3 skall arbetsgivaren vidta de åtgärder som är nödvändiga så att
Artikel 6
Utan att det åsidosätter det enskilda ansvar som varje arbetsgivare har i enlighet med direktiv 89/391/EEG skall den arbetsgivare som i enlighet med nationell lagstiftning och/eller praxis har ansvaret för arbetsplatsen samordna genomförandet av alla åtgärder om arbetstagarnas hälsa och säkerhet samt i sitt explosionsskyddsdokument, som avses i artikel 8, ange målsättningen för denna samordning liksom åtgärderna och förfarandena för genomförandet.
1. Arbetsgivaren skall klassificera områden där explosiv atmosfär kan uppstå i zoner i enlighet med bilaga I.
Artikel 8
Explosionsskyddsdokument skall särskilt innehålla uppgifter om
- de områden som har klassificerats och delats in i zoner i enlighet med bilaga I,
- att åtgärder i enlighet med rådets direktiv 89/655/EEG(10) har vidtagits så att arbetsutrustning används på ett säkert sätt.
Artikel 9
2. Arbetsutrustning, som skall användas i områden där explosiv atmosfär kan uppstå och som tillhandahålls på företaget eller i verksamheten för första gången efter den 30 juni 2003 skall uppfylla de minimikrav som fastställs i bilaga II del A och del B.
5. Om arbetsplatser med områden där explosiv atmosfär kan uppstå förändras, utvidgas eller byggs om efter den 30 juni 2003 skall arbetsgivaren vidta de åtgärder som är nödvändiga så att dessa ändringar, utvidgningar eller ombyggnader överensstämmer med de tillämpliga minimikraven i detta direktiv.
Artikel 10
- antagandet av direktiv om teknisk harmonisering och standardisering avseende området explosionsskydd, och/eller
Artikel 11
Kommissionen skall först samråda med Rådgivande kommittén för arbetarskyddsfrågor i enlighet med rådets direktiv 74/325/EEG(11).
Information till företag
Slutbestämmelser
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de redan har antagit eller antar inom det område som omfattas av detta direktiv.
KOMMISSIONENS DIREKTIV 1999/98/EG
(Text av betydelse för EES)
med beaktande av rådets direktiv 70/156/EEG av den 6 februari 1970 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av motorfordon och släpvagnar till dessa fordon(1), senast ändrat genom Europaparlamentets och rådets direktiv 98/91/EG(2), särskilt artikel 13.2 i detta,
1. Direktiv 96/79/EG är ett av särdirektiven i det förfarande för typgodkännande på gemenskapens nivå som inrättats genom direktiv 70/156/EEG. Bestämmelserna i direktiv 70/156/EEG om system, komponenter och tekniska enheter i fordonet är följaktligen tillämpliga på det här direktivet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
- förbjuda registrering, försäljning eller ibruktagande av ett fordon,
Artikel 3
2. Medlemsstaterna skall till kommissionen överlämna texten till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
av den 25 maj 1999
med hänvisning till rådets slutsatser av den 15 mars 1999, som antogs efter en fördjupad diskussion med företrädare för Europaparlamentet och kommissionen,
(2) Ansvaret för Europeiska byrån för bedrägeribekämpning, som inrättats av kommissionen, förutom skyddet av de ekonomiska intressena även omfattar all verksamhet som har samband med skyddet av gemenskapens intressen mot oegentligheten, som kan leda till administrativa eller straffrättsliga påföljder.
(5) Dessa utredningar skall utföras med iakttagande av tillämpliga bestämmelser i fördragen om upprättandet av Europeiska gemenskaperna, särskilt protokollet om immunitet och privilegier, texter som antagits för deras tillämpning samt tjänsteföreskrifterna.
efter samråd om att införa en gemensam ordning för detta ändamål, och
1. Europaparlamentet, rådet och kommissionen (nedan kallade: institutionerna) beslutar att anta en gemensam ordning för åtgärder som behövs för att underlätta att de utredningar som genomförs av byrån bedrivs på ett korrekt sätt inom institutionerna. Dessa utredningar har som ändamål att
Dessa utredningar skall genomföras med iakttagande av tillämpliga bestämmelser i fördragen om upprättandet av Europeiska gemenskaperna, särskilt protokollet om immunitet och privilegier, texter som antagits för deras tillämpning samt tjänsteföreskrifterna.
3. Institutionerna är eniga om behovet av att till byrån för yttrande överlämna varje begäran om upphävande av immunitet mot rättsliga förfaranden för tjänstemän eller anställda i samband med eventuella fall av bedrägeri, korruption eller all annan olaglig verksamhet. Om en begäran om upphävande av immunitet gäller någon av institutionernas ledamöter skall byrån underrättas.
De andra institutioner, organ och enheter som inrättats genom EG-fördraget och Euratomfördraget eller på grundval av dessa, uppmanas att ansluta sig till detta avtal genom att, var för sig, avge en förklaring som skall lämnas till ordförandena för de institutioner som undertecknat avtalet.
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande (2), och
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
"Organens faktiska utgifter skall för en treårsperiod med början på regleringsåret 1999/2000 till 50 % täckas av gemenskapernas allmänna budget.
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Enligt kompletterande uppgifter som lämnats a
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
Enligt omfattande forskning och vetenskapliga studier bevaras näringsvärdet, särskilt betakarotinhalten, i en produkt av hög kvalitet om torkningen av fodret äger rum vid hög temperatur.
För de tekniska justeringar som är nödvändiga i detta syfte krävs en bekräftelse på att den behöriga myndigheten godkänt företaget.
Förvaltningskommittén för torkat foder har inte avgivet något yttrande inom den tid som dess ordförande har bestämt.
Förordning (EG) nr 785/95 ändras på följande sätt:
1. De tekniska justeringar i torkningsanläggningarna som är nödvändiga enligt bestämmelserna i artikel 1.1 skall göras utan att det påverkar kravet om att underrätta den behöriga myndigheten inom den tidsfrist som anges i artikel 4.1 a sista stycket i förordning (EG) nr 785/95.
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om handelsnormer för morötter
med beaktande av rådets förordning (EEG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom kommissionens förordning (EG) nr 2520/97(2), särskilt artikel 2.2 i denna, och
Syftet med dessa normer är att avlägsna produkter av otillfredsställande kvalitet från marknaden, att styra produktionen på ett sådant sätt att den uppfyller konsumenternas krav samt att underlätta handelsförbindelserna på grundval av sund konkurrens och därigenom bidra till att förbättra lönsamheten.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Dessa normer skall tillämpas i samtliga handelsled och i enlighet med villkoren i förordning (EG) nr 2200/96.
- uppvisa mindre förändringar till följd av sin utveckling och benägenhet att förfaras, dock inte om de klassificerats som klass "Extra".
1) I artikel 1 första stycket skall första strecksatsen utgå.
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om öppnande och förvaltning av tullkvoter för import av tjurar, kor och kvigor av vissa alp- och bergraser som inte är slaktboskap, om upphävande av förordning (EG) nr 1012/98 och om ändring av förordning (EG) nr 1143/98
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött(1), senast ändrad genom förordning (EG) nr 1633/98(2), särskilt artikel 12.1 i denna,
(1) Inom ramen för Världshandelsorganisationen (WTO) har gemenskapen åtagit sig att öppna två tullkvoter med en årlig kvantitet på 5000 djur vardera med en tull på 6 % respektive 4 %. Tullkvoterna gäller tjurar, kor och kvigor av brokig Simmentalras och Schwyz- och Fribourgras som inte är slaktboskap samt kor och kvigor av grå, brun, gul och brokig Simmentalras och Pinzgauras som inte är slaktboskap. Dessa kvoter bör öppnas på flerårsbasis för perioder om tolv månader, nedan kallade importår, som inleds den 1 juli, och tilllämpningsföreskrifter bör fastställas.
(4) För att inte förorsaka alltför stor stelhet i handelsförbindelserna inom sektorn bör dock ytterligare en kvantitet ställas till förfogande för sådana importörer som kan visa att de bedriver seriös verksamhet och handlar med betydande kvantiteter med tredje land. För detta ändamål och för att säkerställa en effektiv förvaltning är det lämpligt att kräva att de berörda aktörerna skall ha importerat minst 15 djur under de tolv månader som föregår importåret i fråga. Ett parti på 15 djur utgör i princip en normal last och erfarenheten har visat att försäljning eller inköp av ett enstaka parti utgör ett minimikrav för att en transaktion skall kunna betraktas som reell och ekonomiskt lönsam.
(7) Det bör föreskrivas att importtillstånden skall fördelas efter en viss betänketid och eventuellt med tillämpning av en enhetlig procentsats för nedsättning.
(10) Kommissionens förordning (EG) nr 1012/98 av den 14 maj 1998 om öppnande och förvaltning av tullkvoter för import av tjurar, kor och kvigor av vissa alp- och bergraser som inte är slaktboskap(12), senast ändrad genom förordning (EG) nr 1143/98(13), bör upphävas.
(13) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för nötkött.
1. För en flerårsperiod skall under perioden 1 juli-30 juni följande år, nedan kallad importåret, följande tullkvoter öppnas:
Undantag kan emellertid beviljas i vederbörligen styrkta fall av force majeure.
- För kor och kvigor: En stamtavla eller ett intyg om registrering i stamboken som styrker rasrenheten.
a) Den första delen av varje kvot om 80 % skall fördelas mellan importörer från gemenskapen som kan styrka att de har importerat djur som omfattas av kvoter med löpnummer 09.0001 och/eller 09.0003 under de 36 månader som föregåJar importåret i fråga.
Importörerna skall vara registrerade i ett nationellt register för mervärdesskatt.
Ansökan om importtillstånd
Ansökningar om importtillstånd för mer än 50 djur skall automatiskt sänkas till detta antal.
Artikel 3
Artikel 4
Om en sökande lämnar in mer än en ansökan för en enskild kvot, skall inga ansökningar från denne sökande för den aktuella kvoten godtas.
- När det gäller den ordning som avses i artikel 2.1 a första stycket, en förteckning över de importörer som uppfyller villkoren för godkännande, med uppgift om deras namn och adress samt antalet importerade djur under den period som avses i artikel 2.2.
Artikel 5
Om den minskning som avses i första stycket resulterar i en kvantitet på mindre än 15 djur per ansökan, skall partier på 15 djur fördelas genom lottdragning av de berörda medlemsstaterna. Om den återstående kvantiteten uppgår till mindre än 15 djur, skall den kvantiteten utgöra ett enda parti.
2. Ansökan om importlicens får endast lämnas in till den behöriga myndigheten i den medlemsstat där den sökande har ansökt om importtillstånd.
5. De utfärdade licenserna skall vara giltiga i hela gemenskapen.
8. Artikel 8.4 i förordning (EEG) nr 3719/88 skall inte tillämpas.
2. För att garantera att skyldigheten enligt punkt 1 att inte slakta djuren efterlevs, och för att säkerställa uppbörden av obetalda tullar om denna skyldighet inte fullgörs, skall en säkerhet ställas hos de behöriga myndigheterna. Denna säkerhet skall motsvara skillnaden mellan de tullar som fastställts i den gemensamma tulltaxan och de tullar som avses i artikel 1.1 och som är tillämpliga den dag då djuren i fråga övergår till fri omsättning.
Artikel 8
b) I fält 16, de KN-nummer som anges i bilaga I.
Artikel 9
3. Kommissionen skall snarast möjligt besluta om dessa återstående kvantiteter.
5. Endast en ansökan per kvot får lämnas in av en och samme aktör.
7. För varje löpnummer skall medlemsstaterna senast den sjunde dagen efter det att den period för inlämnande av ansökningar som anges i punkt 6 gått till ända till kommissionen överlämna en förteckning över de sökande och vilka kvantiteter de har ansökt om.
förordning (EG) nr 1012/98 upphör att gälla.
1) Artikel 2.1 a andra stycket skall ersättas med följande: "Medlemsstaterna får emellertid som referenskvantiteter godkänna importtillstånd som hänför sig till föregående importår men som inte har delats ut om detta beror på ett administrativt fel som begåtts av den nationella behöriga myndigheten."
- Bjergracer (forordning (EF) nr. 1143/98), importår: ...
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av kommissionens förordning (EG) nr 111/1999 om tillämpningsföreskrifter för rådets förordning (EG) nr 2802/98 om ett program för leverans av jordbruksprodukter till Ryska federationen
med beaktande av rådets förordning (EG) nr 2802/98 av den 17 december 1998 om ett program för leverans av jordbruksprodukter till Ryska federationen(1), särskilt artikel 4.2 i denna, och av följande skäl:
(3) Beträffande bearbetade produkter på basis av produkter från interventionslager eller på basis av produkter som anskaffats på gemenskapsmarknaden bör bestämmelserna om intyg om överensstämmelse ändras, särskilt när det gäller hur kontrollerna organiseras, och det bör fastställas mer detaljerade bestämmelser för hur den aktör som innehar kontraktet för transport av varorna utanför gemenskapen skall överta produkterna.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandena från samtliga berörda förvaltningskommittéer.
Förordning (EG) nr 111/1999 ändras på följande sätt:
9) I artikel 5.1 i skall "i enlighet med den förlaga som återfinns i bilaga III" ersättas med "i enlighet med den förlaga som återfinns i bilaga IV".
1. För de leveranser som avser produktion av helt slipat ris eller anskaffande av griskött på gemenskapsmarknaden skall kontraktsinnehavaren erhålla ett fast belopp på 0,45 euro per ton (netto) och dag för ris och på 0,90 euro per ton (netto) och dag för griskött för att täcka alla omkostnader (parkering, försäkring, bevakning, säkerhet, osv.) som uppstår i de fall då transportören utan egen förskyllan inte kan agera inom de föreskrivna tidsramarna.
1. Begäran om betalning för leveransen skall inlämnas till det interventionsorgan som avses i artikel 4 inom två månader från utgången av den leveransperiod som fastställs i anbudsinfordran. Om denna bestämmelse inte iakttas, med undantag för fall av force majeure, skall beloppet minskas med 10 % för den första månadens försening. Vid ytterligare försening skall beloppet minskas med 5 % per månad.
- en kopia av transportdokumenten,
- en kopia av exportlicensen eller exportdeklarationen, i de fall då det enligt lagstiftningen beträffande den gemensamma organisationen av marknaden inte krävs någon exportlicens,
4. Vid anbudsförfarande enligt artikel 2.2 skall den kvantitet interventionsprodukter för vilken anbudsgivaren tilldelats kontrakt ställas till dennes förfogande när det har styrkts att det ställts säkerhet i enlighet med artikel 7.2.
"3. Om det vid leveransstadiet kan konstateras att förseningar har uppstått skall 0,75 euro per ton av leveranssäkerheten förverkas för varje dags försening av den del av kvantiteten som lastats eller levererats för sent. Om sådana förseningar överstiger elva dagar skall avdraget ökas till 1 euro per ton för varje ytterligare dag. Dessa bestämmelser skall tillämpas när kontraktsinnehavaren är ansvarig för förseningen av lastningen eller leveransen."
Exportlicensen skall utfärdas endast om det bevisas att den leveranssäkerhet som avses i artikel 7 har ställts. Ställandet av denna säkerhet skall anses utgöra ställandet av licenssäkerheten. Trots bestämmelserna i avdelning III avsnitt 4 i förordning (EEG) nr 3719/88 skall säkerheten frisläppas på de villkor som fastställs i artikel 12.2."
Artikel 2
av den 16 juni 1999
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(2) I flera medlemsstater har försök i stor skala gjorts med en ny fodertillsats, "natrolit-fonolit" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel". Med hänsyn till de erfarenheter som har gjorts bör denna nya fodertillsats kunna tillåtas.
(5) Det tillfälliga godkännandet av "natrolit-fonolit" slutade gälla redan den 21 april 1999. Av rättssäkerhetsskäl är det därför nödvändigt att denna förordning tillämpas retroaktivt.
Artikel 1
"Hydratiserad kalciumaluminiumsilikat av vulkaniskt ursprung" i gruppen "Bindemedel, klumpförebyggande medel och koaguleringsmedel" får tillåtas enligt direktiv 70/524/EEG som fodertillsats nr 3 på de villkor som anges i bilaga II till den här förordningen.
RÅDETS FÖRORDNING (EG) nr 1258/1999
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europaparlamentets yttrande(2),
av följande skäl: 1. Genom förordning nr 25 om finansieringen av den gemensamma jordbrukspolitiken(5) upprättade rådet Europeiska utvecklings- och garantifonden för jordbruket (EUGFJ), nedan kallad "fonden", som utgör en del av Europeiska gemenskapernas allmänna budget. I den förordningen fastställs de principer som skall tillämpas för finansieringen av den gemensamma jordbrukspolitiken.
4. Kommissionen ansvarar för förvaltningen av fonden. Ett nära samarbete mellan medlemsstaterna och kommissionen i en kommitté för Europeiska utvecklings- och garantifonden för jordbruket föreskrivs.
7. Ett decentraliserat förvaltningssystem för gemenskapens fonder innebär, särskilt efter reformen av den gemensamma jordbrukspolitiken, att flera utbetalningsställen kan utses. När en medlemsstat ackrediterar fler än ett utbetalningsställe måste den därför utse ett enda kontaktorgan för att säkerställa konsekvens av fondernas förvaltning, upprätta kontakter mellan kommissionen och de olika ackrediterade utbetalningsställena och säkerställa att sådana uppgifter om olika utbetalningsställens transaktioner som kommissionen begär skall kunna göras tillgängliga med kort varsel.
10. Granskningen av överensstämmelse och därpå följande beslut om ackreditering kommer således inte längre att vara knutna till verkställandet av budgeten för ett visst budgetår. Det är nödvändigt att fastställa den längsta period som slutsatserna av granskningen av överensstämmelse kan avse. Åtgärderna för landsbygdsutveckling är emellertid fleråriga, vilket gör att det inte är möjligt att tillämpa en sådan längsta period.
13. Det är nödvändigt att i största möjliga utsträckning använda informationsteknik för att få fram den information som skall sändas till kommissionen. När kommissionen utför kontroller måste den ha fullständig och omedelbar tillgång till uppgifter som rör utgifter, både i dokument och i datafiler.
16. Rådets förordning (EEG) nr 729/70 av den 21 april 1970 om finansiering av den gemensamma jordbrukspolitiken(7) har ändrats i betydande omfattning vid ett flertal tillfällen. Nu när nya ändringar görs av nämnda förordning är det önskvärt att bestämmelserna i fråga omarbetas för att förtydliga vissa frågor.
- Garantisektionen.
a) bidrag vid export till tredje land,
d) gemenskapens finansiella bidrag till särskilda veterinära åtgärder, kontrollåtgärder på veterinärområdet och program för bekämpning och övervakning av djursjukdomar (veterinära åtgärder) samt till växtskyddsåtgärder,
4. Utgifter för administration och personal som belastar medlemsstater och mottagare av stöd från fonden skall inte finansieras av fonden.
2. Intervention för att stabilisera jordbruksmarknaderna som görs i enlighet med gemenskapsbestämmelser inom ramen för den gemensamma organisationen av jordbruksmarknaderna skall finansieras enligt artikel 1.2 b.
1. Åtgärder för landsbygdsutveckling utanför mål 1-programmen som vidtas enligt gemenskapsbestämmelser skall finansieras enligt artikel 1.2 c.
4. Tillämpningsföreskrifter för denna artikel skall antas i enlighet med förfarandet i artikel 13.
a) De myndigheter och organ som den ackrediterar för att göra de betalningar som avses i artiklarna 2 och 3, nedan kallade "utbetalningsställen".
a) ansökningarnas berättigande och överensstämmelse med gemenskapsbestämmelserna kontrolleras innan betalningarna godkänns,
3. Utbetalningsställena skall inneha verifikationshandlingar avseende de gjorda utbetalningarna och handlingar som gäller genomförandet av de föreskrivna administrativa och fysiska kontrollerna. Om de relevanta handlingarna förvaras hos de organ som har till uppgift att godkänna utgifterna, skall dessa organ tillställa utbetalningsstället rapporter om antalet genomförda kontroller, dessas innehåll och de åtgärder som har vidtagits mot bakgrund av resultaten.
6. Varje medlemsstat skall till kommissionen överlämna följande upplysningar om utbetalningsställena:
c) Ackrediteringshandlingen.
8. Tillämpningsföreskrifterna för denna artikel skall antas i enlighet med förfarandet i artikel 13.
Förskottsbetalning för genomförande av program inom ramen för de åtgärder för landsbygdsutveckling som avses i artikel 3.1 får beviljas av kommissionen när dessa program godkänns och skall betraktas som utgifter som verkställts den första dagen i månaden efter beslutet om beviljandet.
Artikel 6
b) Årsredovisningen tillsammans med nödvändiga underlag för granskning och godkännande samt ett intyg avseende den vidarebefordrade redovisningens fullständighet, exakthet och sanningsenlighet.
1. Efter att ha hört fondkommittén skall kommissionen fatta de beslut som anges i punkterna 2, 3 och 4.
Ytterligare förskott får göras om fondkommittén underrättas vid nästa samråd.
4. Kommissionen skall besluta om vilka utgifter som inte skall omfattas av gemenskapsfinansiering enligt artiklarna 2 och 3 om den finner att utgifterna inte har verkställts i överensstämmelse med gemenskapsbestämmelserna.
Kommissionen skall göra en bedömning av de belopp som skall undantas, särskilt med hänsyn till hur stor bristen på överensstämmelse är. Kommissionen skall beakta överträdelsens art och betydelse samt den ekonomiska förlust som gemenskapen lidit.
b) De utgifter för åtgärder som avses i artikel 3 och där den slutliga betalningen verkställdes före de tjugofyra månader som föregick kommissionens skriftliga meddelande till den berörda medlemsstaten om resultaten av kontrollerna.
b) av statligt stöd eller överträdelser för vilka förfarandena som anges i artiklarna 88 och 226 i fördraget har inletts.
1. Medlemsstaterna skall i enlighet med nationella bestämmelser i lagar och andra författningar vidta de åtgärder som är nödvändiga för att
c) indriva belopp som förlorats till följd av oegentligheter eller försumlighet.
De indrivna beloppen skall betalas till de ackrediterade utbetalningsställena och dessa organ skall dra av de indrivna beloppen från de utgifter som fonden finansierar. Räntan på de belopp som drivits in eller som betalats för sent skall betalas in till fonden.
1. Medlemsstaterna skall till kommissionens förfogande ställa alla uppgifter som behövs för att fonden skall fungera väl och de skall även vidta alla lämpliga åtgärder för att underlätta den kontroll som kommissionen kan anse vara nödvändig inom ramen för förvaltningen av gemenskapsfinansieringen, inbegripet kontroller på plats.
De får särskilt kontrollera
c) under vilka förhållanden transaktioner som finansieras av fonden genomförs och kontrolleras.
För att effektivisera kontrollen får kommissionen, med de berörda medlemsstaternas samtycke, ombesörja att myndigheter i dessa stater deltar i vissa kontroller eller utredningar.
Före den 1 juli varje år skall kommissionen tillställa Europaparlamentet och rådet en finansiell rapport om förvaltningen av fonden under det föregående räkenskapsåret, särskilt dess ekonomiska ställning och utvecklingen av utgifternas storlek och utgiftsslagen samt förutsättningarna för gemenskapsfinansieringens genomförande.
Artikel 12
1. Om förfarandet i denna artikel skall tillämpas skall ordföranden, antingen på eget initiativ eller på begäran av en företrädare för en medlemsstat, hänskjuta ärendet till fondkommittén.
b) Om beslutet inte är förenligt med fondkommitténs yttrande skall kommissionens emellertid genast underrätta rådet. I sådana fall
Artikel 14
b) angående den bedömning av fondens anslag som skall skrivas in i kommissionens upskattning för kommande budgetår och vid behov i ytterligare budgetsförslag,
Fondkommittén skall regelbundet informeras om fondens verksamheter.
Kommissionen skall ställa sekretariatstjänster till fondkommitténs förfogande.
1. Förordning (EEG) nr 729/70 skall upphävas.
Artikel 15 tredje stycket och artikel 40 i beslut 90/424/EEG skall utgå.
Artikel 19
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
2. Genom undantag från direktiv 70/524/EEG tillåts medlemsstaterna genom rådets direktiv 93/113/EG av den 14 december 1993 om användning och saluföring av enzymer och mikroorganismer och preparat av dessa i djurfoder(3), senast ändrat genom rådets direktiv 97/40/EG(4), att tillfälligt tillåta användning och saluföring av enzymer, mikroorganismer och preparat av dessa i foder.
5. En granskning av de akter som medlemsstaterna har överlämnat i enlighet med artikel 3 i direktiv 93/113/EG ger vid handen att vissa preparat av typen enzymer och mikroorganismer kan godkännas tills vidare.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
om klassificering av vissa varor i Kombinerade nomenklaturen
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom kommissionens förordning (EG) nr 1835/1999(2), särskilt artikel 9 i denna, och
2. I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
5. De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från tullkodexkommittén.
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 3
av den 3 december 1999
med beaktande av rådets direktiv 70/524/EEG av den 23 november 1970 om fodertillsatser(1), senast ändrat genom kommissionens förordning (EG) nr 2439/1999(2), särskilt artiklarna 9h.3 b och 9i.3 b i detta, och
2. Efter den 31 december 1987 skall, särskilt enligt artikel 9h i direktiv 70/524/EEG, de preliminära godkännandena för tillsatser som avses i bilaga I och som hör till gruppen antibiotika och som förts över till bilaga B, kapitel II ersättas med godkännanden som knyts till den som är ansvarig för avyttringen för en tid av tio år.
5. Godkännandet knyts till en person som är ansvarig för avyttringen på grundval av rent administrativa förfaranden och innebär inte någon ny utvärdering av tillsatserna. Även om godkännandena enligt denna förordning beviljas för en viss tid, kan de när som helst återkallas enligt artikel 9m och artikel 11 i direktiv 70/524/EEG. De kan särskilt återkallas mot bakgrund av följande: Vetenskapliga styrkommittén avgav den 28 maj 1999 ett yttrande om antimikrobiell resistens. Användningen av vissa antibiotika i foder håller för närvarande på att utvärderas på nytt enligt artikel 9g i direktiv 70/524/EEG. Sverige har på grundval av artikel 11 i direktiv 70/524/EEG inom sitt territorium förbjudit användningen av alla former av antibiotika som tillsats i foder. Kommissionen håller dessutom på att gå igenom de data som lämnats in och den mer allmänna frågan huruvida användningen av antibiotika som tillsats i foder uppfyller de villkor som föreskrivs i artikel 3a i direktiv 70/524/EEG för att godkännande som tillsats skall meddelas.
Artikel 1
De preliminära godkännandena av de tillsatser som förtecknas i bilaga II till denna förordning skall ersättas med preliminära godkännanden som knyts till den som är ansvarig för avyttringen av tillsatserna och som anges i andra kolumnen i bilaga II.
KOMMISSIONENS FÖRORDNING (EG) nr 2654/1999
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) skummjölk: mjölk från en eller flera kor eller getter, fri från tillsatser och som endast genomgått partiell skumning, så att fetthalten sjunkit till högst 0,10 %,
d) kaseinater: de produkter som erhålls genom torkning av kasein eller råkasein som behandlats med neutraliserande agens."
CENTRALGRUPPENS BESLUT
(SCH/C (99) 25)
KOMMISSIONENS BESLUT
[delgivet med nr K(1999) 4749]
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
2. Villkoren för import av musslor, tagghudingar, manteldjur och marina snäckor och sniglar med ursprung i Chile fastställs i kommissionens beslut 96/675/EG(5).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 9 mars 2000
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(3) I enlighet med artikel 7.1 c i förordning (EEG) nr 3600/92 ingav Förenade kungariket, som utsetts till rapporterande medlemsstat, den 30 april 1996 en rapport till kommissionen om sin utvärdering av de uppgifter som anmälarna lämnat enligt artikel 6.1 i den förordningen.
(6) Den enda anmälaren har informerat kommissionen och den rapporterande medlemsstaten om att denne inte längre önskar delta i arbetsprogrammet för detta verksamma ämne. Viktiga delar av den information som krävs för att uppfylla kraven i direktiv 91/414/EEG kommer därför inte att överlämnas.
(9) Detta beslut påverkar inte de eventuella åtgärder som kommissionen kan vidta i ett senare skede med hänsyn till detta verksamma ämne inom ramen för rådets direktiv 79/117/EEG(7).
Artikel 1
Medlemsstaterna skall garantera att
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
om ändring av bilaga IV till rådets direktiv 90/539/EEG om djurhälsovillkor för handel inom gemenskapen med och för import från tredje land av fjäderfä och kläckningsägg och om ändring av beslut 96/482/EG om djurhälsovillkor och veterinärintyg för import från tredje land av fjäderfä och kläckningsägg, med undantag av strutsfåglar och ägg från strutsfåglar, inbegripet djurhälsoåtgärder som skall vidtas efter sådan import
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av rådets direktiv 91/496/EEG av den 15 juli 1991 om fastställande av regler för hur veterinärkontroller skall organiseras för djur som importeras till gemenskapen från tredje land och om ändring av direktiven 89/662/EEG, 90/425/EEG och 90/675/EEG(3), senast ändrat genom direktiv 96/43/EG(4), särskilt artikel 10 i detta, och
(2) Med hänsyn till de erfarenheter som gjorts vid tillämpningen av de föreskrivna åtgärderna bör villkoren för handel inom gemenskapen med dagsgamla kycklingar från kläckägg som importerats från tredje land ändras. Genom ändringen bör det bli möjligt för medlemsstaterna att sända dagsgamla kycklingar till anläggningar i en annan medlemsstat under förutsättning att kycklingarna isoleras efter import.
(5) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Förlaga 2 i bilaga IV till direktiv 90/539/EEG skall ersättas med bilagan till detta beslut.
Artikel 2
Detta beslut riktar sig till alla medlemsstater.
enligt Europaparlamentets och rådets direktiv 95/46/EG om huruvida ett adekvat skydd säkerställs genom de principer om integritetsskydd (Safe Harbor Privacy Principles) i kombination med frågor och svar som Förenta staternas handelsministerium utfärdat
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Enligt direktiv 95/46/EG skall medlemsstaterna föreskriva att överföring av personuppgifter till tredje land endast får ske om ifrågavarande tredje land säkerställer en adekvat skyddsnivå och om medlemsstatens lagar genom vilka andra bestämmelser i direktivet genomförs, efterlevs före överföringen.
(4) Mot bakgrund av de olika sätten att se på frågan om uppgiftsskydd i olika tredje länder bör bedömningen av om skyddsnivån är adekvat ske, och beslut som grundar sig på artikel 25.6 i direktiv 95/46/EG verkställas, utan godtycklig eller obefogad diskriminering i förhållande till tredje land eller mellan tredje länder där liknande förhållanden råder och så att det inte utgör ett dolt handelshinder. Härvid bör hänsyn tas till gemenskapens nuvarande internationella åtaganden.
(7) För att se till att detta beslut tillämpas korrekt är det nödvändigt att de organisationer som ansluter sig till principerna och FoS kan erkännas av berörda parter, t.ex. de registrerade, exportörer av uppgifter och dataskyddsmyndigheter. I detta syfte bör Förenta staternas handelsministerium, eller det organ som ministeriet bestämmer, förbinda sig att föra och göra tillgänglig för allmänheten en förteckning över de organisationer som förpliktat sig att följa principerna i överensstämmelse med FoS och som lyder under åtminstone en av de myndigheter som nämns i bilaga VII till detta beslut.
(10) Arbetsgruppen för skydd av enskilda med avseende på behandling av personuppgifter som inrättats genom artikel 29 i direktiv 95/46/EG har avgivit yttranden om den skyddsnivå som erbjuds av safe harbor-principerna i Förenta staterna, och vid utarbetandet av föreliggande beslut har hänsyn tagits till dessa yttranden(4).
Artikel 1
b) Ett memorandum om ersättning vid kränkning av enskildas integritet och uttryckliga behörigheter i Förenta staternas lagstiftning, bilaga IV.
2. I samband med varje överföring av uppgifter skall följande villkor vara uppfyllda:
3. De villkor som anges i punkt 2 skall anses vara uppfyllda för varje organisation som genom självcertifiering förbinder sig att följa principerna i överensstämmelse med FoS från den dag då organisationen underrättar Förenta staternas handelsministerium, eller det organ som ministeriet bestämmer, om offentliggörandet av den förpliktelse som avses i punkt 2 a och om namnet på den myndighet som avses i punkt 2 b.
Artikel 3
b) det är i hög grad sannolikt att principerna överträds, det finns välgrundad anledning att tro att den berörda instansen för handläggning av klagomål inte vidtar och inte i rätt tid kommer att vidta de åtgärder som behövs för att lösa problemet, en fortsatt överföring av uppgifterna skulle innebära en överhängande risk för allvarlig skada för registrerade, och de behöriga myndigheterna i medlemsstaten har gjort vad som under rådande omständigheter rimligvis kan krävas för att anmärka mot organisationen och ge den tillfälle att gå i svaromål.
3. Medlemsstaterna och kommissionen skall även underrätta varandra om varje fall där en myndighet, som är ansvarig för att principerna tillämpade i överensstämmelse med FoS följs i Förenta staterna, inte kunnat säkerställa detta.
2. Kommissionen skall om så behövs föreslå åtgärder i enlighet med det förfarande som föreskrivs i artikel 31 i direktivet.
Artikel 6
av den 6 september 2000
(2000/540/EG)
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(1), senast ändrat genom kommissionens direktiv 2000/10/EG(2), särskilt artikel 6.3 i detta, och
(2) Företaget Rohm & Haas France SA lämnade den 2 juni 1999 in en akt med dokumentation för det verksamma ämnet RH-7281 (zoxamid) till myndigheterna i Förenade kungariket för införande av detta verksamma ämne i bilaga I till direktivet.
(5) Företaget Aventis GmbH lämnade den 30 mars 2000 in en akt med dokumentation för det verksamma ämnet AEF130360 (foramsulfuron) till de tyska myndigheterna.
(8) Enligt artikel 6.3 i direktivet krävs en bekräftelse på gemenskapsnivå av att varje akt med dokumentation uppfyller kraven på faktauppgifter och upplysningar enligt bilaga II och, vad beträffar åtminstone ett växtskyddsmedel som innehåller det verksamma ämnet i fråga, enligt bilaga III till direktivet.
(11) Medlemsstaterna och kommissionen har enats om att Förenade kungariket skall fortsätta att noggrant granska dokumentationen om RH-7281 (zoxamid), att Nederländerna skall fortsätta att noggrant granska dokumentationen om B-41; E-187 (milbemectin) och att Tyskland skall fortsätta att noggrant granska dokumentationen om BAS500F (pyraclostrobin) och AEF130360 (foramsulfuron).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Den dokumentation som lämnats in av Rohm & Haas France SA till kommissionen och medlemsstaterna beträffande införandet av RH-7281 (zoxamid) som ett verksamt ämne i bilaga I till direktiv 91/414/EEG, och som överlämnades till Ständiga kommittén för växtskydd den 31 maj 2000.
4. Den dokumentation som lämnats in a
om tillnärmning av medlemsstaternas lagstiftning om märkning och presentation av livsmedel samt om reklam för livsmedel
med beaktande av kommissionens förslag,
av följande skäl:
(3) Det är därför nödvändigt att närma dessa lagstiftningar till varandra för att bidra till att den inre marknaden fungerar smidigare.
(6) Det huvudsakliga syftet med regler om märkning av livsmedel bör vara behovet att informera och skydda konsumenten.
(9) En förteckning bör därför göras upp över alla uppgifter som i princip bör framgå av märkningen på alla livsmedel.
(12) En sådan procedur måste utgöras av ett gemenskapsbeslut, när en medlemsstat önskar att införa ny lagstiftning.
(15) I syfte att underlätta handeln mellan medlemsstaterna får det i handelsleden före försäljningen till konsumenter tillåtas att endast den viktigaste informationen framgår av den yttre förpackningen och att vissa obligatoriska uppgifter som måste finnas på ett färdigförpackat livsmedel behöver framgå endast av handelsdokument som rör detta.
(18) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(5).
2. Detta direktiv gäller även livsmedel avsedda för restauranger, sjukhus; personalrestauranger och andra liknande storkök (i det följande benämnda storkök).
b) färdigförpackat livsmedel: varje enskild vara som i oförändrat skick är avsedd att tillhandahållas konsumenter och storkök och som består av ett livsmedel och den förpackning i vilket det placerades innan det erbjöds till försäljning, oavsett om förpackningen omsluter livsmedlet helt eller endast delvis, men förutsatt att förpackningen omsluter livsmedlet på sådant sätt att innehållet inte kan ändras utan att förpackningen öppnas eller ändras.
a) vara sådan att den på ett avgörande sätt skulle kunna vilseleda köparen, i synnerhet
iii) genom att antyda att livsmedlet har speciella egenskaper, då i själva verket alla liknande livsmedel har sådana egenskaper,
3. De förbud och begränsningar som avses i punkterna 1 och 2 skall gälla också
Artikel 3
2. Ingrediensförteckning.
5. Datum för minsta hållbarhetstid eller, när det gäller livsmedel som ur mikrobiologisk synpunkt är lättfördärvliga, datum för sista förbrukningsdag.
Medlemsstaterna skall dock ha rätt att i fråga om smör som framställts inom deras territorium, kräva uppgift endast om tillverkaren, förpackaren eller säljaren.
9. Bruksanvisning, om det utan en sådan skulle vara omöjligt att använda livsmedlet på rätt sätt.
3. Bestämmelserna i denna artikel skall inte påverka tillämpningen av mer precisa eller långtgående bestämmmelser om mått och vikt.
3. De gemenskapsbestämmelser som avses i punkterna 1 och 2 skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
a) Om gemenskapen saknar bestämmelser skall försäljningsnamnet vara det namn som föreskrivs i lag eller andra författningar som gäller i den medlemsstat i vilken varan säljs till konsumenter eller till institutioner och storkök.
I fall där övriga bestämmelser i detta direktiv, särskilt de i artikel 3, inte är tillräckliga för att säkerställa att konsumenterna i den medlemsstat där produkten saluförs har kännedom om produktens verkliga art och kan särskilja det från produkter som det skulle kunna förväxlas med, skall försäljningsnamnet emellertid kompletteras med ytterligare beskrivande information bredvid namnet.
3. Det namn under vilket varan säljs skall omfatta eller åtföljas av uppgifter om livsmedlets fysiska tillstånd eller den särskilda behandling som livsmedlet fått (t.ex. pulvrisering, frystorkning, djupfrysning, koncentrering, rökning) i samtliga fall då avsaknaden av sådan information skulle kunna skapa förvirring hos köparen.
"irradiado" eller "tratado con radiación ionizante"
- på tyska:
"irradiated" eller "treated with ionizing radiation"
- på italienska:
"doorstraald" eller "door bestraling behandeld" eller "met ioniserende stralen behandeld"
- på finska:
"bestrålad" eller "behandlad med joniserande strålning."
2. Ingredienser behöver inte anges beträffande
- mikrobiellt framställd ättika som utvunnits ur en enda basprodukt coh som inte fillsatts någon annan ingrediens,
- kulturmjölk och syrad grädde,
- om försäljningsnamnet är identiskt med nammet på ingrediensen, eller
4. a) Med ingrediens menas varje ämne, inklusive tillsatser, som använts i tillverkningen eller beredningen av ett livsmedel och som finns kvar i den färdiga produkten, om än i annan form.
i) beståndsdelarna av en ingrediens som under framställningsprocessen tillfälligt avskiljts men senare åter tillförts livsmedlet i proportioner som inte överskrider de ursprungliga,
- som används som processhjälpmedel,
5. Ingrediensförteckningen skall omfatta samtliga ingredienser i livsmedlet i fallande storleksordning efter den vikt som ingrediensen hade vid framställningstidpunkten. Den skall föregås av en lämplig rubrik som innehåller ordet "ingredienser".
- Ingredienser som använts i koncentrerad eller torkad form och som under framställningen rekonstitueras får anges i storleksordning efter den vikt som ingredienserna hade innan de koncentrerades eller torkades.
- Ingredienserna i krydd- eller örtblandningar, i vilka ingen krydda eller ört påtagligt dominerar med hänsyn till vikt får anges i annan ordning, förutsatt att ingrediensförteckningen följs av uttrycket "i varierande proportion" eller liknande uttryck.
- Ingredienser som tillhör någon av de i bilaga 1 uppräknade kategorierna och som är beståndsdelar i ett annat livsmedel, behöver anges endast med namnet på denna kategori.
- Ingredienser som tillhör någon av de i bilaga II uppräknade kategorierna skall alltid anges med namnet på denna kategori åtföljt av deras särskilda beteckning eller E-nummer. Om en ingrediens tillhör mer än en av kategorierna skall den kategori anges som är lämpligast med hänsyn till ingrediensens huvudsakliga funktion i det aktuella livsmedlet.
- Aromer skall benämnas enligt bilaga III.
Det förfarande som fastställs i artikel 19 skall tillämpas på varje sådan nationell bestämmelse.
En sådan förteckning skall dock inte vara obligatorisk i följande fall:
9. Utan hinder av punkt 5 behöver innehållet av vatten inte anges särskilt
Artikel 7
a) om den berörda ingrediensen eller kategorin av ingredienser ingår i försäljningsnamnet eller vanligtvis förknippas med det namnet av konsumenterna, eller
d) i de fall som fastställs i enlighet med det förfarande som anges i artikel 20.2.
- vars avrunna nettovikt anges i enlighet med artikel 8.4,
- som trots att den ingår i försäljningsnamnet inte kommer att styra konsumenternas val i den medlemsstat där saluföringen sker, då variationen i mängd inte är avgörande för att känneteckna livsmedlet eller är sådan att den särskiljer livsmedlet från liknande varor; enligt förfarandet i artikel 20.2 skall det i tveksamma fall avgöras om villkoren i denna strecksats är uppfyllda,
d) i de fall som fastställs i enlighet med det förfarande som anges i artikel 20.2
6. Denna artikel skall tillämpas utan att det påverkar tilllämpningen av gemenskapens regler om näringsvärdesdeklaration.
- i volymenheter i fråga om vätskor,
Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser, som gäller för vissa livsmedel, får avvika från denna regel.
Utan att det påverkar den anmälningsskyldighet som föreskrivs i artikel 24, skall medlemsstaterna underrätta kommissionen och de andra medlemstaterna om varje åtgärd som vidtagits enligt denna punkt.
c) Om en färdigförpackad vara består av två eller flera separata färdigförpackningar som innehåller samma mängd av samma vara, skall nettoinnehållet anges genom uppgift om nettoinnehållet för varje separat förpackning och det totala antalet sådana förpackningar. Dessa uppgifter är dock inte obligatoriska, om det totala antalet separata förpackningar är klart synligt och lätt kan räknas utifrån, och om minst en uppgift om nettoinnehållet i varje enskild förpackning är klart synlig från utsidan.
3. När det gäller livsmedel som normalt säljs styckevis behöver medlemsstaterna inte kräva uppgift om nettoinnehållet under forutsättning att antalet artiklar är klart synliga och lätt räknas utifrån eller, om detta inte är möjligt, framgår av märkningen.
I denna punkt avses med en "lag" följande varor, eventuellt i blandningar och även i fryst eller djupfryst tillstånd, förutsatt att vätskan bara är ett komplement till den aktuella beredningens viktiga beståndsdelar och således inte en för köpet avgörande faktor: vatten, saltlösningar, saltlake; livsmedelssyror lösta i vatten, ättika; sockerlag, vattenlösningar med andra sötningsmedel; i fråga om frukt eller grönsaker, frukt- eller grönsaksjuicer.
5. Det skall inte vara obligatoriskt att ange nettoinnehållet för livsmedel
Gemenskapsbestämmelser eller, om sådana saknas, nationella bestämmelser som gäller för vissa livsmedel får i undantagsfall fastställa gränsvärden som är högre än 5 g eller 5 ml, under förutsättning att detta inte leder till att köparen får bristfällig information.
Artikel 9
2. Datumet skall föregås av orden
3. De ord som anges i punkt 2 skall följas av
Om det behövs, skall dessa uppgifter följas av de förvaringsanvisningar som man måste rätta sig efter för att varan skall hålla sig under den angivna perioden.
- med kortare hållbarhetstid än tre månader tillräckligt att ange dag och månad,
Sättet för att ange datum kan regleras närmare i enlighet med det förfarande som fastställs i artikel 20.2.
- Viner, starkviner, mousserande viner, kryddade starkviner och liknande produkter framställda av andra frukter än druvor samt drycker som faller under KN-numren 22060091, 2206 00 93 och 2206 00 99 och som har framställts av druvor eller druvmust.
- Bageri- eller konditorivaror som med hänsyn till sitt innehåll normalt konsumeras inom 24 timmar efter tillverkningen.
- Tuggummi och liknande produkter.
1. I fråga om livsmedel som från mikrobiologisk synpunkt är lättfördärvliga och som därför efter en kort period kan antas utgära en omedelbar fara för människors hälsa, skall datum för minsta hållbarhetstid ersättas med uppgift om sista förbrukningsdag.
- antingen själva datumet, eller
3. Datumet skall bestå av dag, månad och eventuellt år i denna ordning och i okodad form.
1. Bruksanvisningen till ett livsmedel skall vara utformad så att livsmedlet kan användas på ett ändamålsenligt sätt.
De gemenskapsbestämmelser som avses i denna punkt skall antas i enlighet med det förfarande som fastställs i artikel 20.2.
För andra drycker som innehåller mer än 1,2 volymprocent alkohol skall dessa bestämmelser fastställas i enlighet med det förfarande som föreskrivs i artikel 20.2.
b) Utan hinder av punkt a och utan att det påverkar tilllämpningen av gemenskapsbestämmelser om nominella mängder, är det, om färdigförpackade livsmedel är
2. De uppgifter som anges i artikel 3 och artikel 4.2 skall vara lätta att förstå och markeras på väl synlig plats på sådant sätt att de är lätta att se, klart läsbara och outplånliga.
Detta krav får utvidgas till att omfatta även de uppgifter som avses i artikel 4.2.
5. Irland, Nederländerna och Förenade kungariket får medge undantag från artikel 3.1 och punkt 3 i denna artikel när det är fråga om mjölk och mjölkprodukter i returglas.
För livsmedel som saluhålls till konsumenter eller till storkök utan att vara färdigförpackade, eller för livsmedel som förpackas på försäljningsstället på konsumentens begäran eller är färdigförpackade för direkt försäljning, skall medlemsstaterna anta närmare bestämmelser för hur de uppgifter som omfattas av artikel 3 och artikel 4.2 skall anges.
Detta direktiv skall inte inverka på bestämmelser i nationell lagstiftning, vilka i avsaknad av gemenskapsbestämmelser innebär mindre stränga krav för märkning av livsmedel som presenteras i presentförpackningar som statyetter eller souvenirer.
2. Inom sitt eget territorium får den medlemsstat där saluföringen sker i enlighet med fördragets regler föreskriva att dessa uppgifter i märkningen skall ges på ett eller flera av gemenskapens officiella språk.
I fråga om reglerna för hur uppgifter i artikel 3 och artikel 4.2 skall anges, skall medlemsstaterna inte fastställa krav som är mer detaljerade än de som framgår av artiklarna 3-13.
2. Punkt 1 gäller inte nationella icke harmoniserade bestämmelser som motiveras av att man vill
- skydda industriella och kommersiella äganderätter, uppgifter om ursprung och registrerade ursprungbeteckningar samt att förebygga illojal konkurrens.
Den skall anmäla de planerade åtgärderna och skälen för dessa till kommissionen och de andra medlemsstaterna. Kommissionen skall samråda med medlemsstaterna inom Ständiga livsmedelskommittén, inrättad genom rådets beslut 69/414/EG(6), om den anser att sådant samråd behövs eller om någon medlemsstat begär det.
Artikel 20
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
Om det visar sig nödvändigt att vidta tillfälliga åtgärder för att underlätta tillämpningen av detta direktiv, skall de antas i enlighet med det förfarande som fastställs i artikel 20.2
Varje ändring som är nödvändig för att harmonisera sådana bestämmelser med de regler som fastställs i detta direktiv skall beslutas i enlighet med det förfarande som är tilllämpligt för varje sådan bestämmelse.
Artikel 24
Detta direktiv skall gälla också för Frankrikes utomeuropeiska department.
2. Hänvisningar till det upphävda direktivet skall tolkas som hänvisningar till detta direktiv och skall läsas i enlighet med jämförelsetabellen i bilaga V.
(Text av betydelse för EES)
av följande skäl:
(3) Med hänsyn till den tekniska utvecklingen är det nödvändigt att ändra de renhetskriterier för butylhydroxianisol (BHA) som anges i direktiv 96/77/EG. Det är därför nödvändigt att anpassa detta direktiv.
(6) De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Ständiga livsmedelskommittén.
Direktiv 96/77/EG ändras på följande sätt:
Artikel 2
3) Produkter som släpps ut på marknaden eller som märks före den 31 mars 2001 och som inte uppfyller kraven i detta direktiv får saluföras till dess att lagren är tömda.
av den 16 november 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175.1 i detta,
efter att ha hört Regionkommittén,
(1) På grundval av principerna i artikel 174 i fördraget syftar Europeiska gemenskapens program för politik och åtgärder för miljön och en hållbar utveckling (femte miljöhandlingsprogrammet)(4), kompletterat genom Europaparlamentets och rådets beslut nr 2179/98/EG(5) om en översyn av programmet, särskilt till ändringar i lagstiftningen om luftföroreningar. I programmet rekommenderas att det upprättas långsiktiga mål för luftkvaliteten. Enligt artikel 174 i fördraget skall försiktighetsprincipen tillämpas när det gäller skydd av miljön och av människors hälsa.
(4) Enligt artikel 8 i direktiv 96/62/EG skall det upprättas handlingsplaner för de zoner där koncentrationen av luftförorenande ämnen överskrider gränsvärdena plus tillämpliga tillfälliga toleransmarginaler för att säkerställa att gränsvärdena uppnås inom de fastställda tidsfristerna.
(7) Ändringar som är nödvändiga för anpassning till framsteg som görs på det vetenskapliga och tekniska området får endast gälla kriterier och metoder för att bedöma koncentrationerna av bensen och koloxid eller regler för överlämnandet av information till kommissionen och får inte leda till att gränsvärdena direkt eller indirekt ändras.
(10) När emellertid gränsvärdena för bensen enligt detta direktiv är svåra att uppnå beroende på platsspecifika spridningskarakteristika eller relevanta klimatförhållanden, och om tillämpningen av åtgärderna skulle förorsaka allvarliga socio-ekonomiska problem, kan en medlemsstat be kommissionen om en tidsbegränsad förlängning för en enstaka gång under särskilda förhållanden.
(13) Information om koncentrationer av bensen och koloxid bör översändas till kommissionen som grundval för regelbundna rapporter.
Artikel 1
a) fastställa gränsvärden för koncentrationer av bensen och koloxid i luften, så att skadliga effekter på människors hälsa och på miljön i dess helhet kan undvikas, förebyggas eller minskas,
d) upprätthålla luftkvaliteten, när den är god, och i övriga fall förbättra den med hänsyn till dess halt av bensen och koloxid.
Definitionerna i artikel 2 i direktiv 96/62/EG skall tillämpas.
b) nedre utvärderingströskel: den nivå som avses i bilaga III under vilken enbart modelleringsmetoder eller objektiva skattningsmetoder kan användas för att utvärdera luftkvaliteten, i enlighet med artikel 6.4 i direktiv 96/62/EG,
Bensen
2. När det gränsvärde som anges i bilaga I är svåra att uppnå beroende på platsspecifika spridningskarakteristika eller relevanta klimatförhållanden, t.ex. låg vindhastighet och/eller förhållanden som främjar avdunstning, och om tillämpningen av åtgärderna skulle förorsaka allvarliga socio-ekonomiska problem, kan en medlemsstat be kommissionen om en tidsbegränsad förlängning. Kommissionen kan, i enlighet med det förfarande som anges i artikel 12.2 i direktiv 96/62/EG på begäran av en medlemsstat och utan att det påverkar tillämpningen av artikel 8.3 i detta direktiv, bevilja en enstaka förlängning för en period på upp till fem år om den berörda medlemsstaten
- visar att alla rimliga åtgärder har vidtagits för att sänka koncentrationerna av de berörda föroreningarna och för att begränsa det område i vilket gränsvärdet överskrids, och
Artikel 4
Den toleransmarginal som anges i bilaga II skall tillämpas i enlighet med artikel 8 i direktiv 96/62/EG.
1. De övre och nedre utvärderingströsklarna för bensen och koloxid skall vara de tröskelvärden som anges i avsnitt I i bilaga III.
3. För zoner och tätbebyggelser där uppgifter från fasta mätstationer kompletteras med uppgifter från andra källor, t.ex. utsläppsinventeringar, indikativa mätmetoder och luftkvalitetsmodellering, skall antalet fasta mätstationer som skall upprättas och den rumsliga upplösningen för övriga metoder vara tillräckliga för att göra det möjligt att fastställa koncentrationerna av luftföroreningar i enlighet med avsnitt I i bilaga IV och avsnitt I i bilaga VI.
6. Medlemsstaterna skall underrätta kommissionen om de metoder som används för den preliminära utvärderingen av luftkvaliteten enligt artikel 11.1 d i direktiv 96/62/EG senast den dag som anges i artikel 10 i detta direktiv.
Kommitté
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
Information till allmänheten
Den information som avses i andra stycket skall åtminstone innehålla uppgifter om överskridanden av gränsvärdena för koncentrationerna under de genomsnittsperioder som anges i bilagorna I och II. Den skall även omfatta en kort utvärdering med avseende på gränsvärdena och relevant information om hälsoeffekter.
Artikel 8
2. Den rapport som avses i punkt 1 skall när det gäller bensen och koloxid särskilt ta hänsyn till följande:
c) Förhållandet mellan föroreningar och möjligheter till kombinerade strategier för att uppnå gemenskapens mål i fråga om luftkvalitet och liknande mål.
3. För att upprätthålla en hög skyddsnivå för människors hälsa och för miljön skall rapporten som avses i punkt 1 vid behov kompletteras med förslag till ändringar av detta direktiv som kan inbegripa ytterligare förlängningar av tidsfristen för att uppnå gränsvärdet för bensen enligt bilaga I vilka kan komma att beviljas i enlighet med artikel 3.2.
Medlemsstaterna skall besluta om de påföljder som skall tillämpas vid överträdelser av de nationella bestämmelser som antas i enlighet med detta direktiv. Dessa påföljder skall vara effektiva, proportionella och avskräckande.
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 13 december 2002. De skall genast underrätta kommissionen om detta.
Artikel 11
av den 28 mars 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(3) I artikel 7 i direktiv 86/362/EEG och artikel 4 i direktiv 90/642/EEG föreskrivs det att nödvändiga bestämmelser skall ses över och antas, till exempel om offentliggörande i rapporter från Europeiska gemenskapen av sammanställningar av kontrollen i medlemsstaterna, och att det skall beslutas om åtgärder på gemenskapsnivån vid rapporterade överträdelser av gränsvärdena. Erfarenheterna har bekräftat att de laboratorier som gör analyser med avseende på bekämpningsmedelsrester måste uppfylla höga kvalitetskrav för att deras resultat skall vara tillförlitliga. Laboratoriernas deltagande i regelbundna kvalifikationsprövningar och tillämpning av gemensamnaa riktlinjer för kvalitetskontroll kan användas för att verifiera att de uppfyller ackrediteringskraven enligt artikel 3 i rådets direktiv 93/99/EEG av den 29 oktober 1993(4) om ytterligare åtgärder för offentlig kontroll av livsmedel.
(6) I kommissionens meddelande KOM(97) 183 om konsumenters hälsa och livsmedelssäkerhet beskrivs kontroll- och inspektionsverksamheten på livsmedels-, veterinär- och växtskyddsområdet. Denna bör innefatta kontrollen med avseende på bekämpningsmedelsrester i och på spannmål, frukt och grönsaker.
(9) En sammanfattande översikt av kontrollsystemen i alla medlemsstater krävs för att förbättra kontrollen av bekämpningsmedelsrester i gemenskapen och medverka till att den fungerar på avsett sätt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. För att fleråriga kontrollprogram skall kunna administreras effektivt får kommissionen lämna årliga bekräftelser och kompletteringar till förslag till rekommendationer. Dessa skall, i enlighet med artikel 7.2 b i direktiv 86/362/EEG och artikel 4.2 b i direktiv 90/642/EEG, överlämnas till Ständiga kommittén för växtskydd.
1. Samordna medlemsstaternas verksamhet beträffande kraven för att skapa, registrera, hantera och överföra information om kontroll och kontrollprogram, i tillämpliga fall med hjälp av riktlinjer från Ständiga kommittén för växtskydd, särskilt riktlinjerna för kvalitetskontrollförfaranden vid analys av bekämpningsmedelsrester(5) och vägledningsdokumentet till medlemsstaterna om kommissionens rekommendation om gemenskapens samordnade kontrollprogram(6).
b) utveckling av kvalitetskontrollförfaranden för analys av bekämpningsmedelsrester, i form av anvisningar från Ständiga kommittén för växtskydd, och till regelbunden översyn på expertmöten, i princip vartannat år, av tillämpningen av sådana förfaranden på de laboratorier i medlemsstaterna som utför analyser med avseende på bekämpningsmedelsrester, i syfte att säkerställa kvalitet, noggrannhet och jämförbarhet av de uppgifter som medlemsstaterna lämnar till kommissionen och övriga medlemsstater årligen och som insamlas och sammanställs av kommissionen för offentliggörande i enlighet med artikel 7.3 i direktiv 86/362/EEG och artikel 4.3 i direktiv 90/642/EEG,
Artikel 3
- namnet på mottagaren eller mottagarna av det ekonomiska stödet från gemenskapen,
- en tidsplan för slutförandet av åtgärden.
- uppfyller kraven i artikel 3 i direktiv 93/99/EEG och
Artikel 5
3. Kommissionen skall avtala om dessa besök med nationella tjänstemän inom en lämplig tidsrymd. Förutom experter från den medlemsstat som besöks får kommissionens experter vid kontrollbesöken åtföljas av en eller flera experter från en eller flera av de övriga medlemsstaterna. Under besöken skall experten eller experterna som utsetts av kommissionen från någon medlemsstat följa kommissionens administrativa föreskrifter.
6. Bestämmelserna i denna artikel skall ses över senast den 31 oktober 2001.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
om förstärkt dialog med fiskerisektorn och de grupper som berörs av den gemensamma fiskeripolitiken
med beaktande av kommissionens förslag,
(3) De europeiska branschorganisationerna bör därför få hjälp med att förbereda den rådgivande kommitténs möten i syfte att främja analyser av alla insatser inom den gemensamma fiskeripolitiken och av effekten av dess åtgärder, att stödja olika initiativ från sektorn och att om möjligt söka finna gemensamma ståndpunkter beträffande kommissionens utkast till förslag.
Artikel 1
- förklaring av syften och åtgärder som avser den gemensamma fiskeripolitiken, särskilt förslag från kommissionen, och spridande av relevant information på detta område till fiskerisektorn och andra berörda grupper under upprätthållande av regelbundna kontakter med de berörda organisationerna och grupperna.
Kommissionen kan göra de kontroller den finner vara nödvändiga för att säkerställa efterlevnaden av villkoren för och fullgörandet av de uppgifter som denna förordning ger de europeiska branschorganisationerna, vilka bistår de ombud som kommissionen utser för detta ändamål.
Rådets förordning (EG) nr 813/2000
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel(1), särskilt artikel 17.2 i denna, och
(2) Den i artikel 15 i förordning (EEG) nr 2081/92 angivna kommittén har inte avgivit ett positivt yttrande.
Bilagan till kommissionens förordning (EG) nr 1107/96 skall kompletteras med beteckningarna i bilagan till denna förordning.
Kommissionens förordning (EG) nr 1685/2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
efter att samråd har skett med den kommitté som avses i artikel 147 i fördraget, Kommittén för jordbruksstruktur och landsbygdsutveckling och Kommittén för fiskets och vattenbrukets struktur, och
(2) I artikel 2 i Europaparlamentets och rådets förordning (EG) nr 1783/1999 av den 12 juli 1999 om Europeiska regionala utvecklingsfonden(3) anges vilken typ av åtgärder som ERUF kan delta i finansieringen av.
(5) Enligt artikel 30.3 i förordning (EG) nr 1260/1999 skall nationella regler för stödberättigande utgifter tillämpas om inte kommissionen anser det nödvändigt att anta regler på gemenskapsnivå. För vissa typer av insatser eller projekt anser kommissionen att det är nödvändigt att anta gemensamma regler om stödberättigande utgifter så att en enhetlig och rättvis tillämpning av strukturfonderna kan garanteras över hela gemenskapen. När en regel om någon särskild typ av verksamhet antas, föregriper detta inte frågan enligt vilken av de ovan nämnda fonderna medfinansieringen kan ske. Antagandet av dessa regler bör i vissa fall som bör anges, inte hindra medlemsstaterna från att tillämpa strängare nationella bestämmelser. Reglerna bör vara tillämpliga på alla utgifter som uppstått mellan de tidpunkter som anges i artikel 30.2 i förordning (EG) nr 1260/1999.
(8) De åtgärder som föreskrivs i den här förordningen är förenliga med yttrandet från Kommittén för utveckling och omställning av regioner.
Reglerna i bilagan till den här förordningen skall tillämpas vid bestämmandet av om utgifter kan anses stödberättigande enligt de stödformer som definieras i artikel 9 e i förordning (EG) nr 1260/1999.
Europaparlamentets och rådets förordning (EG) nr 2038/2000
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
efter att ha hört Regionkommittén,
(1) Enligt Europaparlamentets och rådets förordning (EG) nr 2037/2000 av den 29 juni 2000 om ämnen som bryter ned ozonskiktet(3) är export av dosaerosoler till utvecklingsländer och export av läkemedelspumpar som innehåller klorfluorkarboner förbjuden. Exporten av dessa hälsovårdsprodukter som får användas på gemenskapens marknad bör dock inte begränsas.
Artikel 1
Artikel 2
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av kommissionens förslag, och
Artikel 1
a) följande strecksatser läggas till listan i punkt 1 a:
b) följande punkt införas i punkt 1:
- Vanlig valthornssnäcka (Buccinum undatum)".
"1. Produkter enligt artikel 3 skall bedömas efter vikt eller antal per kilo. Hästräkor och krabbor skall dock delas in i storlekskategorier på grundval av skalets omfång. Stora kammusslor och vanliga valthornssnäckor skall delas in i storlekskategorier på grundval av snäckans omfång."
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av rådets förordning (EEG) nr 2913/92 om inrättandet av en tullkodex för gemenskapen
med beaktande av kommissionens förslag(1),
av följande skäl:
(3) Hänsyn bör tas till rådets resolution av den 25 oktober 1996 om förenkling och rationalisering av gemenskapens tullföreskrifter och tullförfaranden(5).
(6) Förfarandena för aktiv förädling, bearbetning under tullkontroll och temporär import bör göras lättare att använda genom att reglerna på området görs flexiblare.
(9) Under vissa omständigheter bör gynnsam behandling i tullhänseende med anledning av varors beskaffenhet eller deras användning för särskilda ändamål samt differenstaxering inom ramen för förfarandet för passiv förädling även tillämpas när en tullskuld har uppkommit av andra skäl än övergång till fri omsättning.
(12) Gemenskapens ekonomiska intressen och gäldenärens rättigheter bör skyddas mot alltför utdragna rättsliga förfaranden.
(15) Förordning (EEG) nr 2913/92 bör ändras i enlighet härmed.
Förordning (EEG) nr 2913/92 ändras på följande sätt:
2. I artikel 35 skall första stycket ersättas med följande:"Om faktorer som används för att fastställa tullvärdet på varor uttrycks i en annan valuta än den som används i den medlemsstat där värderingen görs, skall den växelkurs tillämpas som vederbörligen har offentliggjorts av de på detta område behöriga myndigheterna."
4. I artikel 115 skall punkt 4 ersättas med följande:
6. Artikel 124 skall ersättas med följande:
- importvarorna omfattas av kvantitativa importrestriktioner,
- ett exportbidrag eller en exportavgift har fastställts för förädlingsprodukterna.
7. Artikel 131 skall ersättas med följande:
8. I artikel 133 e skall följande mening läggas till:"De fall där de ekonomiska villkoren skall anses vara uppfyllda får fastställas enligt kommittéförfarandet."
1. Tillämpning av förfarandet för temporär import med partiell befrielse från importtullar skall beviljas för varor som inte omfattas av de bestämmelser som fastställts enligt artikel 141 eller som omfattas av dessa bestämmelser, men inte uppfyller alla de villkor som anges i dem för beviljande av temporär import med fullständig befrielse.
11. I artikel 167 skall punkt 3 ersättas med följande:
"1. Med undantag för de frizoner som utses i enlighet med artikel 168a skall frizonernas och frilagrens gränser samt deras infarter och utfarter övervakas av tullmyndigheterna."
1. Tullmyndigheterna får utse frizoner inom vilka tullkontroller och tullformaliteter skall utföras i enlighet med tullagerförfarandet och inom vilka bestämmelserna om tullskuld skall tillämpas i enlighet med tullagerförfarandet.
14. Artikel 212a skall ersättas med följande:
15. I artikel 215 skall följande punkt läggas till:
"b) Det tullbelopp som enligt lag skall erläggas har inte bokförts på grund av ett misstag från tullmyndigheternas sida och gäldenären kunde inte rimligen ha upptäckt detta, eftersom denne för sin del handlat i god tro och följt bestämmelserna i den gällande lagstiftningen i fråga om tulldeklarationen.
Gäldenären kan åberopa god tro om han kan visa att han under den period då den berörda kommersiella verksamheten pågick visade vederbörlig aktsamhet för att förvissa sig om att samtliga villkor för förmånsbehandling var uppfyllda.
"3. Underrättelse till gäldenären får inte ske senare än tre år efter den dag då tullskulden uppkom. Denna tidsfrist upphör att löpa från det att ett överklagande enligt artikel 243 inges till och med det att överklagandeförfarandet avslutas.
"2. Det kan också enligt kommittéförfarandet fastställas i vilka fall och på vilka villkor gäldenären kan beviljas uppskov med att betala tullarna, nämligen
- när tullskulden uppkom i enlighet med artikel 203 och det finns flera gäldenärer."
De åtgärder som krävs för att genomföra denna kodex, inklusive för tillämpningen av den förordning som avses i artikel 184, med undantag av avdelning VIII och om inte annat följer av artiklarna 9 och 10 i rådets förordning (EEG) nr 2658/87(7) och av artikel 248 i denna förordning, skall antas i enlighet med det föreskrivande förfarande som avses i artikel 247a.2 och med iakttagande av gemenskapens internationella åtaganden.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 248
1. Kommissionen skall biträdas av en tullkodexkommitté (nedan kallad kommittén).
3. Kommittén skall själv anta sin arbetsordning.
Artikel 2
av den 19 december 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Enligt rådets beslut 2000/427/EG av den 19 juni 2000, i enlighet med artikel 122.2 i fördraget om införande av den gemensamma valutan i Grekland den 1 januari 2001(2), uppfyller Grekland de nödvändiga villkoren för att införa den gemensamma valutan.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från EUGFJ-kommittén.
Förordning (EG) nr 296/96 ändras på följande sätt:
Artikel 2
av den 27 december 2000
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I kommissionens förordning (EG) nr 2125/95(4), senast ändrad genom förordning (EG) nr 2493/98(5), fastställs tullkvoterna för svampkonserver från Polen, Rumänien och Bulgarien i bilagorna II, V respektive VI enligt rådets förordning (EG) nr 3066/95 av den 22 december 1995 om införande av vissa koncessioner i form av gemenskapstullkvoter för vissa jordbruksprodukter och om autonom anpassning under en övergångsperiod av vissa jordbrukskoncessioner som föreskrivs i Europaavtalen i syfte att beakta det jordbruksavtal som ingåtts inom ramen för de multilaterala handelsförhandlingarna under Uruguayrundan(6), senast ändrad genom förordning (EG) nr 2435/98(7).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Tullkvoterna för svampkonserver av Agaricus-arter enligt KN-numren 0711 90 40, 2003 10 20 och 2003 10 30, som förtecknas i bilaga I, öppnas i enlighet med de tillämpningsföreskrifter som anges i denna förordning.
om ändring av kapitel 14 i bilaga I till rådets direktiv 92/118/EEG om djurhälso- och hygienkrav för handel inom gemenskapen med produkter, som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A.I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG
(2001/7/EG)
med beaktande av rådets direktiv 92/118/EEG om djurhälso- och hygienkrav för handel inom gemenskapen med produkter, som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A.I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG(1), senast ändrat genom kommissionens beslut 1999/724/EG(2), särskilt artikel 15 i detta, och
(2) Det är nödvändigt att vid förflyttningar över gränser ta hänsyn till sjukdomssituationen i medlemsstaterna.
Artikel 1
kommer från ett område eller en anläggning där det inte finns restriktioner beträffande någon allvarlig transmissibel sjukdom
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
om fastställande av en mall för förteckningarna över de enheter som godkänts av medlemsstaterna när det gäller handeln inom gemenskapen med levande djur, sperma och embryon, samt om bestämmelser avseende överlämnande av dessa förteckningar till kommissionen
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 89/556/EEG av den 25 september 1989 om djurhälsovillkor för handel inom gemenskapen med och import från tredje land av embryon från tamdjur av nötkreatur(4), senast ändrat genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artikel 5.3 i detta,
med beaktande av rådets direktiv 91/68/EEG av den 28 januari 1991 om djurhälsovillkor för handeln med får och getter inom gemenskapen(8), senast ändrat genom beslut 94/953/EG(9), särskilt artikel 2.9 i detta, och
(2) Det är tillåtet att bedriva handel inom gemenskapen med sperma från tama arter av nötkreatur och svin från sådana centraler som godkänts av de behöriga myndigheterna i de medlemsstater där de är belägna.
(5) För att underlätta åtkomsten till uppdaterade förteckningar för gemenskapen är det nödvändigt att harmonisera såväl mallen för dessa förteckningar som det sätt på vilket de skickas.
Artikel 1
Inom ramen för Ständiga veterinärkommitténs arbete skall kommissionen underrätta medlemsstaterna om alla eventuella ändringar av ovanstående format eller av den adress till vilken filerna skall skickas.
Kommissionens beslut
[delgivet med nr K(2001) 108]
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av rådets direktiv 91/689/EEG av den 12 december 1991 om farligt avfall(3), ändrat genom direktiv 94/31/EG(4), särskilt artikel 1.4 andra strecksatsen i detta, och
(2) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som upprättats i enlighet med artikel 18 i direktiv 75/442/EEG.
Beslut 2000/532/EG ändras på följande sätt:
Avfall som klassificeras som farligt anses uppvisa en eller flera av de egenskaper som avses i bilaga 3 till direktiv 91/689/EEG och, vad beträffar H3-H8, H10(6) och H11 i denna bilaga, en eller flera av följande egenskaper:
- ett eller flera ämnen som klassificeras som giftiga vid en total koncentration >= 3 %,
- ett eller flera frätande ämnen som klassificeras som R34 vid en total koncentration >= 5 %,
- ett ämne som är känt för att vara cancerframkallande (kategori 1 eller 2) vid en koncentration >= 0,1 %,
- ett ämne som är skadligt för fortplantningen (kategori 3) och som klassificeras som R62 eller R63 vid en koncentration >= 5 %,
2. Bilagan skall ersättas med texten i bilagan till detta beslut.
Artikel 3
av den 22 februari 2001
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Provtagningsplanerna och de diagnostiska metoderna för påvisande och bekräftelse av vissa fisksjukdomar fastställs i kommissionens beslut 92/532/EEG(3), senast ändrat genom kommissionens beslut 96/240/EG(4).
(4) Gemenskapens referenslaboratorium för fisksjukdomar, som inrättades genom rådets direktiv 93/53/EEG(5), har rådfrågats.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Detta beslut riktar sig till alla medlemsstater.
om ändring av beslut 90/424/EEG om utgifter inom veterinärområdet
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
av följande skäl:
(3) Infektiös laxanemi är en ny sjukdom som första gången förekom i gemenskapen 1998 och som kan orsaka betydande förluster för laxodlingsnäringen.
(6) Bluetongue har konsekvenser på internationell nivå för förflyttning av levande djur av känsliga arter eftersom bluetongue finns upptagen på förteckning A från Internationella byrån för epizootiska sjukdomar.
(9) I beslut 90/424/EEG föreskrivs nödåtgärder som förorsakas av förekomst av bluetongue. Det krävs även ett finansiellt stöd från gemenskapen för övervakning och vissa bekämpningsåtgärder, bland annat vaccinering i högriskområden för bluetongue eller i områden där sjukdomen är endemisk.
(12) Rådets förordning (EG) nr 2792/1999 av den 17 december 1999 om föreskrifter och villkor för gemenskapens strukturstöd inom fiskerisektorn(3), särskilt artikel 15.3 g i denna, utgör den rättsliga grunden för säkerställande av finansiellt stöd när det gäller infektiös laxanemi. Bestämmelserna i avdelning III i rådets förordning (EG) nr 1260/1999 av den 21 juni 1999 om allmänna bestämmelser för strukturfonderna(4) skall därför tillämpas genom undantag från bestämmelserna i artikel 24.5, 24.6, andra meningen, 24.8 och 24.9 i beslut 90/424/EEG.
Artikel 1
Artikel 2
av den 23 juli 2001
med beaktande av rådets direktiv 91/689/EEG av den 12 december 1991 om farligt avfall(1), särskilt artikel 1.4 i detta,
(1) En gemenskapsförteckning över avfall upprättades genom kommissionens beslut 2000/532/EG av den 3 maj 2000 om ersättning av beslut 94/3/EG om en förteckning över avfall i enlighet med artikel 1 a i rådets direktiv 75/442/EEG om avfall, och rådets beslut 94/904/EG om upprättande av en förteckning över farligt avfall i enlighet med artikel 1.4 i rådets direktiv 91/689/EEG om farligt avfall(2).
(4) Beslut 2000/532/EG bör följaktligen ändras.
Artikel 1
Detta beslut skall tillämpas från och med den 1 januari 2002.
Kommissionens beslut
[delgivet med nr K(2001) 2472]
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av rådets beslut 91/666/EEG av den 11 december 1991 om att inom gemenskapen upprätta beredskapslager av vacciner mot mul- och klövsjuka(3), senast ändrat genom kommissionens beslut 2001/181/EG(4), särskilt artiklarna 7 i detta, och
(2) I bilaga I till beslut 91/666/EEG anges närmare vilka mängder och subtyper av antigener till mul- och klövsjukeviruset som skall lagras i gemenskapens beredskapslager.
(5) Genom kommissionens beslut 2000/77/EG(8), fastställs bestämmelser för inköp av ett antal mängder av mul- och klövsjukevirusantigen A Iran 96, A Iran 99, A Malaysia 97, SAT 1, SAT 2 (stammar från östra respektive södra Afrika) och SAT 3.
(8) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
Bilagan till beslut 2000/112/EG skall ersättas med bilagan till detta beslut.
Rådets rambeslut
(2001/413/RIF)
med beaktande av kommissionens initiativ(1),
(1) Bedrägerier och förfalskningar som rör andra betalningsmedel än kontanter sker ofta på internationell nivå.
(4) Eftersom målen för detta rambeslut, nämligen att säkerställa att bedrägeri och förfalskning som rör alla andra betalningsmedel än kontanter anses vara straffbara gärningar som omfattas av effektiva, proportionella och avskräckande påföljder i alla medlemsstater, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna med hänsyn till dessa brotts internationella karaktär utan därför bättre kan uppnås på gemenskapsnivå, får gemenskapen anta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i Fördraget om upprättandet av Europeiska gemenskapen. I enlighet med proportionalitetsprincipen så som den kommer till uttryck i den artikeln går detta rambeslut inte utöver vad som är nödvändigt för att uppnå de målen.
(7) Meddelandet innehåller ett utkast till gemensam åtgärd som är en del av denna övergripande strategi och utgör utgångspunkten för detta rambeslut.
(10) Avsikten med att ge straffrättsligt skydd åt i första hand betalningsinstrument med en särskild form av skydd mot efterbildning eller missbruk är att operatörerna skall uppmuntras att förse de betalningsinstrument de ger ut med detta skydd och att instrumentet därmed förses med en förebyggande faktor.
Artikel 1
a) betalningsinstrument: ett fysiskt instrument annat än lagliga betalningsmedel (legal tender) (sedlar och mynt) som genom sin särskilda karaktär, enskilt eller tillsammans med ett annat (betalnings)instrument, gör det möjligt för innehavaren eller användaren att föra över pengar eller ett penningvärde, t.ex. kreditkort, eurocheckkort, andra av finansinstitut utgivna kort, resecheckar, eurocheckar, andra checkar och växlar som är skyddade mot efterbildning eller bedräglig användning, t.ex. genom sin utformning, kod eller undertecknande,
Brott i samband med betalningsinstrument
b) Hel- eller delförfalskning av ett betalningsinstrument med syfte att använda det för bedrägeri.
Artikel 3
- att utan rätt mata in, ändra, radera, eller undertrycka datoriserade uppgifter, särskilt identifieringsuppgifter, eller
Brottslighet i samband med särskilt anpassad utrustning
- redskap, föremål, datorprogram och alla andra instrument som är särskilt avsedda för att föröva något av de brott som avses i artikel 2 b,
Deltagande, anstiftan och försök
Påföljder
Juridiska personers ansvar
- befogenhet att fatta beslut på den juridiska personens vägnar, eller
2. Utom i de fall som avses i punkt 1 skall varje medlemsstat vidta nödvändiga åtgärder för att säkerställa att en juridisk person kan ställas till ansvar när brister i övervakning eller kontroll som skall utföras av en sådan person som avses i punkt 1 har gjort det möjligt för en person, som är underställd den juridiska personen, att begå ett sådant brott som avses i artikel 2 b-d och artiklarna 3-4.
Påföljder för juridiska personer
b) tillfälligt eller permanent näringsförbud,
2. Varje medlemsstat skall vidta nödvändiga åtgärder för att säkerställa att en juridisk person som har ställts till ansvar i enlighet med artikel 7.2 kan bli föremål för effektiva, proportionella och avskräckande påföljder eller åtgärder.
1. Varje medlemsstat skall vidta nödvändiga åtgärder för att fastställa sin behörighet rörande brott enligt artiklarna 2, 3, 4 och 5 när brott har begåtts
c) till förmån för en juridisk person som har sitt säte inom medlemsstatens territorium.
- punkt 1 c.
Utlämning och åtal
2. I denna artikel skall begreppet medborgare i en medlemsstat tolkas i enlighet med en eventuell förklaring som denna stat avgivit enligt artikel 6.1 b och c i Europeiska utlämningskonventionen.
1. Medlemsstaterna skall i enlighet med tillämpliga konventioner, multilaterala eller bilaterala avtal eller arrangemang i så hög grad som möjligt bistå varandra när det gäller förfaranden som rör brott enligt detta rambeslut.
Informationsutbyte
Artikel 13
Artikel 14
2. Senast den 2 juni 2003 skall medlemsstaterna till rådets generalsekretariat och till Europeiska gemenskapernas kommission överlämna texten till de bestämmelser genom vilka de skyldigheter som åvilar dem enligt detta rambeslut överförs till nationell lag. Senast den 2 september 2003 skall rådet mot bakgrund av en rapport som upprättats på grundval av dessa upplysningar och en skriftlig rapport från kommissionen bedöma i vilken utsträckning medlemsstaterna har vidtagit nödvändiga åtgärder för att följa detta rambeslut.
Detta rambeslut träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
om ändring av rådets direktiv 85/611/EEG om samordning av lagar och andra författningar som avser företag för kollektiva investeringar i överlåtbara värdepapper (fondföretag), vad gäller fondföretags investeringar
med beaktande av kommissionens förslag(1),
av följande skäl:
(3) Den i detta direktiv angivna definitionen av överlåtbara värdepapper gäller endast för detta direktiv och påverkar inte på något sätt de definitioner som används i nationell lagstiftning i andra sammanhang, exempelvis när det gäller beskattning. Denna definition omfattar följaktligen inte aktier och andra värdepapper som motsvarar aktier och som emitteras av sådana organ som hypoteksinstitut och industri- och utvecklingsfonder, där äganderätten i praktiken inte kan överföras på annat sätt än att det emitterande organet återköper dem.
(6) Fondföretag bör tillåtas att investera sina tillgångar i andelar i andra fondföretag och/eller andra företag för kollektiva investeringar av den öppna typen som också investerar i sådana likvida, finansiella tillgångar som omnämns i detta direktiv och som tillämpar principen om riskspridning. Det är nödvändigt att fondföretag och andra företag för kollektiva investeringar som fondföretag investerar i är föremål för effektiv tillsyn.
(9) Utöver det fall då ett fondföretag investerar i banktillgodohavanden i enlighet med sina fondbestämmelser eller sin bolagsordning kan det bli nödvändigt att tillåta alla fondföretag att inneha kompletterande likvida tillgångar, som exempelvis avistakonton. Innehav av sådana kompletterande likvida tillgångar kan exempelvis vara motiverat i följande fall, nämligen för att täcka löpande eller särskilda betalningar, vid försäljningar fram till dess att man kan återinvestera i överlåtbara värdepapper, penningmarknadsinstrument och/eller andra finansiella tillgångar som avses i detta direktiv samt för den tid under vilken det är absolut nödvändigt att uppskjuta investeringen i överlåtbara värdepapper, penningmarknadsinstrument eller andra finansiella tillgångar på grund av ogynnsamma marknadsvillkor.
(12) För OTC-derivat bör ytterligare krav ställas upp för lämplighetsbedömning av motparter och instrument, likviditet och fortlöpande värdering av positionen. Syftet med sådana ytterligare krav är att säkerställa ett tillräckligt skydd för investerarna, liknande det som de erhåller vid förvärv av derivat som handlas på reglerade marknader.
(15) Företag för kollektiva investeringar som omfattas av detta direktiv bör inte användas för andra ändamål än kollektiva investeringar av medel från allmänheten, i enlighet med bestämmelserna i detta direktiv. I de fall som fastställs i detta direktiv får fondföretag ha dotterföretag endast när detta är nödvändigt för att utföra viss, i direktivet angiven verksamhet för fondföretagets räkning. Det är nödvändigt att säkerställa en effektiv tillsyn av fondföretag. Fondföretag skall därför tillåtas att etablera dotterföretag i tredje land endast i de fall och på de villkor som anges i detta direktiv. Den allmänna skyldigheten att uteslutande agera för att tillgodose andelsägarnas intressen och framför allt målet att förbättra kostnadseffektiviteten kan under inga omständigheter rättfärdiga åtgärder från fondföretagets sida som kan hindra de behöriga myndigheterna från att utöva en effektiv tillsyn.
(18) Kommissionen kan komma att överväga att föreslå kodifiering vid lämplig tidpunkt efter det att förslagen har antagits.
Direktiv 85/611/EEG ändras härigenom på följande sätt:
- aktier och andra värdepapper som motsvarar aktier (nedan kallade aktier),
med undantag för den teknik och de instrument som avses i artikel 21.
4. I artikel 19.1 b och c skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
- Följande skall läggas till: "e) andelar i fondföretag som är auktoriserade i enlighet med detta direktiv och/eller andra företag för kollektiva investeringar enligt artikel 1.2 första och andra strecksatsen, oavsett om de är belägna i en medlemsstat eller ej, förutsatt att
- verksamheten i det andra företaget för kollektiva investeringar rapporteras halvårsvis och årsvis, så att det kan ske en värdering av tillgångar och skulder, intäkter och verksamhet under rapporteringsperioden, och
g) finansiella derivat, inklusive motsvarande kontantavräknade instrument, som omsätts på en sådan reglerad marknad som avses i punkterna a, b och c, och/eller finansiella derivatinstrument som handlas direkt mellan parterna (nedan kallade OTC-derivat), förutsatt att
- OTC-derivaten är föremål för tillförlitlig och verifierbar värdering från dag till dag samt att de vid varje tidpunkt, på fondföretagets initiativ, kan säljas, lösas in eller avslutas genom en utjämnande transaktion till ett rimligt värde, och/eller
- emitterats av ett företag, vars värdepapper omsätts på de reglerade marknader som avses i punkterna a, b eller c, eller
6. I artikel 19.2 a skall orden "och penningmarknadsinstrument" läggas till efter orden "överlåtbara värdepapper".
9. Artikel 21 skall ersättas med följande: "Artikel 21
Denna verksamhet får under inga omständigheter leda till att fondföretagen avviker från sina investeringsmål såsom de fastställts i fondföretagens fondbestämmelser, bolagsordning eller prospekt.
Ett fondföretag får inom den gräns som anges i artikel 22.5 investera i finansiella derivatinstrument som ett led i sin investeringspolicy, förutsatt att exponeringen mot de underliggande tillgångarna inte sammanlagt överstiger de investeringsgränser som anges i artikel 22. När ett fondföretag investerar i indexbaserade finansiella derivatinstrument får medlemsstaterna medge att dessa investeringar sammanlagt inte behöver rymmas inom de gränser som anges i artikel 22.
10. Artikel 22 skall ersättas med följande: "Artikel 22
- 10 % av fondföretagets tillgångar när motparten är ett kreditinstitut enligt artikel 19.1 f, eller
Trots de enskilda gränser som fastställs i punkt 1, får ett fondföretag inte kombinera
4. Medlemsstaterna får höja den 5-procentsgräns som anges i punkt 1 första meningen till högst 25 % när det gäller vissa obligationer, om de är emitterade av ett kreditinstitut som har sitt säte i en medlemsstat och enligt lag omfattas av särskild offentlig tillsyn avsedd att skydda obligationsinnehavare. Särskilt skall iakttas att kapital som härrör från emissionen av sådana obligationer enligt lag måste investeras i tillgångar som, under obligationernas hela giltighetstid kan täcka de med obligationerna förenade fordringarna och som i händelse av emittentens oförmåga att fullgöra sina ekonomiska åtaganden skall med prioritet användas för återbetalning av kapital och upplupen ränta.
5. Vid beräkningen av den gräns på 40 % som anges i punkt 2 skall inte de överlåtbara värdepapper och penningmarknadsinstrument som anges i punkterna 3 och 4 beaktas.
Medlemsstaterna kan tillåta investeringar upp till en gräns på 20 % i överlåtbara värdepapper och penningmarknadsinstrument inom samma grupp."
- Det skall ha en tillräckligt diversifierad sammansättning.
2. Medlemsstaterna får höja den gräns som fastställs i punkt 1 till högst 35 % när det visar sig motiverat på grund av exceptionella marknadsvillkor särskilt på reglerade marknader där vissa överlåtbara värdepapper eller penningmarknadsinstrument i hög grad dominerar. Investeringar upp till denna gräns är bara tillåtna för en enda emittent."
1. Ett fondföretag får förvärva andelar i fondföretag och/eller andra företag för kollektiva investeringar enligt artikel 19.1 e, under förutsättning att inte mer än 10 % av dess tillgångar investeras i andelar i ett enda fondföretag eller annat företag för kollektiva investeringar. Medlemsstaterna får höja denna gräns till högst 20 %.
3. När ett fondföretag investerar i andelar i andra fondföretag och/eller andra företag för kollektiva investeringar som direkt eller genom delegering förvaltas av samma förvaltningsbolag eller av ett annat bolag till vilket förvaltningsbolaget är anknutet via gemensam företagsledning eller ägarkontroll eller genom ett betydande direkt eller indirekt ägande får detta förvaltningsbolag eller det andra bolaget inte debitera några avgifter för teckning eller inlösen av fondföretagets investeringar i andelar i dessa andra fondföretag och/eller företag för kollektiva investeringar.
1. I prospektet skall anges vilka kategorier av tillgångar i vilka fondföretaget har tillstånd att investera. Det skall anges om transaktioner med finansiella derivatinstrument är tillåtna; i så fall måste det finnas en tydlig uppgift om huruvida dessa får utföras i syfte att säkra tillgångar eller i avsikt att nå investeringsmål och hur det möjliga resultatet av användningen av finansiella derivatinstrument kan påverka riskprofilen.
4. På begäran av en investerare måste förvaltningsbolaget också tillhandahålla kompletterande information om de kvantitativa gränser som gäller för fondföretagets riskhantering, de metoder som har valts för denna och den senaste utvecklingen av riskerna med och avkastningen från de viktigaste instrumentkategorierna."
2. Följande strecksats skall läggas till: "- 10 % av de penningmarknadsinstrument som emitterats av ett och samma organ."
18. Artikel 25.3 e skall ersättas med följande: "e) Ett eller flera investeringsbolags aktieinnehav i dotterbolag vars verksamhet enbart består i förvaltning, rådgivning eller saluföring i det land där dotterbolaget är beläget, vid återköp av andelar på begäran av andelsägarna, uteslutande för investeringsbolagets eller investeringsbolagens räkning."
20. Artikel 41.2 skall ersättas med följande: "2. Bestämmelserna i punkt 1 skall inte hindra sådana företag från att förvärva överlåtbara värdepapper, penningmarknadsinstrument eller andra finansiella instrument som avses i artikel 19.1 e, g och h och som inte är till fullo betalda."
- Förtydligande av definitionerna för att säkerställa en enhetlig tillämpning av detta direktiv inom hela gemenskapen.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
1. Senast den 13 februari 2005 skall kommissionen lägga fram en rapport för rådet och Europaparlamentet om tillämpningen av det ändrade direktiv 85/611/EEG tillsammans med eventuella förslag till ändringar. Rapporten skall särskilt innehålla
c) en utvärdering av hur fonderna organiseras, inklusive bestämmelser och metoder för delegering samt förhållandet mellan fondförvaltare och förvaringsinstitut,
När kommissionen utarbetar denna rapport skall den i största möjliga utsträckning samråda med de olika branschintressena samt med konsumentorganisationer och tillsynsorgan.
Medlemsstaterna skall anta de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 13 augusti 2003. De skall genast underrätta kommissionen om detta.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
om tillämpningen av artiklarna 87 och 88 i EG-fördraget på statligt stöd till små och medelstora företag
med beaktande av rådets förordning (EG) nr 994/98 av den 7 maj 1998 om tillämpningen av artiklarna 92 och 93 i Fördraget om upprättandet av Europeiska gemenskapen på vissa slag av övergripande statligt stöd(1), särskilt artikel 1 a i och 1 b i denna,
av följande skäl:
(3) Kommissionen har i ett stort antal beslut tillämpat artiklarna 87 och 88 i fördraget på små och medelstora företag både inom och utanför stödområden och har också redogjort för sin politik på området, senast i gemenskapens riktlinjer för statligt stöd till små och medelstora företag(3), och i riktlinjerna för statligt stöd för regionala ändamål(4). För att säkerställa effektiv kontroll och förenklad administration utan att kommissionens kontroll försvagas bör kommissionen, mot bakgrund av dels sin stora erfarenhet av att tillämpa dessa artiklar på små och medelstora företag, dels de allmänna texter om små och medelstora företag och regionalstöd som den antagit på grundval av dessa artiklar, göra bruk av sina befogenheter enligt förordning (EG) nr 994/98.
(6) Genom denna förordning bör undantag medges för alla stöd som uppfyller förordningens samtliga tillämpliga krav, och för alla stödordningar, förutsatt att varje stöd som kan beviljas inom ramen för dessa ordningar uppfyller samtliga tillämpliga krav enligt förordningen. För att säkerställa effektiv kontroll och förenklad administration utan att kommissionens kontroll försvagas bör stödordningar och enskilda stöd som inte omfattas av någon stödordning innehålla en uttrycklig hänvisning till denna förordning.
(9) För att bättre säkerställa att stödet är proportionellt och begränsas till det belopp som är nödvändigt, bör tröskelvärdena i enlighet med kommissionens fastlagda praxis uttryckas som stödnivåer i förhållande till stödberättigande kostnader snarare än som maximala stödbelopp.
(12) Enligt kommissionens erfarenhet bör stödtaken fastställas till en nivå som ger en balans mellan målsättningen att skapa minsta möjliga snedvridning av konkurrensen inom den understödda sektorn och målsättningen att underlätta de små och medelstora företagens ekonomiska utveckling.
(15) För att inte gynna kapitalfaktorn på bekostnad av arbetsfaktorn i samband med en investering, bör i denna förordning föreskrivas en möjlighet att mäta investeringsstöd på grundval av antingen investeringskostnader eller kostnader för nyanställningar i samband med att ett investeringsprojekt genomförs.
(18) För att säkerställa att stödet är nödvändigt och fungerar som ett incitament för att utveckla en viss verksamhet bör undantag enligt denna förordning inte beviljas för verksamhet som stödmottagaren även skulle bedriva på rena marknadsvillkor.
(21) Med hänsyn till kommissionens erfarenhet på detta område, särskilt av hur ofta det i allmänhet är nödvändigt att se över politiken på området för statligt stöd, bör tillämpningsperioden för denna förordning begränsas. Om denna förordnings giltighetstid skulle löpa ut utan att förlängas, bör stödordningar som redan undantagits enligt denna förordning fortsätta att vara undantagna i sex månader.
Tillämpningsområde
a) verksamheter i samband med produktion, bearbetning eller marknadsföring av de produkter som förtecknas i bilaga I till fördraget,
Artikel 2
a) stöd: varje åtgärd som uppfyller samtliga kriterier som anges i artikel 87.1 i fördraget.
d) investering i immateriella tillgångar: investering i överföring av teknik genom förvärv av patenträttigheter, licenser, know-how eller icke patentskyddad teknisk kunskap.
g) antal anställda: antalet arbetskraftsenheter per år, dvs. antalet heltidsanställda under ett år, medan deltidsarbete eller säsongsarbete utgör delar av arbetskraftsenheter.
1. Enskilda stöd som inte omfattas av någon stödordning och som uppfyller samtliga villkor enligt denna förordning skall anses vara förenliga med den gemensamma marknaden enligt artikel 87.3 i fördraget och skall undantas från anmälningskravet enligt artikel 88.3 i fördraget, under förutsättning att stöden innehåller en uttrycklig hänvisning till denna förordning, med angivande av förordningens titel och en hänvisning till dess offentliggörande i Europeiska gemenskapernas officiella tidning.
b) stödordningen innehåller en uttrycklig hänvisning till denna förordning, med angivande av förordningens titel och en hänvisning till dess offentliggörande i Europeiska gemenskapernas officiella tidning.
Investeringar
a) 15 % för små företag, eller
a) 10 procentenheter brutto i de områden som omfattas av artikel 87.3 c, under förutsättning att den totala stödnivån netto inte överstiger 30 %, eller
4. De tak som fastställs i punkterna 2 och 3 skall gälla stödnivån beräknad antingen som en procentandel av investeringens stödberättigande kostnader eller som en procentandel av lönekostnaden för den sysselsättning som skapas till följd av investeringen (stöd till skapande av arbetstillfällen) eller en kombination av båda, under förutsättning att stödet inte överstiger det högsta belopp som endera av beräkningssätten resulterar i.
a) Den skapade sysselsättningen måste ha samband med genomförandet av ett investeringsprojekt i materiella eller immateriella tillgångar. Arbetstillfällena måste skapas inom tre år från det att investeringen har slutförts.
Artikel 5
a) För tjänster som tillhandahålls av utomstående konsulter får stödet brutto inte överstiga 50 % av kostnaderna för dessa tjänster. De berörda tjänsterna får varken vara av fortlöpande eller periodiskt slag eller röra företagets ordinarie driftsutgifter, som t.ex. rutinmässig skatterådgivning, regelbunden juridisk rådgivning eller annonskostnader.
Beviljande av stora enskilda stöd
i) stödnivån brutto i områden som inte är berättigade till regionalstöd är minst 50 % av de stödnivåer som anges i artikel 4.2,
Artikel 7
- har fått en ansökan om stöd från stödmottagaren, eller
Kumulering
Artikel 9
2. Medlemsstaterna skall föra detaljerade register över de stödordningar som undantas genom denna förordning, de enskilda stöd som beviljas enligt dessa stödordningar, och de enskilda stöd som undantas enligt denna förordning och som beviljas vid sidan om en befintlig stödordning. Dessa register skall innehålla alla uppgifter som behövs för att det skall vara möjligt att fastställa att de villkor för beviljande av undantag som anges i denna förordning har uppfyllts inbegripet uppgifter om företagets status som litet eller medelstort företag. Medlemsstaterna skall bevara ett register över ett enskilt stöd under tio år från den dag då stödet beviljades, och, när det gäller en stödordning, under tio år från den dag då det sista enskilda stödet beviljades enligt stödordningen. En berörd medlemsstat skall på skriftlig begäran inom tjugo arbetsdagar, eller inom en längre tidsfrist som anges i begäran, förse kommissionen med alla uppgifter den anser sig behöva för att kunna bedöma om villkoren i denna förordning har följts.
Ikraftträdande och giltighetstid
av den 9 februari 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Genom kommissionens förordning (EG) nr 2734/2000 av den 14 december 2000 om ändring av förordning (EEG) nr 1627/89 om uppköp av nötkött genom anbudsinfordran och om undantag från eller ändring av förordning (EG) nr 562/2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 1254/1999 vad avser systemen för offentliga interventionsuppköp inom nötköttssektorn(2), ändrad genom förordning (EG) nr 3/2001(3), fastställdes ett antal ändringar av eller undantag från kommissionens förordning (EG) nr 562/2000(4) med anledning av den exceptionella situationen på marknaden till följd av den senaste händelseutvecklingen i samband med bovin spongiform encefalopati (BSE).
(4) Med hänsyn till att produkter som köps upp för intervention även får säljas efter den 1 januari 2002, när det obligatoriska märkningssystemet enligt Europaparlamentets och rådets förordning av den 17 juli 2000 om upprättande av ett system för identifiering och registrering av nötkreatur samt märkning av nötkött och nötköttsprodukter och om upphävande av rådets förordning (EG) nr 820/97(5) skall börja tillämpas, bör det för avtal som sluts från och med den 12 februari, dvs. från och med februari månads första anbudsförfarande, vara obligatoriskt att i märkningen ange det eller de länder där de berörda djuren är födda eller har fötts upp enligt artikel 13.5 i förordning (EG) nr 1760/2000, och i förekommande fall de uppgifter som föreskrivs i artikel 2.2 i kommissionens förordning 1825/2000 om tillämpningsföreskrifter för Europaparlamentets och rådets förordning (EG) nr 1760/2000(6).
(7) Med hänsyn till händelseutvecklingen bör denna förordning träda i kraft omedelbart.
Artikel 1
- skall ingen begränsning av den maximala vikten för slaktkroppar tillämpas för de två anbudsförfarandena i februari månad.
Förordning (EG) nr 562/2000 ändras på följande sätt:
2. I bilaga III skall punkt 2 b ersättas med följande:
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
om ändring av bilaga II till rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I enlighet med förordning (EEG) nr 2377/90 måste gränsvärden för högsta tillåtna restmängder successivt fastställas för samtliga farmakologiskt verksamma substanser som används inom gemenskapen veterinärmedicinska läkemedel som är avsedda att ges till livsmedelsproducerande djur.
(4) För kontroll av resthalter bör enligt tillämplig gemenskapslagstiftning gränsvärden vanligtvis fastställas för målvävnaderna lever eller njure. I den internationella handeln avlägsnas dock ofta lever och njure från slaktkroppen, och gränsvärden bör därför alltid fastställas även för muskel- eller fettvävnader.
(7) En tillräckligt lång tidsfrist bör fastställas innan denna förordning träder i kraft så att medlemsstaterna kan göra de nödvändiga anpassningarna till bestämmelserna i denna förordning av tillstånden att släppa ut de berörda veterinärmedicinska läkemedlen på marknaden, vilka beviljats enligt rådets direktiv 81/851/EEG(3), senast ändrat genom kommissionens direktiv 2000/37/EG(4).
Artikel 1
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om tillämpningsföreskrifter till rådets förordning (EG) nr 104/2000 beträffande beviljande av schablonmässigt stöd för vissa fiskeriprodukter
med beaktande av rådets förordning (EG) nr 104/2000 av den 17 december 1999 om den gemensamma organisationen av marknaden för fiskeri- och vattenbruksprodukter(1), särskilt artikel 24.8 i denna, och
(2) I syfte att harmonisera och förenkla bör de förfaranden som krävs inom ramen för det schablonmässiga stödet vara analoga med dem som gäller för den ekonomiska ersättningen och förädlingsstödet, såsom följer av kommissionens förordning (EG) nr 2509/2000 av den 15 november 2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 104/2000 beträffande beviljande av ekonomisk ersättning för återtag från marknaden av vissa fiskeriprodukter(3), och kommissionens förordning (EG) nr 2814/2000 av den 21 december 2000 om tillämpningsföreskrifter till rådets förordning (EG) nr 104/2000 beträffande beviljande av förädlingsstöd för vissa fiskeriprodukter(4). Villkoren för att bevilja schablonmässigt stöd bör följaktligen fastställas på denna grund och kommissionens förordning (EG) nr 4176/88 av den 28 december 1988 om tillämpningsföreskrifter för beviljande av fast stöd för vissa fiskeri- och vattenbruksprodukter(5), senast ändrad genom förordning (EG) nr 3516/93(6), bör upphöra att gälla.
(5) Det schablonmässiga stödet får betalas ut först efter fiskeårets slut. Det bör emellertid införas en möjlighet att bevilja förskott, förutsatt att säkerhet ställs.
(8) Stödmottagarna bör föra lagerbokföring (i kg) över de varor som varje månad bjuds ut till försäljning, återtas och förädlas för att effektiviteten i kontrollerna skall kunna ökas och de bör meddela dessa uppgifter till medlemsstaten. För ett väl fungerande system är det tillräckligt att kräva lagerbokföring under den kortast tillåtna lagringsperioden.
KAPITEL I
Artikel 2
Villkor för att bevilja schablonmässigt stöd enligt artikel 24.2 i förordning (EG) nr 104/2000 (nedan kallat schablonersättning)
Artikel 4
KAPITEL III
1. Schablonbidraget skall fastställas innan fiskeåret börjar enligt artikel 38.2 i förordning (EG) nr 104/2000. Beloppet skall fastställas per viktenhet och gälla för nettovikten av de produkter som anges i bilaga IV till förordning (EG) nr 104/2000.
a) Kostnader för energi.
d) Beredningskostnader (ingredienser).
5. Det schablonbidrag som fastställs för ett fiskeår skall gälla för produkter som började lagras under det året, oavsett när lagringen upphör.
Artikel 7
Slutbestämmelser
2. Efter ansökan av en berörd producentorganisation skall förskott beviljas varje månad för återtagna eller förädlade kvantiteter, under förutsättning att producentorganisationen ställer en säkerhet som minst motsvarar 105 % av förskottsbeloppet.
Artikel 9
3. Producentorganisationen skall i fråga om de produkter som återtagits eller förädlats varje månad underrätta medlemsstaten om datum, art och kvantitet.
Artikel 11
Europaparlamentets och rådets förordning (EG) nr 999/2001
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) Denna förordning har direkt avseende på folkhälsan och har betydelse för hur den inre marknaden fungerar. Den omfattar produkter som ingår i bilaga I till fördraget men även produkter som inte ingår i denna bilaga. Det är därför lämpligt att välja artikel 152.4 b i fördraget som rättslig grund.
(6) Det bör införas bestämmelser om att kommissionen får vidta skyddsåtgärder om den behöriga myndigheten i en medlemsstat eller i ett tredje land inte har hanterat TSE-risken på lämpligt sätt.
(9) Medlemsstaterna måste årligen genomföra ett övervakningsprogram för BSE och scrapie och meddela kommissionen och de övriga medlemsstaterna resultaten härav samt om någon annan form av TSE har uppträtt.
(12) Det bör föreskrivas att varje misstanke om någon form av TSE hos något djur skall anmälas till den behöriga myndigheten, som omedelbart skall vidta alla lämpliga åtgärder, och i synnerhet fastställa restriktioner för förflyttning av det misstänkta djuret i väntan på resultatet av undersökningen eller låta slakta det under officiell övervakning. Om den behöriga myndigheten inte kan utesluta möjligheten att djuret är smittat med TSE, bör den se till att lämpliga undersökningar görs och hålla slaktkroppen under officiell övervakning till dess att en diagnos har ställts.
(15) Det bör fastställas bestämmelser om avyttring av vissa levande djur och animaliska produkter. I nuvarande gemenskapslagstiftning om identifiering och registrering av nötkreatur finns bestämmelser om ett system som gör det möjligt att, enligt internationella normer, spåra djuren tillbaka till moderdjuret och ursprungsbesättningen. Det bör införas bestämmelser om likvärdiga garantier i fråga om nötkreatur som importeras från tredje land. Djur och animaliska produkter som omfattas av nämnda lagstiftning och som förflyttas vid handel inom gemenskapen eller importeras från tredje land bör åtföljas av de intyg som krävs enligt gemenskapslagstiftningen, vid behov kompletterade i enlighet med denna förordning.
(18) Det är nödvändigt att genomföra gemenskapsinspektioner i medlemsstaterna för att garantera en enhetlig tillämpning av kraven när det gäller förebyggande, kontroll och utrotning av TSE samt även föreskriva tillämpning av kontrollförfaranden. För att säkerställa att de garantier som lämnas av tredje land vid import av levande djur och animaliska produkter till gemenskapen är likvärdiga med dem som är i kraft inom gemenskapen bör gemenskapsinspektioner och -kontroller genomföras på plats för att kontrollera att importvillkoren uppfylls av exporterande tredje land.
(21) De övergångsåtgärder som är nödvändiga för att i synnerhet reglera användningen av de typer av riskmaterial som anges i denna förordning bör fastställas.
(24) Eftersom tillämpningsföreskrifterna för denna förordning är åtgärder med allmän räckvidd enligt artikel 2 i rådets beslut 1999/468/EG, bör de antas enligt det föreskrivande förfarandet i artikel 5 i det beslutet.
ALLMÄNNA BESTÄMMELSER
1. I denna förordning fastställs bestämmelser för förebyggande, kontroll och utrotning av transmissibel spongiform encefalopati (TSE) hos djur. Den skall tillämpas på framställning och avyttring, samt i vissa särskilda fall export, av levande djur och animaliska produkter.
b) produkter, eller utgångsmaterial och mellanprodukter till dessa, som inte är avsedda att användas i livsmedel, foder eller gödningsmedel,
Artikel 2
Tillämpningsföreskrifter för denna artikel skall fastställas enligt det förfarande som avses i artikel 24.2.
1. I denna förordning används följande beteckningar med de betydelser som här anges:
c) animaliska produkter: alla produkter som härrör från eller innehåller en produkt som härrör från något av de djur som omfattas av bestämmelserna i direktiv 89/662/EEG(5) eller direktiv 90/425/EEG(6).
f) kategori: någon av de klassificeringskategorier som avses i kapitel C i bilaga II.
i) anläggning: varje anläggning eller plats där djur som omfattas av denna förordning hålls, föds upp och hanteras eller visas upp för allmänheten.
l) snabbtest: de analysmetoder som avses i kapitel C.4 i bilaga X och som ger ett resultat inom 24 timmar.
3. Om en term i denna förordning inte har definierats i punkt 1 eller i bilaga I, skall de relevanta definitionerna i förordning (EG) nr 1760/2000(7) och de definitioner som finns i eller som har fastställts med stöd av direktiven 64/432/EEG(8), 89/662/EEG, 90/425/EEG och 91/68/EEG(9) tillämpas i den utsträckning som det hänvisas till dem i denna text.
1. När det gäller genomförandet av skyddsåtgärder skall principerna och bestämmelserna i artikel 9 i direktiv 89/662/EEG, artikel 10 i direktiv 90/425/EEG, artikel 18 i direktiv 91/496/EEG(10) och artikel 22 i direktiv 97/78/EG(11) tillämpas.
FASTSTÄLLANDE AV BSE-STATUS
1. BSE-status för en medlemsstat, ett tredje land eller en region i en medlemsstat eller ett tredje land (nedan kallade länder eller regioner), kan endast fastställas på grundval av kriterierna i kapitel A i bilaga II och resultaten av en riskanalys som identifierar samtliga potentiella faktorer för uppkomsten av BSE, angivna i kapitel B i bilaga II, samt deras utveckling över tiden.
Detta beslut skall antas inom sex månader efter det att ansökan samt de relevanta upplysningar som avses i punkt 1, andra stycket, har lämnats in. Om kommissionen finner att underlaget inte innehåller den information som fastställs i kapitlen A och B i bilaga II, skall den begära ytterligare information inom en tidsfrist som skall fastställas. Det slutliga beslutet skall sedan fattas inom sex månader efter det att den fullständiga informationen lämnats.
Denna analys skall innehålla en avgörande statistisk undersökning av den epidemiologiska situationen avseende TSE i den ansökande medlemsstaten eller det ansökande tredje landet, vilken skall genomföras med snabbtest med hjälp av ett screeningförfarande. Kommissionen skall beakta de klassificeringskriterier som Internationella byrån för epizootiska sjukdomar har fastställt.
Den berörda medlemsstaten eller det berörda tredje landet skall stå för kostnaderna för detta förfarande.
6. Bibehållandet av ett tredje land i någon av förteckningarna enligt gemenskapens bestämmelser om tillstånd att till Europeiska gemenskapen exportera levande djur och animaliska produkter, för vilka det finns särskilda bestämmelser i denna förordning, beslutas enligt det förfarande som anges i artikel 24.2 och under förutsättning att, med hänsyn till tillgänglig information eller om TSE förmodas förekomma - den information som föreskrivs i punkt 1 lämnas. Om sådan information inte lämnas inom tre månader från det att kommissionen begärt den, skall bestämmelserna i punkt 4 i denna artikel tillämpas så länge informationen inte har lämnats och inte har kunnat utvärderas i enlighet med punkt 2 eller punkt 3.
8. De beslut som avses i punkterna 2, 3, 4, 6 och 7 skall grundas på en riskbedömning med hänsyn till de rekommenderade kriterier som fastställs i kapitlen A och B i bilaga II.
Artikel 6
Snabbtest skall godkännas för detta ändamål enligt det förfarande som avses i artikel 24.2 och införas i en förteckning i kapitel C.4 i bilaga X.
4. Medlemsstaterna skall förelägga kommissionen en årlig rapport som skall innehålla åtminstone den information som avses i kapitel B.I i bilaga III. Rapporten för varje kalenderår skall överlämnas senast den 31 mars nästkommande år. Inom tre månader efter det att de nationella rapporterna har mottagits, skall kommissionen för Ständiga veterinärkommittén lägga fram en sammanfattning av dessa rapporter, som skall innehålla åtminstone den information som avses i kapitel B.II i bilaga III.
1. Det är förbjudet att utfodra idisslare med protein som härrör från däggdjur.
4. De medlemsstater eller regioner i medlemsstaterna som har placerats i kategori 5 skall inte tillåtas att exportera eller lagra sådant foder för livsmedelsproducerande djur som innehåller protein som härrör från däggdjur, eller foder som är avsett för däggdjur, med undantag av hundar och katter, och som innehåller bearbetat protein som härrör från däggdjur.
Artikel 8
Dessa specificerade riskmaterial eller bearbetade material av dessa får endast avyttras eller, i förekommande fall, exporteras för slutlig destruktion i enlighet med punkterna 3 och 4 eller i förekommande fall punkt 7 c eller punkt 8 i bilaga V. De får inte importeras till gemenskapen. Transitering genom gemenskapens territorium skall ske i överensstämmelse med kraven i artikel 3 i direktiv 91/496/EEG.
3. I de medlemsstater eller regioner inom dessa som har placerats i kategorierna 2, 3, 4 och 5 enligt kapitel C i bilaga II får laceration, efter bedövning, av vävnad från centrala nervsystemet med ett avlångt, stavformigt instrument som förs in i hjärnskålen inte användas för nötkreatur, får eller getter vars kött är avsett som livsmedel eller foder.
Trots vad som sägs i artiklarna 1-4, kan efter samråd med den behöriga vetenskapliga kommittén och på grundval av en bedömning av risken för förekomst eller spridning av sjukdomen eller för att människor utsätts för smitta, ett beslut likaså fattas i enlighet med det förfarande som avses i artikel 24.2 om att tillåta att kotpelare och dorsala rotganglier från nötkreatur i eller från de länder eller regioner som placerats i kategori 5, används i livsmedel, foder och gödningsämnen.
Animaliska produkter som härrör från eller innehåller material från idisslare
3. Bestämmelserna i punkterna 1 och 2 skall, när det gäller kriterierna i punkt 5 i bilaga V, inte tillämpas på idisslare som har genomgått ett alternativt test som godkänts enligt det förfarande som avses i artikel 24.2 och där testresultaten är negativa.
Utbildningsprogram
KAPITEL IV
Anmälan
Den behöriga myndigheten skall utan dröjsmål vidta de åtgärder som fastställs i artikel 12 i denna förordning, liksom alla andra nödvändiga åtgärder.
1. Alla djur som misstänks vara smittade med TSE skall vara föremål för officiella restriktioner vad avser förflyttning i avvaktan på att resultaten av den behöriga myndighetens kliniska och epidemiologiska undersökning blir tillgängliga, eller avlivas för laboratorieundersökning under officiell kontroll.
Om det kan styrkas att den anläggning där djuret befann sig när man misstänkte BSE förmodligen inte är den anläggning där djuret kan ha exponerats för BSE, får den behöriga myndigheten besluta att bara det djur som misstänks vara smittat skall vara föremål för en officiell restriktion vad avser förflyttning. Om den behöriga myndigheten anser det nödvändigt, får den också besluta att övriga anläggningar eller endast den anläggning där exponeringen förekom skall ställas under officiell övervakning, beroende på den tillgängliga epidemiologiska informationen.
3. Alla delar av det misstänkta djurets kropp, inklusive huden, skall hållas under officiell övervakning till dess en negativ diagnos har ställts, eller destrueras i enlighet med punkt 3 eller 4 i bilaga V.
Åtgärder vid bekräftad förekomst av TSE
b) En undersökning skall genomföras för att identifiera alla riskdjur i enlighet med punkt 1 i bilaga VII.
2. I avvaktan på att de åtgärder som avses i punkterna 1 b och 1 c genomförs, skall den anläggning där djuret befann sig när förekomsten av TSE bekräftades ställas under officiell övervakning och all förflyttning från eller till anläggningen av djur som riskerar att ha smittats med TSE samt av animaliska produkter från dessa djur godkännas av den behöriga myndigheten, så att djuren och de berörda animaliska produkterna omedelbart skall kunna spåras och identifieras.
4. Ägarna skall utan dröjsmål ersättas för förlusten av de djur som har avlivats och de animaliska produkter som har destruerats i enlighet med artikel 12.2 och punkterna 1 a och 1 c i denna artikel.
Artikel 14
2. Om det är nödvändigt för att möjliggöra en enhetlig tillämpning av gemenskapslagstiftningen får riktlinjerna harmoniseras enligt det förfarande som avses i artikel 24.2.
Artikel 15
2. Avyttring av den första generationen avkomma, sperma, embryon och ägg från djur som misstänks eller bekräftats vara smittade med TSE skall omfattas av de villkor som anges i kapitel B i bilaga VIII.
Avyttring av animaliska produkter
b) i) Rå mjölk enligt definitionen i direktiv 92/46/EEG(13).
iv) Dikalciumfosfat (utan spår av protein eller fett).
vii) Kollagen som härrör från hudar och skinn enligt punkt v.
a) djur som är födda efter den dag då förbudet mot utfodring av idisslare med bearbetat protein som härrör från däggdjur började gälla,
4. Om ett djur förflyttas från ett land eller en region till ett annat land eller en annan region placerade i en annan kategori, skall det klassificeras i den högsta kategorin för de länder eller regioner där det har vistats mer än ett dygn, såvida inte tillräckliga garantier om att djuret inte har utfodrats med foder från detta land eller denna region som klassificerats i den högsta kategorin kan lämnas.
7. Enligt det förfarande som avses i artikel 24.2 får bestämmelserna i punkterna 1-6 utvidgas till att omfatta andra animaliska produkter. Tillämpningsföreskrifter för denna artikel skall fastställas enligt samma förfarande.
Lämpliga handelsdokument för handel med animaliska produkter skall i förekommande fall kompletteras med en uppgift om den kategori som kommissionen i enlighet med artikel 5 placerat medlemsstaten eller ursprungsregionen i.
KAPITEL VI
Referenslaboratorier
Artikel 20
2. När så krävs för att möjliggöra en enhetlig tillämpning av denna artikel, skall tillämpningsföreskrifter - inbegripet metoden för att bekräfta förekomst av BSE hos får och getter - fastställas enligt det förfarande som avses i artikel 24.2.
1. Experter från kommissionen får, när så krävs för en enhetlig tillämpning av denna förordning, i samarbete med de behöriga myndigheterna i medlemsstaterna genomföra kontroller på plats. Den medlemsstat på vars territorium en kontroll utförs skall ge all nödvändig hjälp till experterna så att de kan fullgöra sina uppgifter. Kommissionen skall underrätta den behöriga myndigheten om resultaten av de utförda kontrollerna.
KAPITEL VII
Övergångsbestämmelser för specificerat riskmaterial
3. Detaljerade bestämmelser om denna statistiska undersökning skall, efter samråd med den relevanta vetenskapliga kommittén, antas enligt det förfarande som avses i artikel 24.2.
Ändring av bilagorna och övergångsbestämmelser
Artikel 24
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 25
Artikel 26
Kommissionens förordning (EG) nr 1282/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) För att underlätta förvaltningen av marknaden för vin måste ett datum anges då deklarationerna skall göras. Eftersom skörden äger rum vid olika tidpunkter i de olika medlemsstaterna bör tidsfristerna för inlämning av producenternas deklarationer spridas över en lämplig period. Även de aktörer som levererar vinprodukter före de angivna deklarationsdatumen bör åläggas att lämna deklarationer.
(6) Kategorin "annat vin" bör definieras i förhållande till den klassificering av druvsorter som får odlas inom gemenskapen som fastställs i artikel 19 i förordning (EG) nr 1493/1999.
(9) Tillräcklig information om produktion och lager inom vinsektorn återfinns för närvarande bara i de skörde- och lagerdeklarationer som lämnas av de berörda parterna. Lämpliga åtgärder bör därför vidtas för att säkerställa att dessa deklarationer lämnas av vederbörande och att de är fullständiga och korrekta. Det bör ges möjlighet till påföljder för den händelse att deklarationer inte lämnas eller är felaktiga eller ofullständiga. För att förenkla behandlingen av deklarationsuppgifterna bör varje deklaration som lämnas in i den behöriga administrativa enheten anses vara oberoende av andra deklarationer som samma producent kan ha lämnat in till andra av medlemsstatens administrativa enheter.
(12) I detta sammanhang är det lämpligt att erinra om att det är nödvändigt att respektera de tidsfrister som fastställs för överföring av uppgifterna för att säkerställa marknadsuppföljningen och se till att effektiva åtgärder inom ramen för budgeten kan vidtas i rätt tid.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
2. Följande personer behöver emellertid inte lämna in någon skördedeklaration:
c) Skördare vars jordbruksföretag omfattar mindre än 10 ar vinodlingsareal och som levererar hela skörden till ett vinkooperativ eller en sammanslutning som de tillhör eller är associerade med. I sådana fall skall skördarna till jordbrukskooperativen eller sammanslutningarna lämna deklarationer med uppgift om
iii) den berörda vinodlingens areal och läge.
a) Skördare som själva bearbetar hela sin druvskörd till vin eller som låter bearbeta den för egen räkning.
Artikel 4
3. De skördare som avses i artikel 2.2 samt de producenter som i egna anläggningar av inköpta produkter framställer mindre än tio hektoliter vin, som varken har saluförts eller kommer att saluföras i någon form, är inte skyldiga att lämna någon produktions-, eller i förekommande fall behandlings- eller saluföringsdeklaration.
Artikel 5
Artikel 6
2. I punkt 1 avses med detaljister fysiska eller juridiska personer eller sammanslutningar av sådana personer vars affärsverksamhet omfattar försäljning av vin i små mängder direkt till konsumenten, med undantag för de detaljister som har vinkällare avsedda för lagring och tappning av stora mängder vin.
Artikel 7
Den information som innefattas i de deklarationer som avses i första stycket skall behandlas centralt på nationell nivå.
2. Medlemsstater vars vinodlingsareal inte överstiger 100 ha och som har
De medlemsstater i vilka kapitlen I och II i avdelning II i förordning (EG) nr 1493/1999 inte tillämpas i enlighet med artikel 21 i den förordningen och som har
Artikel 8
Artikel 9
Medlemsstaterna får fastställa koefficienter för konvertering av mängder så att andra produkter kan uttryckas som hektoliter vin. Koefficienterna får anpassas efter olika objektiva kriterier som påverkar konverteringen. Medlemsstaterna skall meddela kommissionen koefficienterna samtidigt som det sammandrag lämnas in som avses i artikel 14.
Denna förordning skall inte påverka medlemsstaternas bestämmelser om skörde-, produktions-, behandlingsoch/eller saluförings- eller lagerdeklarationer som är avsedda att ge mer fullständig information, i synnerhet genom att de omfattar en bredare krets av personer än de som avses i artiklarna 2, 4 och 6.
2. De deklarationer som avses i artikel 6 skall lämnas senast den 10 september för de kvantiteter som innehas den 31 juli. Medlemsstaterna får emellertid fastställa ett eller flera tidigare datum.
Dock gäller att om de frister som avses i första stycket överskrids med högst fem arbetsdagar skall de belopp som skall utbetalas för innevarande vinår minskas med 15 %. Om fristerna överskrids med högst tio arbetsdagar skall beloppen minskas med 30 %.
2. Om medlemsstaternas behöriga myndigheter finner att de deklarationer som avses i denna förordning är ofullständiga eller oriktiga, och om de felaktiga eller ej införda uppgifterna är nödvändiga för en korrekt tillämpning av de åtgärder som avses i punkt 1 skall medlemsstaten, utom i fall av force majeure, tillämpa följande påföljder, utan att det påverkar nationella påföljder.
- två gånger det konstaterade felets procentsats om felet medför att den deklarerade volymen justeras med mer än 5 % men högst 20 %.
b) När det gäller de åtgärder som avses i artiklarna 29 och 30 i förordning (EEG) nr 1493/1999 skall det pris som destillatören skall betala till den deklarerande producenten, om det vin som levereras till destillation ännu inte har betalats, minskas i följande omfattning:
Om den oriktighet som fastställts i deklarationen kan hänföras till information från andra aktörer eller anslutna vilkas namn finns med i de föreskrivna handlingarna och inte kan kontrolleras i förväg av deklaranten skall priserna endast minskas med procentsatsen för justeringen.
Medlemsstaterna skall vid datum som möjliggör för de meddelanden enligt artikel 16 upprätta följande:
c) En bedömning för pågående vinår av den volym vinprodukter som kan förväntas framställas i medlemsstaten.
Artikel 15
3. På de valda platserna skall var fjortonde dag priset på vita och röda bordsviner utan geografisk beteckning och den saluförda volymen av dessa viner noteras på lämpligt sätt.
1. Medlemsstaterna skall meddela kommissionen
c) senast den 30 november, de uppgifter som gör det möjligt att uppskatta de tillgängliga mängderna vinprodukter och deras användning i medlemsstaten enligt artikel 14 d,
2. Medlemsstaterna skall meddela kommissionen
- En beräkning av produktionen under de fem senaste vinåren för de områden som samlats inom produktionsområdet.
b) Från och med den 1 augusti 2001 skall medlemsstaterna varannan tisdag meddela kommissionen priser och volymer för saluförda produkter tillsammans med alla övriga uppgifter som bedöms vara till hjälp för att bedöma marknadsutvecklingen i produktionsområdet.
Artikel 18
Kommissionen ansvarar för att de uppgifter som mottas i enlighet med denna förordning sprids.
a) Producenten har inte lämnat in skörde-, produktions- eller lagerdeklarationen inom fastställda tidsfrister.
Det belopp söm skall återvinnas fastställs enligt reglerna i artikel 13 i förordning (EG) nr 1282/2001.
Artikel 21
Artikel 22
av den 29 juni 2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Vid fastställandet av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemdel i livsmedel med animaliskt ursprung är det nödvändigt att ange de djurarter i vilka restmängder kan förekomma, vilka mängder som kan förekomma i var och en av de relevanta vävnaderna från det behandlade djuret (målvävnad) samt vilket slag av restmängd som är relevant vid övervakningen av restmängder (restmarkör).
(6) Florfenikol bör införas i bilaga I till förordning (EEG) nr 2377/90.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 23 juli 2001
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Vid det nionde sammanträdet med parterna i Konventionen om internationell handel med utrotningshotade arter av vilda djur och växter (CITES) 1994 krävdes att åtgärder för bevakning av uppgifter om fångster av och handel med arter av Elasmobranchii-fiskar (hajar och rockor) skulle vidtas av FN:s livsmedels- och jordbruksorganisation (FAO) och av regionala fiskeorganisationer.
(4) I artikel 4.2 i förordning (EEG) nr 3880/91 föreskrivs att medlemsstaterna efter att i förväg ha inhämtat medgivande från Eurostat, får lämna uppgifter i annan form eller med annat medium än enligt vad som föreskrivs i bilaga IV till förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EG) nr 1623/2000 om tillämpningsföreskrifter för rådets förordning (EG) nr 1493/1999 om den gemensamma organisationen av marknaden för vin, vad beträffar marknadsmekanismerna
med beaktande av rådets förordning (EG) nr 1493/1999 av 17 maj 1999 om den gemensamma organisationen av marknaden för vin(1), senast ändrad genom förordning (EG) nr 2826/2000(2), särskilt artiklarna 33 och 36 i denna, och
(2) I artikel 63 föreskrivs inrättandet av en stödordning för destillation av vin till spritdrycker. Denna ordning tilllämpades första gången under vinåret 2000/2001. Mot bakgrund av de erfarenheter som gjorts under det första tillämpningsåret bör ändringar införas. Bland annat bör destillationen inledas senare på året och andelen av vinproducentens produktion som får gå till denna destillation bör sänkas. Dessutom bör ett slutdatum införas för destillation.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.!
1. Artikel 58 första stycket skall ersättas med följande: "De producenter som omfattas av någon av skyldigheterna enligt artiklarna 45 och 52 i den här förordningen och som före den 15 juli innevarande vinår har levererat minst 90 % av sin ålagda kvantitet kan uppfylla denna skyldighet genom att leverera resterande kvantitet före ett datum som den behöriga nationella myndigheten skall fastställa, dock inte senare än den 31 juli påföljande vinår."
2. Kvantiteten bordsvin, och vin som lämpar sig för framställning av bordsvin, som varje producent får lämna till destillation, skall begränsas till 30 % av dennes maximiproduktion av dessa viner som deklarerats under de tre senaste vinåren, inklusive det innevarande om deklarationen redan lämnats. Om den ovan angivna procentsatsen tillämpas, skall den producerade mängden bordsvin vara den som anges som vin i kolumnen 'bordsvin' i produktionsdeklarationen enligt artikel 18.1 i förordning (EG) nr 1493/1999."
4. Artikel 91.12 skall ersättas med följande: "12. Säkerheten för att garantera att alkoholen exporteras skall, av det interventionsorgan som innehar den, frisläppas för varje kvantitet som bevisligen har exporterats inom föreskriven tidsfrist. Om tidsfristen för export överskrids skall, genom undantag från artikel 23 i förordning (EEG) nr 2220/85, och utom i fall av force majeure, denna exportsäkerhet på 3 euro per hektoliter hundraprocentig alkoholvara förverkas
5. Artikel 95.2 andra och tredje styckerna skall ersättas med följande: "Alkohol i behållare som inte anges i meddelandena om anbudsinfordran och offentlig auktion, eller i det beslut av kommissionen som avses i artiklarna 83-93 i den här förordningen, skall inte omfattas av detta förbud.
a) Punkt 1 skall ersättas med följande: "1. Från och med offentliggörandet av ett meddelande om anbudsförfarande och fram till sista dagen för inlämnande av anbud kan alla intresserade parter, mot betalning av 10 euro per liter, erhålla prover av den alkohol som bjuds ut. Kvantiteten per intresserad part får inte överstiga 5 liter per behållare. För avsättningen enligt delavsnitt III kan varuprovet erhållas, mot samma betalning, inom 30 dagar efter meddelandet om offentlig auktion."
b) får de anbudsgivare som erbjudits en ersättningsmängd enligt artikel 83.3 i den här förordningen erhålla prover av den alkohol som erbjuds som ersättning.
Artikel 2
av den 22 augusti 2001
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
(1) I artikel 1 i kommissionens förordning (EG) nr 174/1999 av den 26 januari 1999 om fastställande av särskilda tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 i fråga om exportlicenser och exportbidrag inom sektorn för mjölk och mjölkprodukter(3), senast ändrad genom förordning (EG) nr 1370/2001(4), fastställs som generell regel att en exportlicens skall uppvisas vid all export av mjölkprodukter för vilken exportbidrag begärs. För att få en effektiv förvaltning av den inre marknaden för skummjölkspulver, en produkt för vilken interventionsåtgärder kan bli aktuella, är det nödvändigt att exportlicensen blir obligatorisk och att medlemsstaterna skall ha skyldighet att meddela kommissionen uppgifter om dessa licenser. Därför bör kommissionens förordning (EG) nr 1498/1999 av den 8 juli 1999 om tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 beträffande meddelanden mellan medlemsstaterna och kommissionen med avseende på mjölk och mjölkprodukter(5), senast ändrad genom förordning (EG) nr 732/2001(6), ändras.
(4) För slutliga licenser för export utan bidrag till Förenta staterna inom den tilläggskvot som är en följd av jordbruksavtalet inom ramen för GATT:s Uruguayrunda(7) (nedan kallat jordbruksavtalet) behöver ingen säkerhet ställas. För att se till att denna kvot i möjligaste mån utnyttjas fullt ut och att de licenser som utfärdats används, bör en säkerhet ställas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 1.1 skall följande stycke läggas till: "Genom undantag från första stycket skall emellertid en exportlicens uppvisas vid all export av sådana produkter som avses i bilaga I kategori II."
4. I artikel 20.2 andra stycket skall "9 euro" ersättas med "6 euro".
Säkerheten för den slutliga licensen får endast frisläppas mot uppvisande av det bevis som avses i artikel 35.5 i förordning (EG) nr 1291/2000(8)."
a) De kvantiteter, fördelade efter nummer i exportbidragsnomenklaturen för mjölkprodukter och efter kod för bestämmelseort, för vilka licens har begärts samma dag,
c) De kvantiteter, fördelade efter nummer i exportbidragsnomenklaturen för mjölkprodukter och efter kod för bestämmelseort, för vilka sådana tillfälliga licenser som avses i artikel 8 i förordning (EG) nr 174/1999 slutligt utfärdats eller dragits in samma dag, med angivande av från vilket organ anbudsinfordran kommer, samt dessutom datum och kvantitet för den tillfälliga licensen.
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av rådets förordning (EG) nr 723/97 om genomförande av medlemsstaternas åtgärdsprogram på området för kontroll av utgifterna för EUGFJ:s garantisektion
med beaktande av kommissionens förslag(1),
(1) Enligt artikel 1 i förordning (EG) nr 723/97(3) skall gemenskapen delta i de kostnader som medlemsstaterna ådragit sig för att genomföra de nya åtgärdsprogram som följer av nya skyldigheter gentemot gemenskapen, vilka har godkänts av kommissionen och vars syfte är att förbättra strukturen hos och effektiviteten av kontrollen när det gäller utgifterna för EUGFJ:s garantisektion. Enligt artikel 4 i förordningen skall det finansiella bidraget från gemenskapen beviljas per kalenderår under en tid av fem år i följd räknat från år 1997. Det skall beviljas inom ramen för de årliga anslag som beviljas av budgetmyndigheten inom ramen för budgetplanen.
(4) Den period under vilken det finansiella bidraget från gemenskapen kan betalas bör därför förlängas med två år.
Artikel 1
Kommissionens förordning (EG) nr 2601/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Inga invändningar enligt artikel 7 i förordning (EEG) nr 2081/92 har framställts till kommissionen till följd av offentliggörandet i Europeiska gemenskapernas officiella tidning(3) av de produktnamn som anges i bilagan till den här förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 4 februari 2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) I kommissionens förordning (EG) nr 194/97 av den 31 januari 1997 om fastställande av högsta tillåtna halt för vissa främmande ämnen i livsmedel(2), senast ändrad genom förordning (EG) nr 1566/1999(3), fastställs högsta tillåtna halter för vissa främmande ämnen i livsmedel, särskilt för aflatoxiner. Dessa gränsvärden har vida överskridits i prov tagna från jordnötter som har sitt ursprung i eller försänds från Kina.
(6) Jordnötter och produkter framställda av jordnötter måste produceras, sorteras, hanteras, bearbetas, förpackas och transporteras under goda hygieniska förhållanden. Halterna av aflatoxin B1 och den totala aflatoxinhalten måste fastställas i prover som tas ur sändningar just innan de lämnar Kina.
(9) För att skydda folkhälsan måste därför de behöriga myndigheterna i den importerande medlemsstaten ta prover på alla sändningar av jordnötter som har sitt ursprung i eller försänds från Kina och som importeras till Europeiska gemenskapen och analysera dessa prover med avseende på aflatoxinhalten, innan jordnötterna släpps ut på marknaden. Eftersom denna åtgärd tar en betydande del av medlemsstaternas kontrollresurser i anspråk, kommer resultaten av åtgärden att utvärderas efter en kort period och åtgärderna ändras vid behov.
Artikel 1
- Jordnötter som omfattas av KN-nummer 2008 11 94 (i förpackningar med en nettovikt på mer än 1 kg) eller 2008 11 98 (i förpackningar med en nettovikt på mindre än 1 kg).
3. Varje sändning skall märkas med samma beteckning som den som anges i hälsointyget och i den bifogade rapporten med resultaten från den officiella provtagningen och analysen som avses i punkt 1.
Artikel 2
om ändring av Europaparlamentets beslut 94/262/EGKS, EG, Euratom om föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 195.4,
med beaktande av Europaparlamentets resolution av den 17 november 2000 om ändring av Europaparlamentets beslut av den 9 mars 1994 om föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning(1),
av följande skäl:
(3) Det är därför nödvändigt att ändra beslut 94/262/EKSG, EG, Euratom och Europaparlamentet av den 9 mars 1994 om föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning(3) eftersom det i detta beslut föreskrivs att ombudsmannens budget skall utgöra bilaga till avsnitt I (Europaparlamentet) i Europeiska gemenskaperna allmänna budget.
Artikel 1
Kommissionens beslut
(Text av betydelse för EES)
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, och
(2) För genomförandet av de regleringsuppgifter som anges i dessa direktiv har nationella regleringsmyndigheter inrättats i samtliga medlemsstater, och dessa myndigheter skall anmälas till kommissionen i enlighet med artikel 3.6 i ramdirektivet. Enligt ramdirektivet skall medlemsstaterna också garantera den oberoende ställningen hos sina nationella regleringsmyndigheter genom att sörja för att de hålls rättsligt åtskilda från och verksamhetsmässigt oberoende av alla organisationer som tillhandahåller nät, utrustning eller tjänster för elektronisk kommunikation. Medlemsstater som behåller äganderätten till eller kontrollen över företag som tillhandahåller elektroniska kommunikationsnät eller kommunikationstjänster skall också sörja för att en praktiskt fungerande organisatorisk åtskillnad görs mellan regleringsverksamhet och sådan verksamhet som har samband med ägande eller kontroll.
(5) En europeisk grupp av regleringsmyndigheter för nät och tjänster inom området elektronisk kommunikation (nedan kallad gruppen) bör bildas. Avsikten är att den skall fungera som förmedlande länk för samråd med och experthjälp åt kommissionen inom området elektronisk kommunikation.
(8) Gruppen bör bedriva nära samarbete med den kommunikationskommitté som inrättats i enlighet med ramdirektivet. Gruppen bör verka på ett sådant sätt så att den inte inkräktar på kommitténs arbete.
Artikel 1
Artikel 2
Artikel 3
Gruppen skall fungera som en förmedlande länk mellan nationella regleringsmyndigheter och kommissionen på sådant sätt att den bidrar till den inre marknadens utveckling och till att regelverket för nät och tjänster inom området elektronisk kommunikation tillämpas på ett enhetligt sätt i alla medlemsstater.
Gruppen skall vara sammansatt av cheferna för respektive medlemsstaters nationella regleringsmyndigheter eller av deras ombud.
Arbetsordning
Ordföranden skall kalla gruppen till sammanträde efter överenskommelse med kommissionen.
Sakkunniga från EES-länder samt från kandidatländerna för anslutning till Europeiska unionen får delta som observatörer i gruppen. Gruppen får kalla andra sakkunniga och observatörer att närvara vid sina möten.
Gruppen skall i ett tidigt skede genomföra omfattande samråd med marknadsaktörer, konsumenter och slutförbrukare på ett sätt som garanterar öppenhet och insyn.
Utan att det påverkar tillämpningen av bestämmelserna i artikel 287 i fördraget, skall gruppens ledamöter, liksom dess observatörer och alla andra personer - i de fall kommissionen upplyser dem om att de rådgivande yttranden som begärts in eller de frågor väckts är av konfidentiell art - vara förpliktade att inte röja uppgifter som har kommit till deras kännedom genom arbetet i gruppen, dess undergrupper eller sakkunniggrupper. Kommissionen får i sådana fall besluta att enbart gruppens ledamöter får närvara vid mötena i fråga.
Gruppen skall lämna en årsberättelse över sin verksamhet till kommissionen. Kommissionen skall överlämna årsberättelsen till Europaparlamentet och rådet, i tillämpliga fall med sina kommentarer bifogade.
Detta beslut träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
om ändring av beslut 94/652/EG om uppdatering av inventeringen och uppgifterna inom ramen för medlemsstaternas samarbete vid den vetenskapliga granskningen av livsmedelsfrågor
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) I kommissionens beslut 94/458/EG(2) fastställs bestämmelser om den administrativa organisationen av samarbetet vid den vetenskapliga granskningen av livsmedelsfrågor.
(4) Uppgifterna bör fördelas med hänsyn till den vetenskapliga kompetens och de resurser som finns i medlemsstaterna och särskilt de institut som kommer att delta i det vetenskapliga samarbetet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 11 mars 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 137.2 i detta,
med beaktande av Regionkommitténs yttrande(3),
(1) Enligt artikel 136 i fördraget skall gemenskapen och medlemsstaterna särskilt ha som mål att främja en dialog mellan arbetsmarknadens parter.
(4) Kommissionen ansåg efter detta samråd att en gemenskapsåtgärd var önskvärd och samrådde på nytt med arbetsmarknadens parter om det planerade förslagets innehåll; arbetsmarknadens parter har inkommit med yttranden till kommissionen.
(7) Det finns behov av att förstärka den sociala dialogen och öka det ömsesidiga förtroendet inom företagen för att göra det lättare att föregripa risker, göra arbetsorganisationen mer flexibel och underlätta arbetstagarnas tillgång till utbildning inom företaget under trygga förhållanden, öka arbetstagarnas medvetenhet om behoven av anpassning, stimulera arbetstagarna att medverka i åtgärder och insatser för att öka deras anställbarhet, främja arbetstagarnas medverkan i företagets verksamhet och framtid samt stärka företagets konkurrenskraft.
(10) Gemenskapen har utarbetat och genomfört en sysselsättningsstrategi som vilar på begreppen "föregripande", "förebyggande" och "anställbarhet", som skall bli hörnstenar i all offentlig politik som kan inverka positivt på sysselsättningen, även den som utformas inom företagen, genom en intensifiering av dialogen mellan arbetsmarknadens parter för att främja sådana förändringar som är förenliga med bibehållandet av det prioriterade sysselsättningsmålet.
(13) Gemenskapens och medlemsstaternas nuvarande rättsliga ramar för information till och samråd med arbetstagare är ofta i alltför hög grad inriktade på hur man hanterar förändringsprocesser i efterhand, samtidigt som de bortser från de ekonomiska aspekterna av besluten och inte främjar ett verkligt föregripande av sysselsättningsutvecklingen i företag eller förebyggande av risker.
(16) Detta direktiv påverkar inte de system som föreskriver direkt deltagande av arbetstagarna, under förutsättning att dessa fortfarande har möjlighet att utöva rätten till information och samråd genom sina representanter.
(19) Denna allmänna ram bör också syfta till att undvika sådana administrativa, ekonomiska och rättsliga förpliktelser som kan motverka etableringen och utvecklingen av små och medelstora företag. Det förefaller därför rimligt att enligt medlemsstaternas val begränsa tillämpningsområdet för detta direktiv till företag med minst 50 arbetstagare eller till driftställen med minst 20 arbetstagare.
(22) Gemenskapsramen för information till och samråd med arbetstagare bör i så hög grad som möjligt begränsa de bördor som läggs på företagen eller driftsställena men likväl säkerställa ett effektivt utövande av rättigheterna.
(25) Företagen och driftställena bör skyddas mot att viss särskilt känslig information lämnas ut.
(28) Administrativa eller rättsliga förfaranden och sanktioner som är effektiva och avskräckande samt står i proportion till hur allvarlig övertädelsen är bör tillämpas när skyldigheterna i detta direktiv inte uppfylls.
(31) Genomförandet av detta direktiv bör inte anses vara ett tillräckligt skäl för att rättfärdiga en sänkning av arbetstagarnas allmänna skyddsnivå på det område som omfattas av direktivet.
Syfte och principer
3. När formerna för information eller samråd fastställs och genomförs, skall arbetsgivaren och arbetstagarrepresentanterna arbeta i samförståndsanda med respekt för varandras ömsesidiga rättigheter och skyldigheter samt med beaktande av såväl företagets eller driftställets intressen som arbetstagarnas intressen.
I detta direktiv avses med
c) arbetsgivare: en fysisk eller juridisk person som är part i ett anställningsavtal eller anställningsförhållande gentemot en arbetstagare i enlighet med nationell lagstiftning och nationell praxis,
f) information: arbetsgivarens överlämnande av uppgifter till arbetstagarrepresentanterna som gör det möjligt för dem att sätta sig in i vad den behandlade frågan avser och att granska densamma,
Räckvidd
b) driftställen som i en medlemsstat sysselsätter minst 20 arbetstagare.
3. Medlemsstaterna får göra undantag från detta direktiv genom särskilda bestämmelser för besättningar på fartyg som trafikerar öppet hav.
1. I enlighet med principerna i artikel 1 och utan att det påverkar tillämpningen av gällande bestämmelser och/eller praxis som är mer gynnsamma för arbetstagarna, skall medlemsstaterna besluta om formerna för rätt till information och samråd på lämplig nivå i enlighet med denna artikel.
b) Information och samråd om situationen, strukturen och den förväntade utvecklingen när det gäller sysselsättningen i företaget eller driftstället samt om eventuella föregripande åtgärder som planeras, bland annat vid hot mot sysselsättningen.
4. Samråd skall äga rum
c) på grundval av de uppgifter som arbetsgivaren lämnat i enlighet med artikel 2 f) och det yttrande som arbetstagarrepresentanterna har rätt att avge,
Artikel 5
Artikel 6
2. I särskilda fall och på de villkor och med de begränsningar som fastställs i nationell lagstiftning skall medlemsstaterna föreskriva att arbetsgivaren inte är skyldig att lämna ut sådan information eller inleda sådant samråd som utifrån objektiva kriterier skulle skada företaget eller driftstället eller vara till allvarligt förfång för dess verksamhet.
Skydd för arbetstagarrepresentanterna
Tillvaratagande av rättigheterna
Artikel 9
2. Detta direktiv skall inte påverka de bestämmelser som antagits i enlighet med direktiv 94/45/EG och direktiv 97/74/EG.
Artikel 10
a) företag med minst 150 anställda eller driftställen med minst 100 anställda till och med den 23 mars 2007, och
Genomförande av direktivet
Artikel 12
Artikel 13
Artikel 14
Europaparlamentets och rådets direktiv 2002/61/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
(1) Arbetet med att upprätta den inre marknaden bör stegvis förbättra livskvaliteten samt hälso- och konsumentskyddet. Åtgärderna i detta direktiv säkerställer en hög hälso- och konsumentskyddsnivå.
(4) Vetenskapliga kommittén för toxicitet, ekotoxicitet och miljö har efter det att kommissionen samrått med den bekräftat att cancerrisken som orsakas av textilier och läderartiklar som färgats med vissa azofärgämnen ger anledning till oro.
(7) Tillämpningen av detta direktiv kräver harmoniserade analysmetoder. Kommissionen bör fastställa sådana metoder i enlighet med artikel 2a i direktiv 76/769/EEG. Analysmetoderna bör företrädesvis utarbetas på europeisk nivå, om så är lämpligt av Europeiska standardiseringskommittén (CEN).
(10) Detta direktiv påverkar inte tillämpningen av gemenskapens lagstiftning om minimikrav för arbetarskydd i rådets direktiv 89/391/EEG(5) och i särdirektiv som grundas på det direktivet, i synnerhet rådets direktiv 90/394/EEG(6) och Europaparlamentets och rådets direktiv 98/24/EG(7).
Bilaga I till direktiv 76/769/EEG ändras härmed i enlighet med bilagan till det här direktivet.
De skall tillämpa dessa bestämmelser från och med 11 september 2003.
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets direktiv 2002/85/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) I rådets direktiv 92/6/EEG(4) anges att kraven på montering och användning av hastighetsbegränsande anordningar senare kan utvidgas till att omfatta lättare nyttofordon, beroende på de tekniska möjligheterna och erfarenheterna i medlemsstaterna.
(6) Eftersom målen för den föreslagna åtgärden, nämligen att ändra gemenskapsbestämmelserna om montering och användning av hastighetsbegränsande anordningar i vissa tunga motorfordonskategorier, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför på grund av åtgärdens omfattning och verkningar bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
Artikel 1
"Artikel 1
Artikel 2
Artikel 3
Artikel 4
b) fordon som registrerats mellan den 1 januari 1988 och den 1 januari 1994,
2. När det gäller motorfordon i kategori M2, fordon i kategori M3 med en totalvikt på över 5 ton men högst 10 ton samt fordon i kategori N2, skall artiklarna 2 och 3 senast tillämpas på
i) från och med den 1 januari 2006, om det rör sig om fordon som används för såväl nationella som internationella transporter,
Artikel 5
2. Följande artikel skall läggas till:
Kommissionen skall vid behov lägga fram lämpliga förslag.".
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 4
av den 16 december 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 47.2 i detta,
efter att ha hört Regionkommittén,
av följande skäl:
(3) I kommissionens handlingsplan för finansiella tjänster utpekas en rad åtgärder som krävs för att fullborda den inre marknaden för finansiella tjänster, och det aviseras att det skall utarbetas lagstiftning om extra tillsyn för finansiella konglomerat i syfte att eliminera kryphål i den nuvarande särlagstiftningen och hantera ytterligare stabilitetsrisker för att på så sätt säkra sunda arrangemang för tillsyn över finansiella grupper med sektorsöverskridande finansiell verksamhet. Ett så ambitiöst mål kan bara uppnås stegvis. Införandet av extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat utgör ett sådant steg.
(6) Beslut att inte låta en viss enhet omfattas av räckvidden för den extra tillsynen bör fattas med beaktande bl.a. av om en sådan enhet omfattas av tillsynen på gruppnivå enligt särreglerna.
(9) Samtliga finansiella konglomerat som omfattas av den extra tillsynen bör ha en samordnare som utses bland berörda behöriga myndigheter.
(12) Det finns ett trängande behov av ett ökat samarbete mellan de myndigheter som ansvarar för tillsynen över kreditinstitut, försäkringsföretag och värdepappersföretag, inbegripet att utveckla särskilda arrangemang för samarbete mellan de myndigheter som är delaktiga i tillsynen över enheter som ingår i samma finansiella konglomerat.
(15) Av detta direktiv följer inte att de behöriga myndigheterna till Kommittén för finansiella konglomerat skall lämna ut information som är belagd med sekretess enligt detta direktiv eller andra sektorsdirektiv.
(18) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(5).
(21) För att man skall kunna bedöma behovet av ytterligare harmonisering av behandlingen av kapitalförvaltningsbolag som omfattas av särregler och förbereda denna harmonisering bör kommissionen rapportera om medlemsstaternas praxis på detta område.
MÅL OCH DEFINITIONER
I detta direktiv fastställs regler för extra tillsyn över reglerade enheter som har erhållit auktorisation enligt artikel 6 i direktiv 73/239/EEG, artikel 6 i direktiv 79/267/EEG, artikel 3.1 i direktiv 93/22/EEG eller artikel 4 i direktiv 2000/12/EG och som ingår i ett finansiellt konglomerat. Genom direktivet ändras också berörda särregler för enheter som regleras av ovannämnda direktiv.
I detta direktiv används följande beteckningar med de betydelser som här anges:
3. värdepappersföretag: ett värdepappersföretag i den mening som avses i artikel 1.2 i direktiv 93/22/EEG, inbegripet företag som avses i artikel 2.4 i direktiv 93/6/EEG.
6. återförsäkringsföretag: ett återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG.
a) Ett kreditinstitut, ett finansiellt institut eller ett företag som tillhandahåller tjänster anknutna till bankverksamhet enligt artikel 1.5 och 1.23 i direktiv 2000/12/EG (banksektorn).
d) Ett blandat finansiellt holdingföretag.
11. ägarintresse: ett ägarintresse i den mening som avses i artikel 17 första meningen i rådets fjärde direktiv 78/660/EEG av den 25 juli 1978 om årsbokslut i vissa typer av bolag(16) eller direkt eller indirekt ägande av 20 % eller mer av rösterna eller kapitalet i ett företag.
a) ägarintresse, innebärande ett innehav, direkt eller genom kontroll av 20 % eller mer av rösterna eller kapitalet i ett företag, eller
14. finansiellt konglomerat: en grupp som uppfyller följande villkor, om inte annat följer av artikel 3:
c) Om ingen reglerad enhet i den mening som avses i artikel 1 finns i toppen av gruppen, bedrivs gruppens verksamhet huvudsakligen inom den finansiella sektorn i den mening som avses i artikel 3.1.
Varje undergrupp till en grupp enligt punkt 12 som uppfyller kriterierna i denna punkt skall anses vara ett finansiellt konglomerat.
17. relevanta behöriga myndigheter:
c) andra berörda behöriga myndigheter, om de myndigheter som anges under a och b anser detta vara relevant. Vid en sådan bedömning skall särskilt beaktas den marknadsandel de reglerade enheterna i konglomeratet har i andra medlemsstater, i synnerhet om den överstiger 5 %, och den betydelse varje reglerad enhet som är etablerad i en annan medlemsstat har inom konglomeratet.
Artikel 3
2. För att verksamheten inom olika finansiella sektorer skall bedömas som betydande i den mening som avses i artikel 2.14 e, skall för varje finansiell sektor genomsnittet av kvoten mellan denna finansiella sektors balansomslutning och den totala balansomslutningen för gruppens enheter inom finansiella sektorer och kvoten mellan solvenskraven för denna finansiella sektor och de totala solvenskraven för gruppens enheter inom finansiella sektorer överstiga 10 %.
a) Den relativa storleken på dess minsta finansiella sektor överstiger inte 5 %, mätt antingen i termer av det genomsnitt som anges i punkt 2 eller i termer av balansomslutningen eller solvenskraven för en sådan finansiell sektor.
4. För tillämpningen av punkterna 1, 2 och 3 får de relevanta behöriga myndigheterna i samförstånd
När ett finansiellt konglomerat har identifierats enligt punkterna 1, 2 och 3 skall de beslut som avses i första stycket och detta stycke fattas på grundval av ett förslag från samordnaren för detta finansiella konglomerat.
Vid tillämpningen av punkt 3 skall, om balansomslutningen för den minsta finansiella sektorn inom gruppen understiger 6 miljarder euro för konglomerat som redan är föremål för extra tillsyn, även ett lägre belopp om 5 miljarder euro tillämpas under de tre följande åren, för att plötsliga byten av tillämpligt regelverk skall kunna undvikas.
De solvenskrav som avses i punkterna 2 och 3 skall beräknas enligt bestämmelserna i de relevanta särreglerna.
1. De behöriga myndigheter som har auktoriserat reglerade enheter skall på grundval av artiklarna 2, 3 och 5 identifiera varje grupp som omfattas av detta direktivs räckvidd.
- skall en behörig myndighet som anser att en av denna myndighet auktoriserad reglerad enhet tillhör en grupp som kan vara ett finansiellt konglomerat, som inte redan har identifierats enligt detta direktiv, underrätta de andra berörda behöriga myndigheterna om sin inställning.
EXTRA TILLSYN
Artikel 5
2. Följande reglerade enheter skall underkastas extra tillsyn på nivån finansiella konglomerat i enlighet med artiklarna 6-17:
c) Varje reglerad enhet som har ett sådant samband med en annan enhet i den finansiella sektorn som avses i artikel 12.1 i direktiv 83/349/EEG.
4. Om personer har ägarintresse i eller kapitalförbindelser med en eller flera reglerade enheter eller utövar ett betydande inflytande över sådana enheter utan att ha ägarintresse eller kapitalförbindelser utöver de fall som avses i punkterna 2 och 3, skall de relevanta behöriga myndigheterna i samförstånd och i enlighet med den nationella lagstiftningen avgöra huruvida och i vilken omfattning extra tillsyn skall utövas över dessa reglerade enheter som om de utgjorde ett finansiellt konglomerat.
5. Utan att det påverkar tillämpningen av artikel 13 skall utövandet av extra tillsyn på nivån finansiellt konglomerat inte på något sätt anses innebära att de behöriga myndigheterna är skyldiga att utöva tillsyn över blandade finansiella holdingföretag, över reglerade enheter i tredje land som tillhör ett finansiellt konglomerat eller över enskilda icke reglerade enheter i ett finansiellt konglomerat.
Artikel 6
2. Medlemsstaterna skall kräva att reglerade enheter i ett finansiellt konglomerat säkerställer att det finns en tillgänglig kapitalbas på nivån finansiellt konglomerat som alltid minst motsvarar de kapitaltäckningskrav som beräknas enligt bilaga I.
Samordnaren skall se till att den beräkning som avses i första stycket utförs minst en gång per år, antingen av de reglerade enheterna eller av det blandade finansiella holdingföretaget.
a) Kreditinstitut, finansiella institut eller företag som tillhandahåller tjänster anknutna till bankverksamhet i den mening som avses i artikel 1.5 och 1.23 i direktiv 2000/12/EG.
d) Blandade finansiella holdingföretag.
5. Samordnaren kan besluta att inte inbegripa en viss enhet vid beräkningen av den extra kapitaltäckningskraven i följande fall:
c) Om det skulle vara olämpligt eller missvisande att inbegripa enheten med hänsyn till målen för den extra tillsynen.
Om samordnaren inte inkluderar en reglerad enhet i tillämpningsområdet med stöd av ett av de fall som anges i b och c i första stycket, får de behöriga myndigheterna i den medlemsstat där denna enhet är belägen begära att den enhet som finns i toppen av det finansiella konglomeratet lämnar upplysningar som underlättar tillsynen över den reglerade enheten.
1. Utan att särreglerna åsidosätts skall extra tillsyn över riskkoncentrationen i de reglerade enheterna i ett finansiellt konglomerat utövas enligt reglerna i artikel 9.2-9.4 i avsnitt 3 i detta kapitel och i bilaga II.
3. Till dess att gemenskapens lagstiftning har samordnats ytterligare får medlemsstaterna fastställa kvantitativa gränser eller tillåta sina behöriga myndigheter att fastställa kvantitativa gränser eller vidta andra tillsynsåtgärder som skulle kunna uppfylla målen för extra tillsyn när det gäller riskkoncentration på nivån finansiellt konglomerat.
Transaktioner inom det finansiella konglomeratet
Den nödvändiga informationen skall överlämnas till samordnaren av den reglerade enhet i den mening som avses i artikel 1 som finns i toppen av det finansiella konglomeratet eller, när det finansiella konglomeratet inte leds av en reglerad enhet i den mening som avses i artikel 1, av det blandade finansiella holdingföretaget eller av den reglerade enhet i det finansiella konglomeratet som identifierats av samordnaren efter samråd med de övriga relevanta behöriga myndigheterna och med det finansiella konglomeratet.
4. När ett finansiellt konglomerat leds av ett blandat finansiellt holdingföretag, skall särregler om transaktioner inom det finansiella konglomeratet i den största finansiella sektorn i det finansiella konglomeratet tillämpas för hela den sektorn, inklusive det blandade finansiella holdingföretaget.
1. Medlemsstaterna skall kräva att det hos reglerade enheter på nivån finansiellt konglomerat finns erforderliga metoder för riskhantering och rutiner för intern kontroll, inbegripet sunda rapporterings- och redovisningsförfaranden.
b) En adekvat kapitaltäckningsstrategi för att kunna förutse den inverkan som deras affärsstrategi har på riskprofilen och kapitalkraven, så som de fastställts i enlighet med artikel 6 och bilaga I.
a) Adekvata mekanismer för kapitaltäckning för att identifiera och mäta samtliga materiella risker och på ett lämpligt sätt ställa kapitalbasen i relation till riskerna.
5. De metoder och mekanismer som avses i punkterna 1-4 skall övervakas av samordnaren.
Artikel 10
2. Utnämningen skall grunda sig på följande kriterier:
i) Om moderföretaget till en reglerad enhet är ett blandat finansiellt holdingföretag, skall samordningen utövas av den behöriga myndighet som har auktoriserat denna reglerade enhet enligt gällande särregler.
Om det finansiella konglomeratet leds av två eller flera blandade finansiella holdingföretag vilka har huvudkontor i olika medlemsstater och det finns en reglerad enhet i var och en av dessa medlemsstater, skall samordningen utövas av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som har den största balansomslutningen, om dessa enheter verkar inom samma finansiella sektor, eller av den behöriga myndighet som ansvarar för tillsynen över den reglerade enhet som verkar inom den största finansiella sektorn.
3. I särskilda fall får de relevanta behöriga myndigheterna i samförstånd bevilja undantag från de kriterier som anges i punkt 2, om det skulle vara olämpligt att tillämpa dessa kriterier, med beaktande av konglomeratets struktur och den relativa betydelsen av dess verksamhet i olika länder, och utse en annan behörig myndighet till samordnare. I dessa fall skall de behöriga myndigheterna innan de fattar sitt beslut ge konglomeratet möjlighet att yttra sig om detta beslut.
1. De uppgifter som samordnaren skall utföra inom ramen för den extra tillsynen skall omfatta följande:
c) Bedömning av huruvida reglerna om kapitaltäckning, riskkoncentration och transaktioner inom det finansiella konglomeratet enligt artiklarna 6, 7 och 8 följs.
f) Andra uppgifter, åtgärder och beslut som har tilldelats samordnaren genom detta direktiv eller som följer av detta direktivs tillämpning.
3. Utan att det påverkar möjligheten att delegera specifika tillsynsbefogenheter och specifikt tillsynsansvar enligt gemenskapslagstiftningen, skall förekomsten av en samordnare som anförtrotts specifika uppgifter i samband med den extra tillsynen över reglerade enheter i ett finansiellt konglomerat inte påverka de behöriga myndigheternas uppgifter och ansvar enligt särreglerna.
1. De behöriga myndigheter som ansvarar för tillsynen över reglerade enheter i ett finansiellt konglomerat och den behöriga myndighet som utses till samordnare för detta skall ha ett nära samarbete med varandra. Utan att det påverkar dessa myndigheters respektive ansvar enligt särreglerna skall de, oavsett om de är inrättade i samma medlemsstat, till varandra överlämna alla uppgifter som är väsentliga eller relevanta för de övriga behöriga myndigheternas utövande av tillsynsuppgifter enligt särreglerna och detta direktiv. Härvid skall de behöriga myndigheterna och samordnaren på begäran överlämna alla relevanta uppgifter och på eget initiativ överlämna alla väsentliga uppgifter.
b) Det finansiella konglomeratets strategier.
e) Organisation, riskhantering och system för intern kontroll på det finansiella konglomeratets nivå.
h) Större sanktioner och exceptionella åtgärder som de behöriga myndigheterna vidtar i enlighet med särreglerna eller detta direktiv.
a) Sådana förändringar av aktieägar-, organisations- eller ledningsstrukturen i reglerade enheter i ett finansiellt konglomerat som kräver de behöriga myndigheternas godkännande eller auktorisation.
3. När de behöriga myndigheterna i den medlemsstat där ett moderföretag har sitt huvudkontor inte själva utövar den extra tillsynen enligt artikel 10, kan samordnaren begära att de av moderföretaget inhämtar alla uppgifter som kan vara relevanta för utövandet av samordningsuppgifterna enligt artikel 11 samt att de överlämnar dessa uppgifter till samordnaren.
Uppgifter som erhålls inom ramen för den extra tillsynen och särskilt varje utbyte av uppgifter mellan behöriga myndigheter eller mellan behöriga myndigheter och andra myndigheter enligt detta direktiv omfattas av särreglernas bestämmelser om tystnadsplikt och överlämnande av förtrolig information.
Medlemsstaterna skall kräva att de personer som faktiskt leder affärsverksamheten i ett blandat finansiellt holdingföretag har ett tillräckligt gott anseende och tillräcklig erfarenhet för att kunna fullgöra sina åligganden.
1. Medlemsstaterna skall säkerställa att det inte finns några rättsliga hinder inom deras jurisdiktion för att de fysiska och juridiska personer, vare sig dessa är reglerade enheter eller ej, som omfattas av extra tillsyn inbördes utbyter uppgifter som kan vara relevanta för den extra tillsynen.
Kontroll
Den behöriga myndighet som har framställt begäran får om den så önskar delta i kontrollen, om den inte själv utför den.
Om de reglerade enheterna i ett finansiellt konglomerat inte uppfyller de krav som anges i artiklarna 6-9 eller om kraven är uppfyllda men enheternas solvens ändå kan vara hotad eller om transaktionerna inom det finansiella konglomeratet eller riskkoncentrationerna utgör ett hot mot de reglerade enheternas finansiella ställning, skall nödvändiga åtgärder vidtas för att avhjälpa situationen så snart som möjligt
Utan att det påverkar tillämpningen av artikel 17.2 får medlemsstaterna bestämma vilka åtgärder som deras behöriga myndigheter får vidta när det gäller blandade finansiella holdingföretag.
De behöriga myndigheternas ytterligare befogenheter
AVSNITT 4
Moderföretag utanför gemenskapen
3. Medlemsstaterna skall tillåta sina behöriga myndigheter att tillämpa andra metoder som säkerställer lämplig extra tillsyn över reglerade enheter i ett finansiellt konglomerat. Metoderna måste godkännas av samordnaren, efter samråd med de andra relevanta behöriga myndigheterna. De behöriga myndigheterna kan särskilt kräva att det inrättas ett blandat finansiellt holdingföretag med huvudkontor inom gemenskapen och tillämpa detta direktiv på de reglerade enheterna i det finansiella konglomerat som leds av detta holdingföretag. Metoderna skall uppfylla de mål för den extra tillsynen som ställs upp i detta direktiv och skall rapporteras till de andra berörda behöriga myndigheterna och kommissionen.
1. Artikel 25.1 och 25.2 i direktiv 2000/12/EG och artikel 10a i direktiv 98/78/EG skall även tillämpas vid förhandlingar om avtal med ett eller flera tredje länder rörande metoder för utövande av extra tillsyn över reglerade enheter i ett finansiellt konglomerat.
KOMMISSIONENS BEFOGENHETER OCH KOMMITTÉFÖRFARANDE
1. Kommissionen skall, i enlighet med det förfarande som avses i artikel 21.2, anta tekniska ändringar av detta direktiv på följande områden:
c) Harmonisering av terminologin och ramarna för definitionerna i direktivet i överensstämmelse med framtida gemenskapsrättsakter om reglerade enheter och närliggande frågor.
2. Kommissionen skall underrätta allmänheten om alla förslag som läggs fram i enlighet med denna artikel och kommer att samråda med de berörda parterna, innan den överlämnar utkastet till åtgärder till den kommitté för finansiella konglomerat som anges i artikel 21.
1. Kommissionen skall bistås av en kommitté för finansiella konglomerat, nedan kallad "kommittén".
3. Kommittén skall själv anta sin arbetsordning.
6. Kommittén skall hållas underrättad av medlemsstaterna om de principer som de tillämpar för tillsynen över transaktioner inom det finansiella konglomeratet och riskkoncentration.
Artikel 22
1. Följande artikel skall läggas till:
a) är dotterföretag till ett försäkringsföretag som är auktoriserat i en annan medlemsstat,
2. Samråd med den behöriga myndigheten i en berörd medlemsstat som ansvarar för tillsynen över kreditinstitut eller värdepappersföretag skall genomföras innan auktorisation beviljas för ett försäkringsföretag som
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen.
"Från den disponibla solvensmarginalen skall även följande dras:
- återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG,
- värdepappersföretag och finansiella institut i den mening som avses i artikel 1.2 i direktiv 93/22/EEG(20) och i artiklarna 2.4 och 2.7 i rådets direktiv 93/6/EEG(21).
- De instrument som avses i artikel 18.3 i direktiv 79/267/EEG.
Som ett alternativ till avdrag av de poster enligt a och b i fjärde stycket som försäkringsföretag innehar i kreditinstitut, värdepappersföretag och finansiella institut, får medlemsstaterna tillåta att deras försäkringsföretag också tillämpar metoderna 1, 2 eller 3 i bilaga I till Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(22). Metod 1 (metod baserad på sammanställd redovisning) skall tillämpas endast om den behöriga myndigheten är säker på graden av samordnad förvaltning och intern kontroll avseende de enheter som skall inbegripas i tillämpningsområdet för sammanställningen. Den valda metoden skall tillämpas konsekvent över tiden.
Artikel 23
1. Följande artikel skall läggas till:
a) är dotterföretag till ett försäkringsföretag som är auktoriserat i en annan medlemsstat,
2. Samråd med den behöriga myndighet som ansvarar för tillsynen över kreditinstitut eller värdepappersföretag skall genomföras innan auktorisation beviljas för ett livförsäkringsföretag som
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett kreditinstitut eller värdepappersföretag som är auktoriserat i gemenskapen.
"Från den disponibla solvensmarginalen skall även följande avdrag göras:
- återförsäkringsföretag i den mening som avses i artikel 1 c i direktiv 98/78/EG,
- värdepappersföretag och finansiella institut i den mening som avses i artikel 1.2 i direktiv 93/22/EEG(26) och i artiklarna 2.4 och 2.7 i direktiv 93/6/EEG(27).
- De instrument som avses i artikel 16.3 i direktiv 73/239/EEG.
Med det avdrag av ägarintresse som anges i denna punkt menas här ägarintresse i den mening som avses i artikel 1 f i direktiv 98/78/EG.".
Direktiv 92/49/EEG ändras på följande sätt:
2. Artikel 16.5c skall ersättas med följande:
- i förekommande fall till andra myndigheter med ansvar för övervakning av betalningssystem,
Ändring av direktiv 92/96/EEG
"1a. Om köparen av det innehav som avses i punkt 1 är ett försäkringsföretag, ett kreditinstitut eller ett värdepappersföretag med auktorisation i en annan medlemsstat eller moderföretag till en sådan enhet, eller en fysisk eller juridisk person som har ägarkontroll över en sådan enhet, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av ett sådant samråd som avses i artikel 12a i direktiv 79/267/EEG.".
- till centralbanker och andra organ med liknande funktion i egenskap av monetära myndigheter,
Artikel 26
"- finansiellt holdingföretag: ett finansiellt institut vars dotterföretag antingen uteslutande eller huvudsakligen är värdepappersföretag eller andra finansiella institut av vilka åtminstone ett är ett värdepappersföretag, vilket inte är ett finansiellt holdingföretag med blandad verksamhet i den mening som avses i Europaparlamentets och rådets direktiv 2002/87/EG av den 16 december 2002 om extra tillsyn över kreditinstitut, försäkringsföretag och värdepappersföretag i ett finansiellt konglomerat(29).
Ändringar av direktiv 93/22/EEG
"Samråd med den behöriga myndighet i en berörd medlemsstat som har ansvar för tillsynen över kreditinstitut eller försäkringsföretag skall genomföras innan auktorisation beviljas för ett värdepappersföretag som
c) står under ägarkontroll av samma fysiska eller juridiska personer som har ägarkontrollen över ett kreditinstitut eller ett försäkringsföretag som är auktoriserat i gemenskapen.
"2. Om förvärvaren av det innehav som avses i punkt 1 är ett värdepappersföretag, ett kreditinstitut eller ett försäkringsföretag med auktorisation i en annan medlemsstat eller moderföretag till ett värdepappersföretag, ett kreditinstitut eller ett försäkringsföretag med auktorisation i en annan medlemsstat, eller en fysisk eller juridisk person som har ägarkontroll över ett värdepappersföretag, ett kreditinstitut eller ett försäkringsföretag med auktorisation i en annan medlemsstat, och om det företag som köparen vill förvärva ett innehav i som resultat av detta förvärv skulle komma att bli ett dotterföretag till köparen eller hamna under dennas ägarkontroll, skall bedömningen av förvärvet föregås av sådant samråd som avses i artikel 6.".
Direktiv 98/78/EG ändras på följande sätt:
h) anknutet företag: ett företag som är antingen ett dotterföretag eller ett annat företag som är föremål för ägarintresse eller ett företag som är knutet till ett annat företag genom ett sådant förhållande som avses i artikel 12.1 i direktiv 83/349/EEG.
2. I artikel 6.3 skall följande mening läggas till:
"Medlemsstaterna skall kräva att försäkringsföretagen följer adekvata metoder för riskhantering och rutiner för intern kontroll, inbegripet sunda rapporterings- och redovisningsförfaranden, för att på ett lämpligt sätt identifiera, mäta, övervaka och kontrollera transaktioner enligt bestämmelserna i punkt 1. Medlemsstaterna skall också kräva att försäkringsföretagen minst en gång om året rapporterar betydande transaktioner till de behöriga myndigheterna. Dessa förfaranden och betydande transaktioner skall övervakas av de behöriga myndigheterna.".
Samarbete med behöriga myndigheter i tredje land
b) försäkringsföretag i ett icke-medlemsland bland vars delägare det finns företag i den mening som avses i artikel 2 med huvudkontor inom gemenskapen.
b) att de behöriga myndigheterna i tredje land kan få fram den information som krävs för att utöva extra tillsyn över försäkringsföretag med huvudkontor inom deras territorier och med dotterföretag eller ägarintressen i företag i en eller flera medlemsstater.
Ledningsorgan för holdingföretag med blandad verksamhet
"Om det inte finns några kapitalband mellan vissa av företagen i en försäkringsgrupp, skall den behöriga myndigheten fastställa vilken proportionell andel som det skall tas hänsyn till.".
Reglerna om avdrag av ett sådant ägarintresse enligt artikel 16.1 i direktiv 73/239/EEG och artikel 18 i direktiv 79/267/EEG samt bestämmelserna om medlemsstaternas möjlighet att under vissa villkor tillåta alternativa metoder och att tillåta att ett sådant ägarintresse inte skall dras av, skall även tillämpas vid beräkningen av jämkad solvens hos ett försäkringsföretag som är ett företag med ägarintresse i ett kreditinstitut, ett värdepappersföretag eller ett finansiellt institut.".
Direktiv 2000/12/EG ändras på följande sätt:
"9. ägarintresse vid tillämpningen av gruppbaserad tillsyn och vid tillämpningen av artikel 34.2.15 och 34.2.16: ägarintresse i den mening som avses i artikel 17 första meningen i direktiv 78/660/EEG eller direkt eller indirekt innehav av 20 % eller mer av rösterna eller kapitalet i ett företag.".
22. holdingföretag med blandad verksamhet: ett moderföretag som inte är ett finansiellt holdingföretag, ett kreditinstitut eller ett blandat finansiellt holdingföretag i den mening som avses i direktiv 2002/87/EG, vilket har minst ett kreditinstitut bland sina dotterföretag.".
a) är dotterföretag till ett försäkringsföretag som är auktoriserat i gemenskapen,
De relevanta behöriga myndigheter som avses i första och andra stycket skall samråda med varandra särskilt när de bedömer aktieägarnas lämplighet och det goda anseendet och erfarenheten hos chefer som ingår i ledningen för en annan enhet i samma grupp. De skall till varandra överlämna alla uppgifter om aktieägarnas lämplighet och ledningens goda anseende och erfarenhet vilka är relevanta för övriga berörda behöriga myndigheter när det gäller att bevilja auktorisation samt fortlöpande bedöma efterlevnaden av uppställda verksamhetsvillkor.".
4. Artikel 34.2 skall ändras på följande sätt:
13. Fordringar med efterställd rätt till betalning och sådana instrument som avses i artikel 35 och artikel 36.3 som ett kreditinstitut innehar hos kreditinstitut och finansiella institut, i vilka kreditinstitutet har en ägarandel som i varje enskilt fall motsvarar mer än 10 % av kapitalet.
- försäkringsföretag i den mening som avses i artikel 6 i direktiv 73/239/EEG, artikel 6 i direktiv 79/267/EEG eller artikel 1 b i Europaparlamentets och rådets direktiv 98/78/EG(32),
16. Var och en av följande poster som ett kreditinstitut innehar i de enheter som definieras i punkt 15 i vilka det har ägarintresse
b) Andra stycket skall ersättas med följande:
Medlemsstaterna får föreskriva att kreditinstitut som är föremål för gruppbaserad tillsyn enligt kapitel 3 eller extra tillsyn enligt ovan nämnda direktiv 2002/87/EG, vid beräkning av den egna icke gruppbaserade kapitalbasen inte behöver dra ifrån poster enligt punkterna 15 och 16 i de kreditinstitut, finansiella institut eller försäkrings- eller återförsäkringsföretag eller försäkringsholdingföretag som omfattas av den gruppbaserade tillsynen eller av den extra tillsynen.
"3. Medlemsstaterna behöver inte tillämpa begränsningarna enligt punkterna 1 och 2 för ägarposter i försäkringsföretag enligt definitionen i direktiv 73/239/EEG och direktiv 79/267/EEG eller i återförsäkringsföretag enligt definitionen i direktiv 98/78/EG.".
7. Artikel 54 skall ändras på följande sätt:
b) I punkt 4 första stycket skall tredje strecksatsen utgå.
Ledningsorgan för finansiella holdingföretag
"Artikel 55a
De behöriga myndigheterna skall kräva att kreditinstituten följer adekvata metoder för riskhantering och rutiner för intern kontroll, inbegripet sunda rapporterings- och redovisningsförfaranden, för att på ett lämpligt sätt identifiera, mäta, övervaka och kontrollera transaktionerna med det holdingföretag med blandad verksamhet som är moderföretag och dess dotterföretag. De behöriga myndigheterna skall kräva att kreditinstituten rapporterar varje annan betydande transaktion med dessa enheter än den som avses i artikel 48. Dessa förfaranden och betydande transaktioner skall övervakas av de behöriga myndigheterna.
"Den behöriga myndighet som har framställt begäran får om den så önskar delta i kontrollen, om den inte själv utför den.".
Moderföretag i tredje land
Alternativt skall medlemsstaterna tillåta sina behöriga myndigheter att använda andra lämpliga metoder för tillsyn vilka uppfyller målen för den gruppbaserade tillsynen över kreditinstitut. De myndigheter som skulle vara ansvariga för gruppbaserad tillsyn måste enas om dessa metoder efter att ha samrått med andra berörda behöriga myndigheter. De behöriga myndigheterna kan särskilt kräva att det inrättas ett finansiellt holdingföretag med huvudkontor inom gemenskapen och tillämpa bestämmelserna om gruppbaserad tillsyn på det finansiella holdingföretagets ställning på gruppnivå. Metoderna måste uppfylla de mål för den gruppbaserade tillsynen som ställs upp i detta kapitel och rapporteras till de andra berörda behöriga myndigheterna och kommissionen.".
Artikel 30
a) tillämpningsområdet för gruppbaserad tillsyn av kreditinstitut eller värdepappersföretag och/eller tillämpningsområdet för extra tillsyn över sådana försäkringsföretag som ingår i en försäkringsgrupp, och
Om ett kapitalförvaltningsbolag utgör en del av ett finansiellt konglomerat skall hänvisningar till begreppet reglerad enhet och till begreppet behöriga myndigheter och relevanta behöriga myndigheter i detta direktiv anses inbegripa kapitalförvaltningsbolag respektive de behöriga myndigheter som ansvarar för tillsynen över kapitalförvaltningsbolag. Detta skall också tillämpas på sådana grupper som avses i första stycket a.
Artikel 31
- huruvida kapitalförvaltningsbolag bör omfattas av tillsynen på gruppnivå,
- hur ofta finansiella konglomerat skall beräkna kapitaltäckningskraven enligt artikel 6.2 och rapportera till samordnaren om betydande riskkoncentrationer enligt artikel 7.2.
Artikel 32
Artikel 33
Artikel 34
Kommissionens direktiv 2002/97/EG
(Text av betydelse för EES)
med beaktande av rådets direktiv 86/362/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på spannmål(1), senast ändrat genom kommissionens direktiv 2002/79/EG(2), särskilt artikel 10 i detta,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(5), senast ändrat genom kommissionens direktiv 2002/81/EG(6), särskilt artikel 4.1 f i detta, och
(2) Nämnda införande i bilaga I till direktiv 91/414/EEG av dessa verksamma ämnen grundades på en utvärdering av de uppgifter som lämnats in om det föreslagna användningsområdet. Uppgifterna om användningen har lämnats in av vissa medlemsstater i enlighet med artikel 4.1 f i direktiv 91/414/EEG. Tillgängliga uppgifter har nu gåtts igenom, och de har befunnits vara tillräckliga för att vissa gränsvärden för bekämpningsmedelsrester skall kunna fastställas.
(5) För att konsumenterna skall kunna skyddas från exponering av bekämpningsmedelsrester i eller på produkter som inte har godkänts, bör de provisoriska gränsvärden som fastställs motsvara den lägsta analytiska bestämningsgränsen för samtliga produkter som omfattas av direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG.
(8) Kommissionen anmälde utkastet till detta direktiv till Världshandelsorganisationen (WTO), vars synpunkter beaktats vid den slutliga utformningen av direktivet. Möjligheten att för import fastställa gränsvärden för bekämpningsmedelsrester för vissa särskilda kombinationer av bekämpningsmedel och grödor kommer att undersökas av kommissionen, förutsatt att relevanta data lämnas in.
Artikel 1
Artikel 2
Artikel 3
Medlemsstaterna skall senast den 30 juni 2003 sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv. De skall omedelbart underrätta kommissionen om detta.
Artikel 5
Detta beslut riktar sig till medlemsstaterna.
om ändring av rådets förordning (EEG) nr 3696/93 om den statistiska indelningen av produkter efter näringsgren (CPA) inom Europeiska ekonomiska gemenskapen
med beaktande av rådets förordning (EEG) nr 3696/93 av den 29 oktober 1993 om den statistiska indelningen av produkter efter näringsgren (CPA) inom Europeiska ekonomiska gemenskapen(1), ändrad genom kommissionens förordning (EG) nr 1232/98(2), särskilt artikel 5 b och artikel 6 i denna, och
(2) Med anledning av uppdateringen av den statistiska näringsgrensindelningen i gemenskapen (vanligen kallad NACE Rev. 1) är det nödvändigt att göra ändringar i CPA.
(5) Förordning (EEG) nr 3696/93 bör därför ändras.
Artikel 1
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om notering av priserna för färska och kylda slaktkroppar av får på gemenskapens representativa marknader
med beaktande av rådets förordning (EG) nr 2529/2001 av den 19 december 2001 om den gemensamma organisationen av marknaden för får- och getkött(1), särskilt artiklarna 20 och 24 i denna, och
(2) Enligt artikel 20 i förordning (EG) nr 2529/2001 skall medlemsstaterna registrera priserna på får och fårkött. Närmare bestämmelser för prisrapporteringen bör fastställas.
(5) I vissa medlemsstater grundar sig dessa priser på priserna för levande djur. I de fallen bör priserna räknas om med hjälp av lämpliga koefficienter. I de områden där det görs en individuell värdering av levande djur för att uppskatta den slaktade vikten, kan dock omräkningen baseras på denna värdering.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
2. Priserna skall vara de som noterats i de prisnoteringsområden som avses i artikel 12 i förordning (EG) nr 2529/2001 av medlemsstater som uppfyller kraven som infördes genom punkt 1. De skall vara grossistpriser som noteras av dessa medlemsstater på den eller de representativa marknaderna under den vecka som föregår den vecka då uppgifterna lämnas. Den eller de representativa marknaderna skall beslutas av medlemsstaterna som nämns ovan. Prisberäkningen skall grunda sig på marknadspriserna exklusive mervärdeskatt.
Då priset är noterat enligt olika kategorier av slaktkroppar skall priset på den representativa marknaden vara lika med genomsnittet, viktat med koefficienter som har fastställts av medlemstaten för att avspegla den relativa betydelsen av varje kategori, av de priser som har noterats för dessa kategorier under en period på sju dagar i grossistled.
I de områden där priserna noteras på grundval av en individuell uppskattning av vikten på slaktkroppen av lammet skall omräkningen grundas på denna värdering.
2. Priset i medlemsstaten skall vara genomsnittet av de priser som noteras på de aktuella marknaderna, viktat med koefficienter som avspeglar den relativa betydelsen av varje marknad eller av varje kategori.
Senast den 1 mars år 2002 skall medlemsstaterna meddela kommissionen:
c) De koefficienter för viktning och omräkning som avses i artiklarna 2 och 3.
Förordning (EEG) nr 1481/86 upphör att gälla.
Kommissionens förordning (EG) nr 538/2002
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
av följande skäl:
(3) Inga invändningar enligt artikel 7 i förordning (EEG) nr 2081/92 har framställts till kommissionen till följd av offentliggörandet i Europeiska gemenskapernas officiella tidning(3) av det produktnamn som anges i bilagan till den här förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 8 maj 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Genom förordning (EEG) nr 2019/93 inrättades för de mindre Egeiska öarna en ordning med stöd för bikupor med produktion av kvalitetshonung. Eftersom artikel 12 i förordningen i dess ändrade lydelse enligt förordning (EG) nr 442/2002 numera hänvisar till "sammanslutningar av producenter" bör följaktligen terminologin i kommissionens förordning (EG) nr 3063/93(3) anpassas.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fjäderfäkött och ägg.
3. Artikel 3 skall ändras på följande sätt:
4. I artikel 4 skall andra stycket utgå.
- Antal bikupor för vilka sammanslutningar av biodlare eller enskilda biodlare ansökt om och beviljats stöd."
7. Artikel 8 skall utgå.
Europaparlamentets och rådets förordning (EG) nr 1460/2002
(Text av betydelse för EES)
med beaktande av kommissionens förslag(1),
i enlighet med det förfarande som anges i artikel 251 i fördraget(4), och
(2) Vissa av de arbetsuppgifter som nu utförs på gemenskapsnivå eller nationell nivå skulle kunna utföras av ett specialiserat expertorgan. Det behövs tekniskt och vetenskapligt stöd och en fast engagerad sakkunskap på hög nivå för att gemenskapens lagstiftning på områdena för sjösäkerhet och förhindrande av förorening från fartyg skall tillämpas korrekt och för att tillämpningen av lagstiftningen skall kunna bevakas och befintliga åtgärders effektivitet utvärderas. Det finns därför ett behov av att inrätta en europeisk sjösäkerhetsbyrå (byrån) inom gemenskapens befintliga institutionsstruktur och befogenhetsfördelning.
(5) Byrån bör arbeta för att förbättra samarbetet mellan medlemsstaterna och utarbeta bra metoder och sprida kunskap om dessa i gemenskapen. Detta bör i sin tur leda till att sjösäkerhetssystemet i gemenskapen blir bättre och att risken för olyckor, förorening och dödsfall till sjöss minskar.
(8) När det gäller byråns avtalsrättsliga ansvar, som regleras av den lagstiftning som är tillämplig på det avtal som byrån ingått, bör domstolen vara behörig att träffa avgöranden med stöd av en skiljedomsklausul i avtalet. Domstolen skall också vara behörig i tvister som gäller byråns utomobligatoriska ersättningsansvar.
(11) För att garantera byråns fullständiga oberoende och självständighet anses det nödvändigt att den har en egen budget, där intäkterna främst utgörs av ett bidrag från gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
2. Byrån skall ge medlemsstaterna och kommissionen tekniskt och vetenskapligt stöd och tillhandahålla sakkunskap på hög nivå för att hjälpa dem att på ett korrekt sätt tillämpa gemenskapslagstiftningen på området för sjösäkerhet och förhindrande av förorening från fartyg, att bevaka genomförandet av denna och att utvärdera befintliga åtgärders effektivitet.
För att säkerställa att de mål som anges i artikel 1 uppnås på ett lämpligt sätt skall byrån utföra följande uppgifter:
i) kontrollera att hela gemenskapssystemet för hamnstatskontroll fungerar, eventuellt genom besök i medlemsstaterna, och föreslå kommissionen förbättringar av systemet,
c) Den skall i samarbete med medlemsstaterna
d) Den skall underlätta samarbetet mellan medlemsstaterna och kommissionen på det område som omfattas av direktiv 2002/59/EG. Den skall särskilt
e) Den skall underlätta samarbetet mellan medlemsstaterna och kommissionen vid utarbetandet, med beaktande av medlemsstaternas olika rättssystem, av en gemensam metod för utredning av sjöolyckor i enlighet med internationellt överenskomna principer, vid tillhandahållande av stöd till medlemsstaterna vid utredning av allvarliga sjöolyckor och vid analys av befintliga olycksrapporter.
Artikel 3
2. Byrån skall underrätta den berörda medlemsstaten om det planerade besöket, namnen på de bemyndigade tjänstemännen och vilken dag besöket skall inledas. De bemyndigade tjänstemännen skall genomföra besöket efter uppvisande av ett beslut från byråns verkställande direktör, där syftet och målet med besöket anges.
Öppenhet och skydd av information
3. Styrelsen skall fastställa de interna regler som är nödvändiga för tillämpningen av punkterna 1 och 2.
BYRÅNS ORGANISATION OCH VERKSAMHET
1. Byrån skall vara ett gemenskapsorgan. Den skall vara en juridisk person.
4. Byrån skall företrädas av den verkställande direktören.
1. Tjänsteföreskrifterna för tjänstemän i Europeiska gemenskaperna, anställningsvillkoren för övriga anställda i Europeiska gemenskaperna och bestämmelser som antagits gemensamt av Europeiska gemenskapernas institutioner för tillämpningen av tjänsteföreskrifterna och anställningsvillkoren skall gälla för byråns personal. Styrelsen skall i samförstånd med kommissionen utfärda nödvändiga tillämpningsföreskrifter.
Artikel 7
Artikel 8
2. Domstolen skall vara behörig att träffa avgöranden på grundval av skiljedomsklausuler i de avtal som ingåtts av byrån.
5. De anställdas personliga ansvar gentemot byrån skall regleras av bestämmelserna i de tjänsteföreskrifter eller de anställningsvillkor som gäller för dem.
1. Bestämmelserna i förordning nr 1 av den 15 april 1958 om vilka språk som skall användas i Europeiska ekonomiska gemenskapen(11) skall gälla för byrån.
Styrelsens inrättande och dess befogenheter
a) utnämna den verkställande direktören i enlighet med artikel 16,
d) senast den 31 oktober varje år, efter att ha beaktat kommissionens yttrande, anta byråns arbetsprogram för det kommande året och skicka det till medlemsstaterna, Europaparlamentet, rådet och kommissionen.
f) utarbeta förfaranden för de beslut som skall fattas av den verkställande direktören,
i) ha disciplinär bestämmanderätt över den verkställande direktören och de enhetschefer som avses i artikel 15.3,
Styrelsens sammansättning
2. Varje medlemsstat och kommissionen skall utse sina företrädare i styrelsen samt en suppleant, som skall företräda ledamoten i dennes frånvaro.
Artikel 12
2. Mandatperioden för ordföranden och vice ordföranden skall vara tre år och skall upphöra om uppdraget som styrelseledamot upphör. Mandatet skall kunna förnyas en gång.
1. Styrelsens ordförande skall sammankalla till styrelsens sammanträden.
4. Styrelsen får, om det är fråga om konfidentiella uppgifter eller intressekonflikter, besluta att ta upp särskilda frågor på sin dagordning utan närvaro av de ledamöter som har utsetts i sin egenskap av yrkesverksamma personer från de mest berörda sektorerna. Närmare regler för tillämpningen av denna bestämmelse får fastställas i arbetsordningen.
7. Styrelsens sekretariat skall tillhandahållas av byrån.
1. Styrelsen skall fatta sina beslut med två tredjedelars majoritet av alla ledamöter som har rösträtt.
3. Röstningsförfarandena skall fastställas utförligare i arbetsordningen, särskilt villkoren för en ledamot att agera på en annan ledamots vägnar.
1. Byrån skall ledas av den verkställande direktören, som skall vara fullständigt oavhängig i sin tjänsteutövning, utan att det påverkar kommissionens och styrelsens respektive befogenheter.
b) Han/hon skall efter att ha hört kommissionen besluta om genomförandet av sådana besök som avses i artikel 3, i enlighet med de riktlinjer som fastställts av styrelsen i enlighet med artikel 10.2 g.
e) Han/hon skall utöva de befogenheter i förhållande till personalen som anges i artikel 6.2.
Artikel 16
Den verkställande direktören kan avsättas av styrelsen enligt samma förfarande.
Tredje lands deltagande
KAPITEL III
Budget
b) eventuella bidrag från de tredjeländer som deltar i byråns arbete i enlighet med artikel 17,
3. Den verkställande direktören skall göra en beräkning av byråns intäkter och utgifter för påföljande budgetår och överlämna denna till styrelsen tillsammans med en tjänsteförteckning.
På grundval av detta budgetförslag skall kommissionen fastställa motsvarande beräkningar i det preliminära förslag till Europeiska unionens allmänna budget som den skall förelägga rådet enligt artikel 272 i fördraget. Ramarna för gemenskapens godkända budgetprognos för de kommande åren måste iakttas.
Genomförande och kontroll av budgeten
3. Den verkställande direktören skall senast den 31 mars varje år översända utförliga räkenskaper över intäkter och utgifter under föregående räkenskapsår till kommissionen, styrelsen och revisionsrätten.
Artikel 20
2. Byrån skall ansluta sig till det interinstitutionella avtalet av den 25 maj 1999 om interna utredningar som utförs av OLAF och skall utan dröjsmål utfärda lämpliga föreskrifter, som skall gälla all dess personal.
Finansiella bestämmelser
SLUTBESTÄMMELSER
1. Senast fem år efter det att byrån inlett sin verksamhet skall styrelsen beställa en oberoende extern utvärdering av förordningens tillämpning. Kommissionen skall tillhandahålla byrån all den information som denna anser sig behöva för att kunna genomföra denna utvärdering.
Artikel 23
Artikel 24
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
om hälsobestämmelser för animaliska biprodukter som inte är avsedda att användas som livsmedel
med beaktande av kommissionens förslag(1),
enligt förfarandet i artikel 251 i fördraget(3), mot bakgrund av det gemensamma utkast som förlikningskommittén godkände den 12 september 2002, och
(2) Den vetenskapliga styrkommittén har antagit flera yttranden i denna fråga sedan det direktivet antogs. Den viktigaste slutsatsen i dessa är att animaliska biprodukter från djur som vid en hälsobesiktning inte bedöms vara lämpliga för användning som livsmedel inte heller bör få komma in i näringskedjan för djur.
(5) Genom den internationella vetenskapliga konferens om kött- och benmjöl som kommissionen och Europaparlamentet arrangerade i Bryssel den 1-2 juli 1997, inleddes en debatt om produktionen av kött- och benmjöl och om dess användning som foder. Det framhölls vid denna konferens att den framtida politiken på området behövde diskuteras ytterligare. För att kunna skapa så bred offentlig debatt som möjligt om gemenskapens framtida foderlagstiftning, färdigställde kommissionen i november 1997 ett samrådsdokument om kött- och benmjöl. Efter detta samråd verkar det råda samsyn kring behovet av att ändra direktiv 90/667/EEG så att dess bestämmelser anpassas till de nya vetenskapliga rönen.
(8) Matavfall som innehåller produkter av animaliskt ursprung kan också vara en vektor för sjukdomsspridning. Allt matavfall från transportmedel i internationell trafik bör bortskaffas på ett säkert sätt. Matavfall som produceras inom gemenskapen bör inte användas för utfodring av produktionsdjur, med undantag av pälsdjur.
(11) Europaparlamentets och rådets direktiv 2000/76/EG av den 4 december 2000 om förbränning av avfall(6) skall inte tillämpas på förbränningsanläggningar om det avfall som hanteras endast består av slaktkroppar av djur. Det är nödvändigt att fastställa minimikrav för sådana förbränningsanläggningar för att skydda djurs och människors hälsa. I väntan på att gemenskapen skall införa dessa krav får medlemsstaterna anta miljölagar för sådana anläggningar. Mindre strikta krav bör tillämpas på förbränningsanläggningar med låg kapacitet, exempelvis sådana som är belägna på jordbruksföretag och krematorier för sällskapsdjur, eftersom det material som hanteras där utgör en lägre risk och för att undvika onödiga transporter av animaliska biprodukter.
(14) Undantag kan även vara lämpliga för att göra det möjligt att bortskaffa animaliska biprodukter på plats under övervakning. Kommissionen bör få den information som behövs för att kunna övervaka situationen och fastställa tillämpningsföreskrifter om så är lämpligt.
(17) Medlemsstaterna använder sig av ett stort antal system för finansiellt stöd för bearbetning, insamling, lagring och bortskaffande av animaliska biprodukter. För att detta inte skall påverka konkurrensvillkoren för jordbruksprodukter, är det nödvändigt att genomföra en undersökning på området och, vid behov, vidta lämpliga åtgärder på gemenskapsnivå.
(20) För att säkerställa att produkter som importeras från tredje land uppfyller hälsokrav som är minst likvärdiga med eller motsvarande dem som tillämpas i gemenskapen, bör det inrättas ett system för godkännande av tredje länder och anläggningar i dessa, liksom bestämmelser om gemenskapsinspektioner för att se till att villkoren för godkännande efterlevs. Import från tredje land av sällskapsdjursfoder och råvaror för sådant foder får göras på villkor som avviker från dem som gäller samma typer av material som producerats i gemenskapen, särskilt när det gäller de garantier som krävs beträffande restsubstanser som är förbjudna enligt rådets direktiv 96/22/EG av den 29 april 1996 om förbud mot användning av vissa ämnen med hormonell och tyreostatisk verkan samt av B-agonister vid animalieproduktion och om upphävande av direktiv 81/602/EEG, 88/146/EEG och 88/299/EEG(9). För att det skall vara möjligt att garantera att sådant sällskapsdjursfoder och sådana råvaror bara används i avsett syfte är det nödvändigt att fastställa kontrollåtgärder för import av sådant material som omfattas av dessa undantagsbestämmelser.
(23) Rådets direktiv 92/118/EEG av den 17 december 1992 om djurhälso- och hygienkrav för handel inom gemenskapen med produkter, som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A.I till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG, samt för import till gemenskapen av sådana produkter(10) syftar till att uppfylla ovannämnda mål.
(26) De berörda produkterna bör omfattas av bestämmelserna om veterinära kontroller, inklusive kontroller av experter från kommissionen, och av de skyddsåtgärder som anges i rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att fullborda den inre marknaden(11).
(29) För att kunna ta hänsyn till den tekniska och vetenskapliga utvecklingen bör ett nära och välfungerande samarbete mellan kommissionen och medlemsstaterna säkerställas inom ramen för den ständiga kommitté, som inrättats genom Europaparlamentets och rådets förordning (EG) nr 178/2002 av den 28 januari 2002 om allmänna principer och krav för livsmedelslagstiftning, om inrättande av Europeiska myndigheten för livsmedelssäkerhet och om förfaranden i frågor som gäller livsmedelssäkerhet(15).
a) insamling, transport, lagring, hantering, bearbetning och användning eller bortskaffande av animaliska biprodukter, så att dessa produkter inte innebär några risker för folk- eller djurhälsan,
a) Färskt sällskapsdjursfoder från detaljhandelsledet eller i anläggningar vid försäljningsställen, där styckning och lagring enbart sker i samband med försäljning direkt till konsumenten.
d) Färskt sällskapsdjursfoder som skall användas inom det ursprungliga jordbruksföretaget, om detta foder framställts från djur som slaktats inom detta företag i syfte att användas enbart för jordbrukaren och dennes familj, i enlighet med nationell lagstiftning (husbehovsslakt).
ii) är avsett som foder, eller
g) Transitering med båt eller flyg.
Definitioner
b) kategori 1-material: animaliska biprodukter som avses i artikel 4.
e) djur: alla ryggradsdjur och ryggradslösa djur (inklusive fiskar, kräldjur och groddjur).
h) sällskapsdjur: djur av sådana arter som, utan att användas som livsmedel, i normala fall hålls och föds upp av människor i annat syfte än användning som produktionsdjur.
k) handel: handel med varor mellan medlemsstaterna enligt artikel 23.2 i fördraget.
n) transmissibel spongiform encefalopati (TSE): alla typer av transmissibel spongiform encefalopati, utom de som förekommer hos människor.
Artikel 3
2. Medlemsstaterna får dock reglera import och utsläppande på marknaden av produkter som inte anges i bilagorna VII och VIII i sin nationella lagstiftning i väntan på att ett beslut skall fattas i enlighet med det förfarande som avses i artikel 33.2. De skall omedelbart informera kommissionen om de använder sig av den möjligheten.
a) Alla delar av kroppen, inklusive hudar och skinn, från följande djur:
iii) Andra djur än produktionsdjur och vilda djur, särskilt inbegripet sällskapsdjur, djurparksdjur och cirkusdjur.
b) i) Specificerat riskmaterial.
d) Allt animaliskt material som samlas in vid rening av avloppsvatten från bearbetningsanläggningar för kategori 1-material samt från andra lokaler där specificerat riskmaterial avlägsnas, inbegripet material som avskiljts genom siktning eller i sandfång, fett- och oljeblandningar, slam och material som avlägsnats från dessa anläggningars avloppssystem, utom i de fall då detta material inte innehåller specificerat riskmaterial eller delar av sådant material.
2. Kategori 1-material skall utan onödigt dröjsmål samlas in, transporteras bort och identifieras i enlighet med artikel 7, och skall, om inte annat föreskrivs i artiklarna 23 och 24,
c) med undantag av material som avses i punkt 1 a i och ii, bearbetas enligt bearbetningsmetod 1 i en bearbetningsanläggning som godkänts i enlighet med artikel 13, och då skall det därav uppkomna materialet märkas permanent, med lukt om detta är tekniskt möjligt, i enlighet med kapitel I i bilaga VI och slutligen bortskaffas som avfall genom nedgrävning på en deponi som godkänts i enlighet med rådets direktiv 1999/31/EG av den 26 april 1999 om deponering av avfall(20),
3. Mellanhantering eller mellanlagring av kategori 1-material får bara genomföras på hanteringsställen för kategori 1 som godkänts enligt artikel 10.
Kategori 2-material
b) Allt slags animaliskt material som samlats in vid rening av avloppssvatten från slakterier, utom sådana slakterier som omfattas av artikel 4.1 d, eller från bearbetningsanläggningar för kategori 2-material, inbegripet material som avskiljts genom siktning eller i sandfång, fett- och oljeblandningar, slam och material som avlägsnats från dessa anläggningars avloppssystem.
e) Djur och delar av djur, med undantag av dem som avses i artikel 4, som dött på annat sätt än genom slakt för användning som livsmedel, inbegripet djur som avlivats för att utrota någon epizootisk sjukdom.
2. Kategori 2-material skall utan onödigt dröjsmål samlas in, transporteras bort och identifieras i enlighet med artikel 7, och skall, om inte annat föreskrivs i artiklarna 23 och 24,
i) omedelbart bortskaffas som avfall genom förbränning eller samförbränning i en förbrännings- eller samförbränningsanläggning som godkänts i enlighet med artikel 12, eller,
i) när det gäller uppkommet proteinhaltigt material, användas som organiskt gödningsmedel eller jordförbättringsmedel i enlighet med eventuella krav som har fastställts enligt förfarandet i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén,
d) när det gäller material som kommer från fisk, ensileras eller komposteras i enlighet med bestämmelser som har antagits enligt förfarandet i artikel 33.2,
ii) användas på mark i enlighet med denna förordning, eller
g) bortskaffas med någon annan metod, eller användas på något annat sätt, i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2 efter samråd med den berörda vetenskapliga kommittén. Denna metod eller detta sätt får antingen komplettera eller ersätta dem som föreskrivs i punkterna a-f.
Artikel 6
a) Delar från slaktade djur som är tjänliga som livsmedel i enlighet med gemenskapslagstiftningen, men som av kommersiella skäl inte är avsedda som livsmedel.
d) Blod från andra djur än idisslare som slaktas i ett slakteri och som har genomgått en före slaktbesiktning där de befunnits lämpade för slakt för att användas som livsmedel i enlighet med gemenskapslagstiftningen.
g) Färsk mjölk från djur som inte visar några kliniska tecken på sådana sjukdomar som kan överföras till människor eller djur via produkten i fråga.
j) Skal, biprodukter från kläckerier samt biprodukter i form av knäckägg från djur som inte visat några kliniska tecken på sådana sjukdomar som kan överföras till människor eller djur via produkten i fråga.
2. Kategori 3-material skall utan onödigt dröjsmål samlas in, transporteras bort och identifieras i enlighet med artikel 7, och skall, om inte annat föreskrivs i artiklarna 23 och 24,
c) bearbetas i en bearbetningsanläggning som godkänts i enlighet med artikel 17,
f) omvandlas i en biogas- eller komposteringsanläggning som godkänts i enlighet med artikel 15,
i) bortskaffas med någon annan metod, eller användas på något annat sätt, i enlighet med bestämmelser som har fastställts enligt förfarandet i artikel 33.2, efter samråd med berörd vetenskaplig kommitté. Denna metod eller detta sätt får komplettera eller ersätta dem som föreskrivs i punkterna a-h.
Insamling, transport och lagring
3. Medlemsstaterna skall säkerställa ändamålsenliga arrangemang för att garantera att insamling och transport av kategori 1- och kategori 2-material genomförs i enlighet med bilaga II.
6. Medlemsstaterna får emellertid besluta att inte tillämpa bestämmelserna i denna artikel på naturgödsel som transporteras mellan två platser inom samma jordbruksföretag, eller mellan jordbruksföretag och användare som är etablerade i samma medlemsstat.
1. Animaliska biprodukter och bearbetade produkter får sändas till andra medlemsstater endast på de villkor som anges i punkterna 2-6.
a) åtföljas av ett handelsdokument eller, när det krävs enligt denna förordning, ett hälsointyg, och
5. När den behöriga myndigheten på bestämmelseorten underrättats om en sändning i enlighet med punkt 4, skall den underrätta den behöriga myndigheten på ursprungsorten om varje sändnings ankomst via Animo-systemet, eller med hjälp av någon annan överenskommen metod.
Register
Godkännande av hanteringsställen
a) uppfylla kraven i kapitel I i bilaga III,
d) kontrolleras av den behöriga myndigheten i enlighet med artikel 26.
b) kunna hantera och lagra kategori 3-material i enlighet med kapitel II del A i bilaga III,
Artikel 11
2. För att kunna godkännas skall en lagringsanläggning
Artikel 12
2. För att godkännas av den behöriga myndigheten för bortskaffande av animaliska biprodukter, skall en förbränningsanläggning eller samförbränningsanläggning med hög kapacitet som inte omfattas av direktiv 2000/76/EG uppfylla
c) kraven i kapitel III i bilaga IV beträffande utsläpp i vattnet,
f) bestämmelserna för onormala driftsförhållanden i kapitel VI i bilaga IV.
b) när den ligger på ett jordbruksföretag endast användas för bortskaffande av material från det jordbruksföretaget,
e) uppfylla kraven i kapitel V i bilaga IV beträffande restsubstanser,
4. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
Godkännande av bearbetningsanläggningar för kategori 1- och kategori 2-material
a) uppfylla kraven i kapitel I i bilaga V,
d) genomgå anläggningens egenkontroll på det sätt som föreskrivs i artikel 25,
3. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
1. Oleokemiska anläggningar skall godkännas av den behöriga myndigheten.
c) föra register över de uppgifter som erhållits genom de åtgärder som anges i punkt b så att de kan läggas fram för den behöriga myndigheten,
4. Godkännandet skall dras in omedelbart om villkoren för godkännandet inte längre är uppfyllda.
1. Biogas- och komposteringsanläggningar skall godkännas av den behöriga myndigheten.
b) hantera och bearbeta animaliska biprodukter i enlighet med kapitel II delarna B och C i bilaga VI,
e) säkerställa att rötrest och, om tillämpligt, kompost uppfyller de mikrobiologiska krav som anges i kapitel II del D i bilaga VI.
Allmänna djurhälsobestämmelser
a) kommer från ett jordbruksföretag, ett område, en del av ett område eller, när det gäller vattenbruksprodukter, från en fiskodling, en zon eller en del av en zon som inte är föremål för djurhälsorestriktioner som gäller de berörda djuren och produkterna; detta gäller särskilt restriktioner som införts i samband med åtgärder för sjukdomsbekämpning enligt gemenskapslagstiftningen eller restriktioner till följd av en allvarlig överförbar sjukdom som förtecknas i rådets direktiv 92/119/EEG av den 17 december 1992 om införande av allmänna gemenskapsåtgärder för bekämpning av vissa djursjukdomar och särskilda åtgärder mot vesikulär svinsjuka(22),
a) har framställts, hanterats, transporterats och lagrats avskilt från, eller vid andra tidpunkter än produkter som uppfyller alla djurhälsovillkor,
d) uppfyller de särskilda krav som anges i bilagorna VII och VIII, eller de närmare bestämmelser som skall fastställas i enlighet med förfarandet i artikel 33.2.
Godkännande av bearbetningsanläggningar för kategori 3-material
a) uppfylla kraven i kapitel I i bilaga V och kapitel I i bilaga VII,
d) genomgå anläggningens egenkontroll på det sätt som föreskrivs i artikel 25,
3. Godkännandet skall omedelbart återkallas om villkoren för godkännandet inte längre uppfylls.
1. Anläggningar för tillverkning av sällskapsdjursfoder och tekniska anläggningar skall godkännas av den behöriga myndigheten.
i) uppfylla de särskilda krav på produktionen som ställs i denna förordning,
iv) föra register över de uppgifter som erhållits i enlighet med ii och iii och hålla dem tillgängliga för den behöriga myndigheten. Resultaten från kontroller och tester skall sparas i minst två år,
3. Godkännandet skall omedelbart återkallas om villkoren för godkännandet inte längre uppfylls.
Medlemsstaterna skall se till att bearbetat animaliskt protein och andra bearbetade produkter som skulle kunna användas som foderråvara släpps ut på marknaden eller exporteras endast om de
c) har hanterats, bearbetats, lagrats och transporterats i enlighet med bilaga VII och på ett sådant sätt att det säkerställs att artikel 22 följs,
Utsläppande på marknaden och export av sällskapsdjursfoder, tuggben och tekniska produkter
i) uppfyller de särskilda kraven i bilaga VIII, eller
2. Medlemsstaterna skall se till att organiska gödningsmedel och jordförbättringsmedel som är framställda av bearbetade produkter, såvida de inte framställts av naturgödsel och mag- och tarminnehåll, släpps ut på marknaden eller exporteras endast om de uppfyller eventuella krav som fastställts i enlighet med det förfarande som avses i artikel 33.2, efter samråd med den berörda vetenskapliga kommittén.
b) har hanterats, bearbetats, lagrats och transporterats i enlighet med bilaga VI,
Skyddsåtgärder
Begränsningar i användningen
b) Utfodring av produktionsdjur, med undantag av pälsdjur, med matavfall eller foderråvara som innehåller eller framställts av matavfall.
Artikel 23
a) Användning av animaliska biprodukter för diagnostisk verksamhet samt i undervisnings- och forskningssyfte.
b) De animaliska biprodukter som avses i stycke a är följande:
c) De djur som avses i stycke a är följande:
iii) andra kräldjur och rovfåglar än djurparksdjur och cirkusdjur,
vi) hundar från etablerade kennlar eller grupper av sådana hundar som jakt- eller draghundar,
3. Medlemsstaterna skall informera kommissionen om
4. Varje medlemsstat skall upprätta en förteckning över de användare och uppsamlingscentraler i det egna landet som godkänts och registrerats i enlighet med punkt 2 c iv, vi och vii. Varje användare och uppsamlingscentral skall tilldelas ett officiellt nummer för kontrolländamål och för att produkterna i fråga skall kunna spåras till sitt ursprung.
5. Närmare bestämmelser om kontrollåtgärder får antas i enlighet med det förfarande som avses i artikel 33.2.
1. Den behöriga myndigheten får vid behov besluta att
i) kategori 1-material som avses i artikel 4.1 b ii,
c) animaliska biprodukter får bortskaffas som avfall genom förbränning eller nedgrävning på platsen vid utbrott av en sjukdom som anges i A-listan från Internationella byrån för epizootiska sjukdomar (OIE) om den behöriga myndigheten avvisar transport till närmaste förbrännings- eller bearbetningsanläggning på grund av risken för spridning av hälsorisker eller på grund av att ett omfattande utbrott av en epizootisk sjukdom leder till kapacitetsbrist på sådana anläggningar.
4. Medlemsstaterna skall informera kommissionen om
5. Den behöriga myndigheten skall vidta nödvändiga åtgärder för att
6. Närmare bestämmelser för genomförandet av denna artikel får fastställas i enlighet med förfarandet i artikel 33.2.
1. Ansvariga för eller ägare till hanteringsställen och bearbetningsanläggningar eller deras företrädare skall vidta alla nödvändiga åtgärder för att uppfylla kraven i denna förordning. De skall införa, genomföra och upprätthålla ett permanent förfarande som utarbetats i enlighet med principerna för systemet för riskbedömning och kritiska kontrollpunkter (HACCP). De skall särskilt
c) när det gäller bearbetningsanläggningar, ta representativa prov för att kontrollera att
d) föra register över resultaten av de kontroller och tester som avses i styckena b och c, och bevara dessa i minst två år, så att de behöriga myndigheterna kan ta del av dem,
a) omedelbart ge den behöriga myndigheten all relevant information om typen av prov och om det parti från vilket det tagits,
d) se till att inget material som konstaterats eller misstänks vara smittat avlägsnas från anläggningen innan det genomgått förnyad bearbetning under den behöriga myndighetens tillsyn samt förnyad officiell provtagning, så att kraven i denna förordning uppfylls, såvida det inte skall bortskaffas,
g) införa lämpliga dekontaminerings- och rengöringsmetoder på anläggningen.
Officiella kontroller och förteckningar över godkända anläggningar
3. Om de besiktningar som utförs av den behöriga myndigheten visar att ett eller flera krav i denna förordning inte har uppfyllts, skall den behöriga myndigheten vidta lämpliga åtgärder.
Artikel 27
Artikel 28
Det skall dock vara tillåtet att importera sällskapsdjursfoder och råvaror för produktion av sådant foder från tredje land även om detta foder och dessa råvaror kommer från djur som har behandlats med vissa ämnen som är förbjudna enligt direktiv 96/22/EG, under förutsättning att dessa råvaror är permanent märkta och i enlighet med vissa särskilda villkor, som fastställts i enlighet med förfarandet i artikel 33.2.
1. Det skall vara förbjudet att importera eller transitera animaliska biprodukter och bearbetade produkter om det inte sker i enlighet med denna förordning.
Förteckningen får samordnas med andra förteckningar som upprättats av folk- och djurhälsoskäl.
b) Hur den behöriga myndigheten i det tredje landet och dess inspektörer är organiserade, vilka befogenheter som inspektörerna har, vilken tillsyn inspektörerna är underkastade, samt inspektörernas behörighet att effektivt övervaka hur landets lagstiftning tillämpas.
e) Erfarenheter från saluföringen av produkten från det tredje landet samt resultaten av de införselkontroller som genomförts.
h) Hur snabbt och regelbundet det tredje landet tillhandahåller uppgifter om förekomsten av infektiösa eller smittsamma djursjukdomar på dess territorium, särskilt de sjukdomar som anges i OIE:s A-lista och B-lista eller, beträffande sjukdomar hos vattenbruksdjur, de anmälningspliktiga sjukdomar som förtecknas i OIE:s hälsokodex för vattenlevande djur.
Godkända förteckningar skall ändras enligt följande:
c) Om minst en medlemsstat har lämnat skriftliga synpunkter skall kommissionen inom fem arbetsdagar underrätta övriga medlemsstater om detta samt föra upp ärendet som en punkt på dagordningen till Ständiga kommitténs för livsmedelskedjan och djurhälsa nästa sammanträde för avgörande, i enlighet med förfarandet i artikel 33.2.
6. Sändningar av de produkter som avses i bilagorna VII och VIII skall, om inte något annat anges i dessa bilagor, åtföljas av ett hälsointyg som utformats enligt förlagan i bilaga X och som bestyrker att produkterna uppfyller de villkor som avses i dessa bilagor samt att de kommer från anläggningar som säkerställer att dessa villkor uppfylls.
Likvärdighet
2. De villkor som avses i punkt 1 skall omfatta
c) vid behov, förfaranden för att upprätta och ändra förteckningar över regioner eller anläggningar från vilka import och/eller transitering är tillåten.
Gemenskapens inspektioner och granskningar
b) kontrollera efterlevnaden av
iii) villkoren för erkännande av att åtgärder är likvärdiga,
2. De kontroller som avses i punkt 1 skall utföras på gemenskapens vägnar och på gemenskapens bekostnad.
Artikel 32
2. När det gäller förbudet mot utfodring med matavfall som fastställs i artikel 22 skall, i medlemsstater där lämpliga kontrollsystem finns innan denna förordning börjar tillämpas, övergångsåtgärder vidtas, i enlighet med första stycket, för att tillåta fortsatt användning av vissa typer av matavfall under noga kontrollerade förhållanden under en period på högst fyra år från och med den 1 november 2002. Genom åtgärderna skall det garanteras att det inte finns några onödiga risker för djurs hälsa eller folkhälsan under övergångsperioden.
1. Kommissionen skall biträdas av Ständiga kommittén för livsmedelskedjan och djurhälsa, nedan kallad "kommittén".
3. Kommittén skall själv anta sin arbetsordning.
Samråd skall genomföras med de berörda vetenskapliga kommittéerna i alla frågor inom denna förordnings tillämpningsområde som kan påverka människors eller djurs hälsa.
1. Medlemsstaterna skall till kommissionen överlämna texterna till nationell lagstiftning som de antar inom det område som omfattas av denna förordning.
Artikel 36
Artikel 37
Hänvisningar till direktiv 90/667/EEG skall från den dagen förstås som hänvisningar till denna förordning.
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om rättelse av förordning (EG) nr 1282/2002 om ändring av bilagorna till rådets direktiv 92/65/EEG om fastställande av djurhälsokrav i handeln inom och importen till gemenskapen av djur, sperma, ägg (ova) och embryon som inte faller under de krav som fastställs i de specifika gemenskapsregler som avses i bilaga A.I till direktiv 90/425/EEG
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Förordning (EG) nr 1282/2002 om ändring av direktiv 92/65/EEG antogs den 15 juli 2002.
(4) Förordning (EG) nr 1282/2002 bör därför rättas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 14 oktober 2002
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
(2) I artikel 13.1 i förordning (EG) nr 2200/96 fastställs att det datum då de två- och femåriga övergångsperioderna inleds skall vara det datum förordningen träder i kraft, dvs. den 21 november 1996. Detta är ett misstag; faktum är att det skulle ha varit meningslöst att låta övergångsåtgärder vara stödberättigande från och med datumet för ikraftträdande av förordning (EG) nr 2200/96, eftersom förordning (EEG) nr 1035/72 gällde fram till och med den 31 december 1996. Övergångsperioderna i fråga borde ha inletts i och med tillämpningsdatumet för förordning (EG) nr 2200/96.
Artikel 1
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EEG) nr 3149/92 om närmare bestämmelser för leverans av livsmedel från interventionslager till förmån för de sämst ställda i gemenskapen
med beaktande av rådets förordning (EEG) nr 3730/87 av den 10 december 1987 om allmänna bestämmelser för leverans av livsmedel från interventionslager till utsedda organisationer för utdelning till de sämst ställda i gemenskapen(1), ändrad genom förordning (EG) nr 2535/95(2), särskilt artikel 6 i denna, och
(2) I artikel 5 i förordning (EEG) nr 3149/92 fastställs bokföringsvärdet för de produkter som ställs till förfogande. Denna bestämmelse bör ändras för att hänsyn skall kunna tas till de ändringar som gjorts i interventionssystemet inom den gemensamma organisationen av marknaden för nötkött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 3.1 skall följande läggas till som andra stycke:"Uttag av produkter från interventionslagren skall ske från och med den 1 oktober till och med den 31 augusti följande år."
1. I EUGFJ:s (garantisektionen) bokföring, och utan att det påverkar tillämpningen av artikel 8 i förordning (EEG) nr 1883/78(5), skall bokföringsvärdet för de interventionsprodukter som ställs till förfogande enligt den här förordningen vara detsamma som gällande interventionspris den 1 oktober varje räkenskapsår.
2. Om interventionsprodukter transporteras från en medlemsstat till en annan skall den levererande medlemsstaten bokföra den levererade produkten till ett värde av noll, och destinationsmedlemsstaten skall bokföra produkten som intäkt under uttagsmånaden, till det pris som fastställs enligt punkt 1."
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om ändring av förordning (EG) nr 3223/94 om tillämpningsföreskrifter till importsystemet för frukt och grönsaker
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom förordning (EG) nr 545/2002(2), särskilt artikel 32.5 i denna, och
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för färsk frukt och färska grönsaker.
2. Åttonde strecksatsen skall ersättas med följande:
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS) och om ändring av förordningarna om sjösäkerhet och förhindrande av förorening från fartyg
med beaktande av kommissionens förslag(1),
i enlighet med förfarandet i artikel 251 i fördraget(4), och
(2) I sin resolution av den 8 juni 1993 om en gemensam politik för säkerhet till sjöss(7) godkände rådet i princip att det inrättas en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS) och uppmanade kommissionen att lägga fram ett förslag om att inrätta en sådan kommitté.
(5) Beslut 87/373/EEG har ersatts med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(8), vars bestämmelser bör tillämpas på COSS. Syftet med beslut 1999/468/EG är att fastställa tillämpliga kommittéförfaranden och att garantera mer uttömmande information till Europaparlamentet och allmänheten om kommittéernas arbete.
(8) Nämnda lagstiftning grundar sig på tillämpningen av regler som härrör från sådana internationella instrument som är i kraft vid tidpunkten för antagandet av den aktuella gemenskapsrättsakten eller vid en tidpunkt som anges i denna. Detta innebär att medlemsstaterna inte kan tillämpa senare ändringar av dessa internationella instrument, om inte gemenskapens direktiv eller förordningar ändras. Svårigheten att få tidpunkten för ikraftträdandet av ändringen på internationell nivå att sammanfalla med tidpunkten för ikraftträdandet av den förordning genom vilken ändringen infogas i gemenskapsrätten orsakar stora problem, och framför allt försenas tillämpningen av nyare och strängare internationella säkerhetsnormer inom gemenskapen.
(11) För insynens skull bör relevanta ändringar av de internationella instrument som är införlivade i gemenskapens sjöfartslagstiftning offentliggöras i gemenskapen genom Europeiska gemenskapernas officiella tidning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Syftet med denna förordning är att förbättra genomförandet av den gemenskapslagstiftning som avses i artikel 2.2 om sjösäkerhet, förhindrande av förorening från fartyg samt boende- och arbetsförhållanden ombord på fartyg genom att
Artikel 2
a) Rådets förordning (EEG) nr 613/91.
d) Rådets direktiv 94/57/EG av den 22 november 1994 om gemensamma regler och standarder för organisationer som utför inspektioner och utövar tillsyn av fartyg och för sjöfartsadministrationernas verksamhet i förbindelse därmed.(13)
g) Rådets direktiv 96/98/EG av den 20 december 1996 om marin utrustning.(15)
j) Rådets direktiv nr 98/41/EG av den 18 juni 1998 om registrering av personer som färdas ombord på passagerarfartyg som ankommer till eller avgår från hamnar i gemenskapens medlemsstater.(18)
m) Europaparlamentets och rådets direktiv 2001/25/EG av den 4 april 2001 om minimikrav på utbildning för sjöfolk.(21)
Artikel 3
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 4
Artikel 5
2. Ett förfarande för kontroll av överensstämmelse inrättas härmed i syfte att från tillämpningsområdet för gemenskapens sjöfartslagstiftning undanta en ändring av ett internationellt instrument endast om det, på grundval av en bedömning från kommissionens sida, finns en uppenbar risk att den internationella ändringen, inom ramen för tillämpningsområdet för de förordningar eller direktiv som avses i artikel 2.2, kommer att försämra den nivå på sjösäkerheten, förhindrandet av förorening från fartyg eller skydd av boende- och arbetsförhållandena ombord på fartyg som fastställs i gemenskapens sjöfartslagstiftning, eller vara oförenlig med denna lagstiftning.
Kommissionen skall snarast efter antagandet av en ändring av ett internationellt instrument för COSS lägga fram ett förslag till åtgärder som syftar till att undanta den aktuella ändringen från den gemenskapstext som berörs.
Artikel 6
Artikel 7
Artikel 8
1. Artikel 1 a skall ersättas med följande:
"Artikel 6
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara två månader.
Ändringarna av de internationella instrument som avses i artikel 1 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i förordning (EG) nr 2099/2002."
Förordning (EG) nr 2978/94 ändras på följande sätt:
2. Följande stycke skall läggas till i artikel 6:"Ändringarna av de internationella instrument som avses i artikel 3 får undantas från denna förordnings tillämpningsområde i enlighet med artikel 5 i Europaparlamentets och rådets förordning (EG) nr 2099/2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(25)."
1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i förordning (EG) nr 2099/2002.
3. Kommittén skall själv anta sin arbetsordning."
Förordning (EG) nr 3051/95 ändras på följande sätt:
"Artikel 10
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara två månader.
Ändring av förordning (EG) nr 417/2002
"1. Kommissionen skall biträdas av Kommittén för sjösäkerhet och förhindrande av förorening från fartyg (COSS), inrättad genom artikel 3 i Europaparlamentets och rådets förordning (EG) nr 2099/2002 av den 5 november 2002 om inrättande av en kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS)(29)."
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
om anpassning av rådets förordning (EG) nr 577/98 om anordnande av statistiska urvalsundersökningar av arbetskraften i gemenskapen och kommissionens förordning (EG) nr 1575/2000 om genomförande av rådets förordning (EG) nr 577/98 vad gäller förteckningen över variabler för utbildning samt deras kodning för användning vid överföring av data från och med 2003
med beaktande av rådets förordning (EG) nr 577/98 av den 9 mars 1998 om anordnande av statistiska urvalsundersökningar av arbetskraften i gemenskapen(1), ändrad genom Europarlamentets och rådets förordning (EG) nr 1991/2002(2), särskilt artikel 4.3 i denna, och
(2) Härav följer att koderna för dessa variabler enligt vad som anges i bilagan till kommissionens förordning (EG) nr 1575/2000 av den 19 juli 2000(3) också skall anpassas. Den nya förteckningen och kodningen skall genomföras redan under 2003 så att full kompatibilitet med ad hoc-modulen för 2003 om livslångt lärande(4) kan garanteras.
Artikel 1
deltagande i formell utbildning under de närmast föregående fyra veckorna
deltagande i kurser och annan undervisningsaktivitet under de närmast föregående fyra veckorna
- inriktning på den senaste undervisningsaktiviteten
- högsta nivå för med framgång avslutad utbildning
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
om tillämpning av rådets förordning (EEG) nr 1612/68 med avseende på förmedling av lediga platser och platsansökningar
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
av följande skäl:
(3) Med hänsyn till den kommande utvidgningen av Europeiska unionen bör införandet av EURES-nätverket i kandidatländerna beaktas i full utsträckning samtidigt som man ser till att systemet fortfarande är effektivt och hanterbart.
(6) Den yrkesmässiga och geografiska rörligheten behöver stimuleras i enlighet med den europeiska sysselsättningsstrategin med sikte på att genomföra handlingsplanen för kompetens och rörlighet(4) och rådets resolution av den 3 juni 2002 i samma fråga(5).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Kommissionen, medlemsstaternas arbetsförmedlingar och övriga nationella partner som de kan ha skall upprätta ett europeiskt nätverk för arbetsförmedlingar, som skall betecknas "EURES-nätverket" (EURopean Employment Services) och ansvara för utvecklingen av det informationsutbyte och samarbete som föreskrivs i del II i förordning (EEG) nr 1612/68.
EURES-nätverket skall bidra till en samordnad tillämpning av bestämmelserna i del II i förordning (EEG) nr 1612/68. Nätverket skall stödja den europeiska sysselsättningsstrategin och bidra till att stärka EU:s gemensamma marknad.
b) förmedling av lediga platser och platsansökningar mellan olika länder och regioner och i gränstrakter,
Artikel 3
a) EURES-medlemmar, som skall vara särskilda förmedlingar som medlemsstaterna utser enligt artikel 13.2 i förordning (EEG) nr 1612/68, och Europeiska samordningsbyrån, enligt artiklarna 21, 22 och 23 i den förordningen, och
ii) arbetsförmedlingar som ansvarar för gränstrakter,
Artikel 4
Europeiska samordningsbyrån (nedan kallad "EURES samordningsbyrå") skall övervaka iakttagandet av bestämmelserna i del II i förordning (EEG) nr 1612/68 och hjälpa nätverket att genomföra sin verksamhet.
b) utforma en samstämmig och övergripande metod samt lämpliga former för att främja samarbete och samordning mellan medlemsstaterna,
EURES-logotypen
Artikel 6
Kommissionen skall samråda med högnivågruppen i frågor som rör strategisk planering, utveckling, genomförande, övervakning och utvärdering när det gäller de tjänster och verksamheter som avses i det här beslutet, inklusive
c) kommissionens utkast till årsrapport som föreskrivs enligt artikel 19.1 i förordning (EEG) nr 1612/68,
Gruppen skall själv fastställa sina arbetsmetoder och anta sin arbetsordning. Gruppen skall sammankallas av ordföranden minst två gånger per år. Den skall anta sina yttranden med enkel majoritet.
Arbetsgrupp
EURES-stadga
a) Beskrivningar av den verksamhet som EURES medlemmar och samarbetspartner skall bedriva, vilket inbegriper
iii) främjande av en samordnad övervakning och bedömning av hinder för rörligheten, överskott och brist på kunskaper samt migrationsströmmar.
ii) typ av information, t.ex. information om arbetsmarknaden, levnad- och arbetsvillkor, lediga platser och platsansökningar samt hinder för rörlighet, som de måste lämna till sina kunder och till nätverket,
v) villkor för användning av EURES-logotypen för medlemmar och samarbetspartner,
Artikel 9
I riktlinjerna skall villkoren för det ekonomiska stöd som Europeiska gemenskapen kan lämna i enlighet med punkt 4 anges.
b) den personal och de ekonomiska resurser som tilldelats för tillämpningen av del II i förordning (EEG) nr 1612/68,
3. EURES samordningsbyrå skall granska verksamhetsplanerna och den information som lämnats om deras genomförande för att bedöma om de följer riktlinjerna och bestämmelserna i del II i förordning (EEG) nr 1612/68. Resultaten av denna bedömning skall granskas tillsammans med EURES-medlemmarna varje år i enlighet med artikel 19.1 i den förordningen samt inbegripas i den rapport som kommissionen vartannat år skall lämna till Europaparlamentet, rådet och Ekonomiska och sociala kommittén i enlighet med artikel 19.3 i den förordningen.
Upphävande
Datum för tillämpning
Adressater
av den 14 april 2003
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2 i detta,
efter att ha hört Regionkommittén,
(1) Genom rådets direktiv 98/18/EG av den 17 mars 1998 om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg(4) införs en enhetlig säkerhetsnivå för människoliv och egendom på nya och existerande passagerarfartyg och höghastighetspassagerarfartyg när dessa typer av fartyg används på inrikes resor, och fastställs förfaranden för förhandlingar på internationell nivå i syfte att harmonisera bestämmelserna för passagerarfartyg som används på internationella resor.
(4) Genom Europaparlamentets och rådets direktiv 2003/25/EG av den 14 april 2003 om särskilda stabilitetskrav för ro-ro-passagerarfartyg(5) införs skärpta stabilitetskrav för ro-ro-passagerarfartyg som går i internationell trafik till och från hamnar i gemenskapen; dessa krav bör även omfatta vissa kategorier av fartyg som går i inrikes trafik under motsvarande sjöförhållanden. Ro-ro-passagerarfartyg som inte uppfyller dessa stabilitetskrav bör tas ur trafik efter ett visst antal år i drift.
(7) Enligt direktiv 98/18/EG är den internationella säkerhetskoden för höghastighetsfartyg - fastställd i IMO:s sjösäkerhetskommittés resolution MSC 36 (63) av den 20 maj 1994 - tillämplig på alla höghastighetspassagerarfartyg som går i inrikes trafik. IMO har antagit en ny kod för höghastighetsfartyg - Internationella säkerhetskoden för höghastighetsfartyg 2000 (HSC-koden 2000), fastställd i IMO:s sjösäkerhetskommittés resolution MSC 97 (73) av den 5 december 2000 - som är tillämplig på alla höghastighetsfartyg byggda den 1 juli 2002 eller senare. Det är viktigt att se till att direktiv 98/18/EG kan uppdateras på ett flexibelt sätt så att sådan utveckling på internationell nivå kan tillämpas, även på höghastighetspassagerarfartyg som går i inrikes trafik.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. I artikel 2 skall följande punkter läggas till:
"w) personer med nedsatt rörlighet: alla personer som har särskilda problem med att använda allmänna transportmedel, inbegripet äldre, personer med funktionshinder, personer med sensoriska funktionshinder och rullstolsburna, gravida, och personer i sällskap med små barn."
a) fastställa och vid behov uppdatera en förteckning över de fartområden som omfattas av deras jurisdiktion och fastställa zonerna för åretrunttrafik och, i förekommande fall, begränsad periodisk trafik för de olika fartygsklasserna enligt klassificeringskriterierna i punkt 1,
3. Följande artiklar skall införas:
1. Ro-ro-passagerarfartyg i klasserna A-C som kölsträcks eller är på motsvarande byggnadsstadium den 1 oktober 2004 eller senare skall uppfylla artiklarna 6, 8 och 9 i Europaparlamentets och rådets direktiv 2003/25/EG av den 14 april 2003 om särskilda stabilitetskrav för ro-ro-passagerarfartyg(6).
Säkerhetskrav för personer med nedsatt rörlighet
3. När det gäller ombyggnaden av passagerarfartyg i klasserna A-D och höghastighetspassagerarfartyg som används för allmänna transporter och som kölsträcks eller befinner sig på motsvarande byggnadsstadium före den 1 oktober 2004, skall medlemsstaterna tillämpa riktlinjerna i bilaga III, i den mån det är rimligt och praktiskt möjligt i ekonomiskt hänseende.
4. Bilagan till detta direktiv skall läggas till som bilaga III.
Artikel 3
Artikel 4
om anpassning till den tekniska utvecklingen av Europaparlamentets och rådets direktiv 2000/30/EG i fråga om hastighetsbegränsande anordningar och avgasutsläpp från nyttofordon
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Direktiv 2000/30/EG rör den rättsliga ram för vägkontroller av nyttofordon, oavsett om de fraktar passagerare eller gods. Direktivet innehåller krav på att medlemsstaterna skall komplettera de årliga trafiksäkerhetsprovningarna med oanmälda vägkontroller av en representativ del av nyttofordonen varje år.
(4) De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från den kommitté för anpassning till den tekniska utvecklingen som inrättats genom artikel 8 i direktiv 96/96/EG.
Bilagorna I och II till direktiv 2000/30/EG ändras enligt bilagan till detta direktiv.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Europaparlamentets och rådets direktiv 2003/30/EG
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande(2),
av följande skäl:
(3) Det finns dock ett brett spektrum av biomassa som kan användas för att producera biodrivmedel och som härrör från jordbruks- och skogsbruksprodukter liksom från restprodukter och avfall från skogsbruk och skogs- och jordbrukslivsmedelsindustrin.
(6) En ökad användning av biodrivmedel utgör en del av det åtgärdspaket som krävs för att följa Kyotoprotokollet, liksom av andra strategier för att uppfylla ytterligare åtaganden i detta hänseende.
(9) Avgränsade fordonsflottor erbjuder möjligheten att använda biodrivmedel i högre koncentration. I vissa städer finns det redan avgränsade fordonsflottor som drivs med rent biodrivmedel, vilket i vissa fall har bidragit till att förbättra luftkvaliteten i städerna. Medlemsstaterna skulle därför ytterligare kunna främja användningen av biodrivmedel i offentliga transportmedel.
(12) Ren vegetabilisk olja från oljeväxter som framställs genom pressning, extraktion eller jämförbara metoder, rå eller raffinerad men kemiskt oförändrad, kan också användas som biodrivmedel i vissa fall där användningen är förenlig med motortyperna och motsvarande utsläppskrav.
(15) Att främja användningen av biodrivmedel i enlighet med hållbara jordbruks- och skogsbruksmetoder som föreskrivs i bestämmelserna inom den gemensamma jordbrukspolitiken kan skapa nya möjligheter till hållbar utveckling av landsbygden inom ramen för en mer marknadsinriktad gemensam jordbrukspolitik som är mer inriktad på den europeiska marknadens behov, en levande landsbygd och ett mångsidigare jordbruk och kan öppna en ny marknad för innovativa jordbruksprodukter i de nuvarande och framtida medlemsstaterna.
(18) Om alternativa drivmedel skall lyckas komma in på marknaden, måste de vara lättillgängliga och konkurrenskraftiga.
(21) Nationell politik för att främja användningen av biodrivmedel får inte hindra den fria rörligheten för drivmedel som uppfyller de harmoniserade miljöspecifikationerna i gemenskapslagstiftningen.
(24) Forskning och teknisk utveckling när det gäller biodrivmedlens hållbarhet bör främjas.
(27) Åtgärder bör vidtas för att snabbt utveckla kvalitetsstandarderna för biodrivmedel som används inom fordonssektorn, både som rena biodrivmedel och som blandningskomponenter i konventionella drivmedel. Även om den biologiskt nedbrytbara delen av avfall är en potentiellt användbar källa för framställning av biodrivmedel, måste det i kvalitetsstandarderna tas hänsyn till att avfallet eventuellt kan vara kontaminerat, så att inte vissa komponenter skadar fordonet eller förvärrar utsläppen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
b) biomassa: den biologiskt nedbrytbara delen av produkter, avfall och restprodukter från jordbruk (inklusive material av vegetabiliskt och animaliskt ursprung), skogsbruk och därmed förknippad industri, liksom den biologiskt nedbrytbara delen av industriavfall och kommunalt avfall,
2. Åtminstone de produkter som förtecknas nedan skall anses vara biodrivmedel:
c) biogas: en bränslegas som framställs av biomassa och/eller den biologiskt nedbrytbara delen av avfall som kan renas till naturgaskvalitet och som skall användas som biodrivmedel, eller vedgas.
f) bio-ETBE (etyltertiärbutyleter): ETBE som framställs av bioetanol. Volymandelen biodrivmedel i bio-ETBE beräknas till 47 %.
i) bioväte: vätgas som framställs av biomassa och/eller den biologiskt nedbrytbara delen av avfall, och som skall användas som biodrivmedel.
1. a) Medlemsstaterna bör se till att en minsta andel biodrivmedel och andra förnybara bränslen släpps ut på deras marknader och skall fastställa nationella vägledande mål för detta.
2. Biodrivmedel får tillhandahållas i följande form:
c) Vätskor som framställs av biodrivmedel, t.ex. ETBE (etyltertiärbutyleter), som innehåller den procentandel biodrivmedel som anges i artikel 2.2.
5. Medlemsstaterna skall se till att allmänheten upplyses om att biodrivmedel och andra förnybara drivmedel finns tillgängliga. Det skall föreskrivas att biodrivmedel som blandats i mineraloljederivat och som överstiger gränsvärdet på 5 % för fettsyrametylestrar (FAME) eller 5 % för bioetanol skall förses med en särskild märkning vid försäljningsställena.
- vilka åtgärder som vidtagits för att främja användningen av biodrivmedel eller andra förnybara drivmedel som skall ersätta diesel eller bensin för transportändamål,
I sin första rapport efter ikraftträdandet av detta direktiv skall medlemsstaterna ange nivån på sina nationella vägledande mål för den första fasen. I rapporten för år 2006 skall medlemsstaterna ange sina nationella vägledande mål för den andra fasen.
b) Storleken på de resurser som anslås till produktion av biomassa för annan energianvändning än transport samt de särskilda tekniska eller klimatmässiga förhållanden som kännetecknar den nationella marknaden för drivmedel.
Denna rapport skall åtminstone omfatta följande:
c) Biodrivmedel och andra förnybara drivmedel i ett livscykelperspektiv, för att ange möjliga åtgärder för det framtida främjandet av de av dem som är klimat- och miljövänliga och som kan bli konkurrenskraftiga och kostnadseffektiva.
f) En genomgång av ytterligare mer långsiktiga alternativ när det gäller åtgärder för energieffektivitet på transportområdet.
Förteckningen i artikel 2.2 får anpassas till den tekniska utvecklingen i enlighet med förfarandet i artikel 6.2. Vid anpassning av förteckningen skall biodrivmedlens inverkan på miljön beaktas.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Artikel 7
2. Medlemsstaterna skall till kommissionen överlämna texten till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 9
av den 18 juni 2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av rådets direktiv 86/362/EEG av den 24 juli 1986 om fastställande av gränsvärden för bekämpningsmedelsrester i och på spannmål(3), senast ändrat genom direktiv 2002/79/EG, särskilt artikel 10 i detta,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(7), senast ändrat genom kommissionens direktiv 2003/39/EG(8), särskilt artikel 4.1 f i detta, och
(2) De nya verksamma ämnena fenhexamid, acibenzolar-S-metyl, cyklanilid, pyraflufenetyl, iprovalikarb, prosulfuron, sulfosulfuron, cinidonetyl, cyhalofopbutyl, famoxadon, florasulam, metalaxyl-M, pikolinafen och flumioxazin infördes i bilaga I till direktiv 91/414/EEG genom kommissionens direktiv 2001/28/EG(12), 2001/87/EG(13), 2002/48/EG(14), 2002/64/EG(15) och 2002/81/EG(16).
(5) För de verksamma ämnena klorfenapyr, fentinacetat och fentinhydroxid fattades beslut om att inte införa dem i bilaga I till direktiv 91/414/EEG genom kommissionens direktiv 2001/697/EG(17), 2002/478/EG(18) respektive 2002/479/EG(19). I besluten föreskrivs att användningen av växtskyddsmedel som innehåller dessa verksamma ämnen inte längre skall vara tillåten i gemenskapen. Det är därför nödvändigt att alla bekämpningsmedelsrester som uppstår genom användning av dessa växtskyddsmedel läggs till i bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG för att möjliggöra en ordentlig övervakning och kontroll av förbuden mot användning och för att skydda konsumenterna.
(8) I samband med att de berörda verksamma ämnena infördes i eller uteslöts från bilaga I till direktiv 91/414/EEG avslutades de tekniska och vetenskapliga utvärderingarna genom kommissionens granskningsrapport. Utvärderingsrapporterna för de nämnda ämnena avslutades de datum som anges i de kommissions direktiv som anförs i skäl 1 och 2 samt i de kommissionsbeslut som anförs i skäl 5. I dessa rapporter fastställdes acceptabelt dagligt intag (ADI) och om nödvändigt akut referensdos (ARfD) för de berörda ämnena. Konsumenternas livstidsexponering genom livsmedel som behandlats med det berörda verksamma ämnet har uppskattats och utvärderats med hjälp av de metoder som används inom gemenskapen. Hänsyn har också tagits till de riktlinjer som offentliggjorts av Världshälsoorganisationen(20) samt yttrandet om de använda metoderna från den Vetenskapliga kommittén för växter(21). Slutsatsen har dragits att de föreslagna gränsvärdena inte leder till att acceptabla dagliga intag eller akuta referensdoser överskrids.
(11) Det är därför nödvändigt att förteckna samtliga de bekämpningsmedelsrester som härrör från användningen av dessa växtskyddsprodukter i bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG för att möjliggöra en ändamålsenlig övervakning och kontroll av användningsförbudet och för att skydda konsumenterna. Bilagorna till direktiv 86/362/EEG, 86/363/EEG och 90/642/EEG bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
De gränsvärden för bekämpningsmedelsrester som anges i bilagorna II och III till detta direktiv skall läggas till i del A och B i bilaga II till direktiv 86/363/EEG.
Artikel 5
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 7
av den 28 mars 2003
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Det är fel i de engelska och nederländska versionerna av kommissionens förordning (EG) nr 2603/1999(2), senast ändrad genom förordning (EG) nr 2055/2001(3). Dessa språkversioner bör därför rättas.
1. Rättelsen rör bara den nederländska versionen.
Kommissionens förordning (EG) nr 1053/2003
(Text av betydelse för EES)
med beaktande av Europaparlamentets och rådets förordning (EG) nr 999/2001 av den 22 maj 2001 om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati(1), senast ändrad genom kommissionens förordning (EG) nr 260/2003(2), särskilt första stycket i artikel 23 i denna, och
(2) I förordning (EG) nr 999/2001 fastställs även en förteckning över snabbtest som har godkänts för övervakning av TSE.
(5) För att garantera att godkända snabbtest håller samma prestandanivå efter godkännandet bör ett förfarande fastställas för eventuella ändringar av testet eller testprotokollet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 2
av den 27 juni 2003
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
(1) Förordning (EG) nr 999/2001 innehåller bestämmelser om övervakning av transmissibel spongiform encefalopati (TSE) hos får och getter, inklusive övervakning av ett urval av djur som inte slaktas för att användas som livsmedel. Det är nödvändigt att klargöra definitionen av denna grupp av djur för att undvika olämplig riktning av proven.
(4) I Vetenskapliga styrkommitténs yttrande av den 7 och 8 november 2002 om TSE-infektivitetens distribution i vävnader från idisslare rekommenderas att tonsiller från nötkreatur i alla åldrar bör anses medföra risk för BSE.
(7) Bestämmelserna om sändning av slaktkroppar, halva slaktkroppar och kvartsparter av slaktkroppar som inte innehåller annat specificerat riskmaterial än ryggraden till övriga medlemsstater utan deras förhandsgodkännande bör utvidgas till att omfatta halva slaktkroppar som styckats i högst tre grossistdelar för att återspegla den faktiska handeln mellan medlemsstater.
(10) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
Bilagorna III och XI till förordning (EG) nr 999/2001 skall ändras i enlighet med bilagan till denna förordning.
Europaparlamentets och rådets förordning (EG) nr 1267/2003
(Text av betydelse för EES)
med beaktande av kommissionens förslag(1),
av följande skäl:
(3) I rapporten betonades att man inom EMU kommer att behöva ägna större uppmärksamhet åt jämförelser mellan de olika ländernas arbetsmarknader.
(6) I handlingsplanen avseende den statistik som krävs i samband med den ekonomiska och monetära unionen, godkänd av Ekofin-rådet den 29 september 2000, fastställs att leverans av sysselsättningsuppgifter i nationalräkenskaperna i enheten "arbetade timmar" prioriteras.
Artikel 1
a) Texten till "Tabellöversikt" skall ersättas med texten i bilaga I.
Artikel 2
av den 30 oktober 2003
med beaktande av rådets förordning (EG) nr 3448/93 av den 6 december 1993 om systemet för handeln med vissa varor som framställs genom bearbetning av jordbruksprodukter(1), senast ändrad genom förordning (EG) nr 2580/2000(2), särskilt artikel 11.1 tredje stycket i denna, och
(2) Kommissionens förordning (EG) nr 1488/2001(5), bör ändras för att klargöra att de förfaranden som avses i artikel 16 i förordning (EG) nr 3448/93 är tillämpliga för att fastställa vilka basjordbruksprodukter som skall hänföras till förfarandet för aktiv förädling samt för att kontrollera och planera kvantiteterna av dessa produkter.
Artikel 1
"2. Om behoven av bidrag beräknas bli större än de tillgängliga ekonomiska medlen, skall kvantiteterna av de olika produkter som anges med sin åttasiffriga KN-kod, fastställas i enlighet med artikel 11.1 i förordning (EG) nr 3448/93 och med hjälp av prognosen."
"Artikel 24
av den 16 december 2003
med beaktande av Europaparlamentets och rådets förordning (EG) nr 2195/2002 av den 5 november 2002 om en gemensam terminologi vid offentlig upphandling (CPV)(1), särskilt artikel 2 i denna, och
(2) Uppbyggnaden av och koderna i CPV kan behöva anpassas, eller till och med ändras, i enlighet med marknadens utveckling och användarnas behov.
(5) I sitt yttrande(2) om förslaget till en förordning om CPV poängterade Regionkommittén att klassificeringen av läkemedel måste förbättras och rekommenderade att Världshälsoorganisationens klassificeringssystem, ATC (Anatomic Therapeutic Chemical), används för att komplettera CPV-systemet och dess koder för läkemedel.
(8) För tydlighetens skull bör CPV och konverteringstabellen mellan CPV och CPC Prov. ersättas i sin helhet. Alla ändringar i CPV-koderna eller i deras beskrivningar bör anges i en separat ny bilaga till förordning (EG) nr 2195/2002.
(11) Konverteringstabellen mellan CPV och CPA 96 i bilaga II till förordning (EG) nr 2195/2002 behöver därför inte uppdateras. Bilagan bör därför utgå.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Bilaga I skall ersättas med texten i bilaga I till denna förordning.
Bilaga IV skall ändras i enlighet med bilaga IV till denna förordning.
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
om antagande av undantag för Österrike, Frankrike och Luxemburg från bestämmelserna i Europaparlamentets och rådets förordning (EG) nr 2150/2002 om avfallsstatistik
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Frankrikes begäran av den 12 juni 2003,
(1) I enlighet med artikel 4.1 i förordning (EG) nr 2150/2002 får kommissionen under en övergångsperiod bevilja undantag från vissa bestämmelser i bilagorna till förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
a) Österrike beviljas undantag för redovisning av resultat avseende avsnitt 8.1.1, post 1 (jordbruk, jakt och skogsbruk) i bilaga I.
2. De undantag som beviljas i punkt 1 gäller endast uppgifter från det första referensåret, dvs. 2004.
Denna förordning träder i kraft den tjugonde dagen efter det att den offentliggjorts i Europeiska unionens officiella tidning.
